
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pc, property_invalid_acc, property_invalid_iram);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire [7:0] ACC_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [7:0] \oc8051_golden_model_1.n0994 ;
  wire [3:0] \oc8051_golden_model_1.n1071 ;
  wire [3:0] \oc8051_golden_model_1.n1073 ;
  wire [3:0] \oc8051_golden_model_1.n1075 ;
  wire [3:0] \oc8051_golden_model_1.n1076 ;
  wire [3:0] \oc8051_golden_model_1.n1077 ;
  wire [3:0] \oc8051_golden_model_1.n1078 ;
  wire [3:0] \oc8051_golden_model_1.n1079 ;
  wire [3:0] \oc8051_golden_model_1.n1080 ;
  wire [3:0] \oc8051_golden_model_1.n1081 ;
  wire \oc8051_golden_model_1.n1118 ;
  wire \oc8051_golden_model_1.n1146 ;
  wire [8:0] \oc8051_golden_model_1.n1147 ;
  wire [8:0] \oc8051_golden_model_1.n1148 ;
  wire [7:0] \oc8051_golden_model_1.n1149 ;
  wire \oc8051_golden_model_1.n1150 ;
  wire \oc8051_golden_model_1.n1151 ;
  wire [2:0] \oc8051_golden_model_1.n1152 ;
  wire \oc8051_golden_model_1.n1153 ;
  wire [1:0] \oc8051_golden_model_1.n1154 ;
  wire [7:0] \oc8051_golden_model_1.n1155 ;
  wire [15:0] \oc8051_golden_model_1.n1181 ;
  wire [7:0] \oc8051_golden_model_1.n1183 ;
  wire [8:0] \oc8051_golden_model_1.n1185 ;
  wire [8:0] \oc8051_golden_model_1.n1189 ;
  wire \oc8051_golden_model_1.n1190 ;
  wire [3:0] \oc8051_golden_model_1.n1191 ;
  wire [4:0] \oc8051_golden_model_1.n1192 ;
  wire [4:0] \oc8051_golden_model_1.n1196 ;
  wire \oc8051_golden_model_1.n1197 ;
  wire [8:0] \oc8051_golden_model_1.n1198 ;
  wire \oc8051_golden_model_1.n1206 ;
  wire [7:0] \oc8051_golden_model_1.n1207 ;
  wire [8:0] \oc8051_golden_model_1.n1211 ;
  wire \oc8051_golden_model_1.n1212 ;
  wire [4:0] \oc8051_golden_model_1.n1217 ;
  wire \oc8051_golden_model_1.n1218 ;
  wire \oc8051_golden_model_1.n1226 ;
  wire [7:0] \oc8051_golden_model_1.n1227 ;
  wire [8:0] \oc8051_golden_model_1.n1229 ;
  wire [8:0] \oc8051_golden_model_1.n1231 ;
  wire \oc8051_golden_model_1.n1232 ;
  wire [3:0] \oc8051_golden_model_1.n1233 ;
  wire [4:0] \oc8051_golden_model_1.n1234 ;
  wire [4:0] \oc8051_golden_model_1.n1236 ;
  wire \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1238 ;
  wire \oc8051_golden_model_1.n1245 ;
  wire [7:0] \oc8051_golden_model_1.n1246 ;
  wire [8:0] \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1257 ;
  wire [7:0] \oc8051_golden_model_1.n1258 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [4:0] \oc8051_golden_model_1.n1264 ;
  wire [4:0] \oc8051_golden_model_1.n1266 ;
  wire \oc8051_golden_model_1.n1267 ;
  wire [8:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire [7:0] \oc8051_golden_model_1.n1276 ;
  wire [4:0] \oc8051_golden_model_1.n1278 ;
  wire \oc8051_golden_model_1.n1279 ;
  wire [7:0] \oc8051_golden_model_1.n1280 ;
  wire [8:0] \oc8051_golden_model_1.n1282 ;
  wire \oc8051_golden_model_1.n1283 ;
  wire \oc8051_golden_model_1.n1290 ;
  wire [7:0] \oc8051_golden_model_1.n1291 ;
  wire [7:0] \oc8051_golden_model_1.n1292 ;
  wire [8:0] \oc8051_golden_model_1.n1295 ;
  wire [8:0] \oc8051_golden_model_1.n1296 ;
  wire [7:0] \oc8051_golden_model_1.n1297 ;
  wire \oc8051_golden_model_1.n1298 ;
  wire [7:0] \oc8051_golden_model_1.n1299 ;
  wire [7:0] \oc8051_golden_model_1.n1300 ;
  wire [8:0] \oc8051_golden_model_1.n1303 ;
  wire [8:0] \oc8051_golden_model_1.n1305 ;
  wire \oc8051_golden_model_1.n1306 ;
  wire [4:0] \oc8051_golden_model_1.n1307 ;
  wire [4:0] \oc8051_golden_model_1.n1309 ;
  wire \oc8051_golden_model_1.n1310 ;
  wire \oc8051_golden_model_1.n1317 ;
  wire [7:0] \oc8051_golden_model_1.n1318 ;
  wire [8:0] \oc8051_golden_model_1.n1322 ;
  wire \oc8051_golden_model_1.n1323 ;
  wire [4:0] \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1333 ;
  wire [7:0] \oc8051_golden_model_1.n1334 ;
  wire [8:0] \oc8051_golden_model_1.n1338 ;
  wire \oc8051_golden_model_1.n1339 ;
  wire [4:0] \oc8051_golden_model_1.n1341 ;
  wire \oc8051_golden_model_1.n1342 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire [7:0] \oc8051_golden_model_1.n1350 ;
  wire [8:0] \oc8051_golden_model_1.n1354 ;
  wire \oc8051_golden_model_1.n1355 ;
  wire [4:0] \oc8051_golden_model_1.n1357 ;
  wire \oc8051_golden_model_1.n1358 ;
  wire \oc8051_golden_model_1.n1365 ;
  wire [7:0] \oc8051_golden_model_1.n1366 ;
  wire \oc8051_golden_model_1.n1520 ;
  wire [6:0] \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [3:0] \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire [7:0] \oc8051_golden_model_1.n1555 ;
  wire [7:0] \oc8051_golden_model_1.n1680 ;
  wire \oc8051_golden_model_1.n1683 ;
  wire \oc8051_golden_model_1.n1685 ;
  wire \oc8051_golden_model_1.n1691 ;
  wire [7:0] \oc8051_golden_model_1.n1692 ;
  wire \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1698 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire \oc8051_golden_model_1.n1709 ;
  wire \oc8051_golden_model_1.n1711 ;
  wire \oc8051_golden_model_1.n1717 ;
  wire [7:0] \oc8051_golden_model_1.n1718 ;
  wire \oc8051_golden_model_1.n1722 ;
  wire \oc8051_golden_model_1.n1724 ;
  wire \oc8051_golden_model_1.n1730 ;
  wire [7:0] \oc8051_golden_model_1.n1731 ;
  wire \oc8051_golden_model_1.n1733 ;
  wire [7:0] \oc8051_golden_model_1.n1734 ;
  wire [7:0] \oc8051_golden_model_1.n1735 ;
  wire [15:0] \oc8051_golden_model_1.n1739 ;
  wire \oc8051_golden_model_1.n1745 ;
  wire [7:0] \oc8051_golden_model_1.n1746 ;
  wire \oc8051_golden_model_1.n1749 ;
  wire [7:0] \oc8051_golden_model_1.n1750 ;
  wire \oc8051_golden_model_1.n1765 ;
  wire [7:0] \oc8051_golden_model_1.n1766 ;
  wire \oc8051_golden_model_1.n1771 ;
  wire [7:0] \oc8051_golden_model_1.n1772 ;
  wire \oc8051_golden_model_1.n1777 ;
  wire [7:0] \oc8051_golden_model_1.n1778 ;
  wire \oc8051_golden_model_1.n1783 ;
  wire [7:0] \oc8051_golden_model_1.n1784 ;
  wire \oc8051_golden_model_1.n1789 ;
  wire [7:0] \oc8051_golden_model_1.n1790 ;
  wire [7:0] \oc8051_golden_model_1.n1791 ;
  wire [3:0] \oc8051_golden_model_1.n1792 ;
  wire [7:0] \oc8051_golden_model_1.n1793 ;
  wire [7:0] \oc8051_golden_model_1.n1828 ;
  wire \oc8051_golden_model_1.n1847 ;
  wire [7:0] \oc8051_golden_model_1.n1848 ;
  wire [7:0] \oc8051_golden_model_1.n1852 ;
  wire [3:0] \oc8051_golden_model_1.n1853 ;
  wire [7:0] \oc8051_golden_model_1.n1854 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff0 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff1 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff2 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff3 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_iram;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_42882_, rst);
  not (_18188_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_18199_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_18210_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _18199_);
  and (_18221_, _18210_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_18232_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _18199_);
  and (_18243_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _18199_);
  nor (_18254_, _18243_, _18232_);
  and (_18265_, _18254_, _18221_);
  nor (_18276_, _18265_, _18188_);
  and (_18287_, _18188_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18298_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_18309_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _18298_);
  nor (_18320_, _18309_, _18287_);
  not (_18331_, _18320_);
  and (_18342_, _18331_, _18265_);
  or (_18353_, _18342_, _18276_);
  and (_22216_, _18353_, _42882_);
  nor (_18374_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18385_, _18374_);
  and (_18396_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_18407_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_18418_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_18429_, _18418_);
  not (_18440_, _18309_);
  nor (_18451_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_18462_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_18473_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _18462_);
  nor (_18483_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_18494_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_18505_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _18494_);
  nor (_18516_, _18505_, _18483_);
  nor (_18527_, _18516_, _18473_);
  not (_18538_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_18549_, _18473_, _18538_);
  nor (_18560_, _18549_, _18527_);
  and (_18571_, _18560_, _18451_);
  not (_18582_, _18571_);
  and (_18593_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_18604_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_18615_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_18626_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _18615_);
  and (_18637_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_18648_, _18637_, _18604_);
  and (_18669_, _18648_, _18582_);
  nor (_18670_, _18669_, _18440_);
  not (_18681_, _18287_);
  nor (_18702_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_18703_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _18494_);
  nor (_18714_, _18703_, _18702_);
  nor (_18735_, _18714_, _18473_);
  not (_18736_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_18747_, _18473_, _18736_);
  nor (_18768_, _18747_, _18735_);
  and (_18769_, _18768_, _18451_);
  not (_18780_, _18769_);
  and (_18801_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_18802_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_18813_, _18802_, _18801_);
  and (_18834_, _18813_, _18780_);
  nor (_18835_, _18834_, _18681_);
  nor (_18845_, _18835_, _18670_);
  nor (_18866_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_18867_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _18494_);
  nor (_18878_, _18867_, _18866_);
  nor (_18889_, _18878_, _18473_);
  not (_18900_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_18911_, _18473_, _18900_);
  nor (_18922_, _18911_, _18889_);
  and (_18933_, _18922_, _18451_);
  not (_18944_, _18933_);
  and (_18955_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_18966_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_18977_, _18966_, _18955_);
  and (_18988_, _18977_, _18944_);
  nor (_18999_, _18988_, _18331_);
  nor (_19010_, _18999_, _18374_);
  and (_19021_, _19010_, _18845_);
  nor (_19032_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_19043_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _18494_);
  nor (_19054_, _19043_, _19032_);
  nor (_19065_, _19054_, _18473_);
  not (_19076_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_19087_, _18473_, _19076_);
  nor (_19098_, _19087_, _19065_);
  and (_19109_, _19098_, _18451_);
  not (_19120_, _19109_);
  and (_19131_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_19142_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_19153_, _19142_, _19131_);
  and (_19164_, _19153_, _19120_);
  and (_19175_, _19164_, _18374_);
  nor (_19185_, _19175_, _19021_);
  not (_19196_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19207_, _19196_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19218_, _19207_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19229_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_19240_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19251_, _19240_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19262_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_19272_, _19262_, _19229_);
  nor (_19283_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19294_, _19283_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19305_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_19316_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19327_, _19207_, _19316_);
  and (_19338_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_19349_, _19338_, _19305_);
  and (_19359_, _19349_, _19272_);
  and (_19370_, _19283_, _19196_);
  and (_19381_, _19370_, _19098_);
  and (_19392_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19403_, _19392_, _19316_);
  and (_19414_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_19425_, _19392_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19436_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_19446_, _19436_, _19414_);
  not (_19457_, _19446_);
  nor (_19468_, _19457_, _19381_);
  and (_19479_, _19468_, _19359_);
  not (_19490_, _19479_);
  and (_19501_, _19490_, _19185_);
  not (_19512_, _19501_);
  nor (_19522_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_19533_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _18494_);
  nor (_19544_, _19533_, _19522_);
  nor (_19555_, _19544_, _18473_);
  not (_19566_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_19577_, _18473_, _19566_);
  nor (_19588_, _19577_, _19555_);
  and (_19599_, _19588_, _18451_);
  not (_19609_, _19599_);
  and (_19620_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_19631_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_19642_, _19631_, _19620_);
  and (_19653_, _19642_, _19609_);
  nor (_19664_, _19653_, _18440_);
  nor (_19675_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_19686_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _18494_);
  nor (_19696_, _19686_, _19675_);
  nor (_19707_, _19696_, _18473_);
  not (_19718_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_19729_, _18473_, _19718_);
  nor (_19740_, _19729_, _19707_);
  and (_19751_, _19740_, _18451_);
  not (_19762_, _19751_);
  and (_19773_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_19783_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_19794_, _19783_, _19773_);
  and (_19805_, _19794_, _19762_);
  nor (_19816_, _19805_, _18681_);
  nor (_19827_, _19816_, _19664_);
  nor (_19838_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_19859_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _18494_);
  nor (_19871_, _19859_, _19838_);
  nor (_19883_, _19871_, _18473_);
  not (_19895_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_19907_, _18473_, _19895_);
  nor (_19919_, _19907_, _19883_);
  and (_19931_, _19919_, _18451_);
  not (_19932_, _19931_);
  and (_19943_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_19953_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_19964_, _19953_, _19943_);
  and (_19975_, _19964_, _19932_);
  nor (_19986_, _19975_, _18331_);
  nor (_19997_, _19986_, _18374_);
  and (_20008_, _19997_, _19827_);
  nor (_20019_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_20030_, _18494_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_20040_, _20030_, _20019_);
  nor (_20051_, _20040_, _18473_);
  not (_20062_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_20073_, _18473_, _20062_);
  nor (_20084_, _20073_, _20051_);
  and (_20095_, _20084_, _18451_);
  not (_20106_, _20095_);
  and (_20116_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_20127_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_20138_, _20127_, _20116_);
  and (_20149_, _20138_, _20106_);
  and (_20160_, _20149_, _18374_);
  nor (_20171_, _20160_, _20008_);
  and (_20182_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_20193_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_20203_, _20193_, _20182_);
  and (_20214_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_20225_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_20236_, _20225_, _20214_);
  and (_20247_, _20236_, _20203_);
  and (_20258_, _20084_, _19370_);
  and (_20269_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_20280_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_20290_, _20280_, _20269_);
  not (_20301_, _20290_);
  nor (_20312_, _20301_, _20258_);
  and (_20323_, _20312_, _20247_);
  not (_20334_, _20323_);
  and (_20345_, _20334_, _20171_);
  and (_20356_, _20345_, _19512_);
  not (_20366_, _20356_);
  and (_20377_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_20388_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_20399_, _20388_, _20377_);
  and (_20410_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_20421_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_20432_, _20421_, _20410_);
  and (_20443_, _20432_, _20399_);
  and (_20453_, _19740_, _19370_);
  and (_20464_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_20475_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_20486_, _20475_, _20464_);
  not (_20497_, _20486_);
  nor (_20508_, _20497_, _20453_);
  and (_20519_, _20508_, _20443_);
  not (_20530_, _20519_);
  and (_20541_, _20530_, _20171_);
  and (_20551_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_20562_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_20573_, _20562_, _20551_);
  and (_20584_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_20595_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_20606_, _20595_, _20584_);
  and (_20617_, _20606_, _20573_);
  and (_20628_, _19370_, _18768_);
  and (_20639_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_20649_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_20660_, _20649_, _20639_);
  not (_20671_, _20660_);
  nor (_20682_, _20671_, _20628_);
  and (_20693_, _20682_, _20617_);
  not (_20704_, _20693_);
  and (_20715_, _20704_, _19185_);
  and (_20726_, _20541_, _20715_);
  and (_20736_, _19490_, _20726_);
  nor (_20747_, _19501_, _20726_);
  nor (_20768_, _20747_, _20736_);
  and (_20779_, _20768_, _20541_);
  and (_20780_, _20345_, _19501_);
  and (_20791_, _19490_, _20171_);
  and (_20812_, _20334_, _19185_);
  nor (_20823_, _20812_, _20791_);
  nor (_20824_, _20823_, _20780_);
  and (_20844_, _20824_, _20779_);
  nor (_20855_, _20824_, _20779_);
  nor (_20856_, _20855_, _20844_);
  and (_20867_, _20856_, _20736_);
  nor (_20878_, _20867_, _20844_);
  nor (_20889_, _20878_, _20366_);
  and (_20910_, _20171_, _20704_);
  and (_20911_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_20921_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_20932_, _20921_, _20911_);
  and (_20943_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_20954_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_20965_, _20954_, _20943_);
  and (_20976_, _20965_, _20932_);
  and (_20987_, _19588_, _19370_);
  and (_20998_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_21009_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_21019_, _21009_, _20998_);
  not (_21040_, _21019_);
  nor (_21041_, _21040_, _20987_);
  and (_21052_, _21041_, _20976_);
  not (_21063_, _21052_);
  and (_21074_, _21063_, _19185_);
  and (_21085_, _21074_, _20910_);
  and (_21096_, _20530_, _19185_);
  nor (_21106_, _21096_, _20910_);
  nor (_21117_, _21106_, _20726_);
  and (_21128_, _21117_, _21085_);
  nor (_21139_, _19501_, _20541_);
  nor (_21150_, _21139_, _20779_);
  and (_21161_, _21150_, _21128_);
  nor (_21172_, _20856_, _20736_);
  nor (_21183_, _21172_, _20867_);
  and (_21194_, _21183_, _21161_);
  nor (_21214_, _21183_, _21161_);
  nor (_21215_, _21214_, _21194_);
  not (_21226_, _21215_);
  and (_21237_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_21248_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_21259_, _21248_, _21237_);
  and (_21270_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_21281_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_21291_, _21281_, _21270_);
  and (_21302_, _21291_, _21259_);
  and (_21313_, _19919_, _19370_);
  and (_21324_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_21335_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_21346_, _21335_, _21324_);
  not (_21357_, _21346_);
  nor (_21368_, _21357_, _21313_);
  and (_21379_, _21368_, _21302_);
  not (_21389_, _21379_);
  and (_21410_, _21389_, _20171_);
  and (_21411_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_21422_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_21433_, _21422_, _21411_);
  and (_21444_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_21455_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_21466_, _21455_, _21444_);
  and (_21476_, _21466_, _21433_);
  and (_21487_, _19370_, _18560_);
  and (_21498_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_21509_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_21520_, _21509_, _21498_);
  not (_21531_, _21520_);
  nor (_21542_, _21531_, _21487_);
  and (_21553_, _21542_, _21476_);
  not (_21564_, _21553_);
  and (_21574_, _21564_, _19185_);
  and (_21585_, _21574_, _21410_);
  and (_21596_, _21389_, _19185_);
  not (_21607_, _21596_);
  and (_21618_, _21564_, _20171_);
  and (_21629_, _21618_, _21607_);
  and (_21640_, _21629_, _21074_);
  nor (_21651_, _21640_, _21585_);
  and (_21661_, _21063_, _20171_);
  nor (_21672_, _21661_, _20715_);
  nor (_21683_, _21672_, _21085_);
  not (_21694_, _21683_);
  nor (_21705_, _21694_, _21651_);
  nor (_21716_, _21117_, _21085_);
  nor (_21727_, _21716_, _21128_);
  and (_21737_, _21727_, _21705_);
  nor (_21758_, _21150_, _21128_);
  nor (_21759_, _21758_, _21161_);
  and (_21770_, _21759_, _21737_);
  and (_21781_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_21792_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_21803_, _21792_, _21781_);
  and (_21814_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_21824_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_21835_, _21824_, _21814_);
  and (_21846_, _21835_, _21803_);
  and (_21867_, _19370_, _18922_);
  and (_21868_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_21879_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_21890_, _21879_, _21868_);
  not (_21901_, _21890_);
  nor (_21911_, _21901_, _21867_);
  and (_21922_, _21911_, _21846_);
  not (_21933_, _21922_);
  and (_21944_, _21933_, _20171_);
  and (_21955_, _21944_, _21596_);
  nor (_21966_, _21574_, _21410_);
  nor (_21977_, _21966_, _21585_);
  and (_21988_, _21977_, _21955_);
  nor (_21998_, _21629_, _21074_);
  nor (_22009_, _21998_, _21640_);
  and (_22020_, _22009_, _21988_);
  and (_22031_, _21694_, _21651_);
  nor (_22042_, _22031_, _21705_);
  and (_22053_, _22042_, _22020_);
  nor (_22064_, _21727_, _21705_);
  nor (_22075_, _22064_, _21737_);
  and (_22085_, _22075_, _22053_);
  nor (_22096_, _21759_, _21737_);
  nor (_22107_, _22096_, _21770_);
  and (_22118_, _22107_, _22085_);
  nor (_22129_, _22118_, _21770_);
  nor (_22140_, _22129_, _21226_);
  nor (_22151_, _22140_, _21194_);
  and (_22161_, _20878_, _20366_);
  nor (_22172_, _22161_, _20889_);
  not (_22183_, _22172_);
  nor (_22194_, _22183_, _22151_);
  or (_22205_, _22194_, _20780_);
  nor (_22217_, _22205_, _20889_);
  nor (_22228_, _22217_, _18429_);
  and (_22239_, _22217_, _18429_);
  nor (_22249_, _22239_, _22228_);
  not (_22260_, _22249_);
  and (_22271_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_22282_, _22183_, _22151_);
  nor (_22293_, _22282_, _22194_);
  and (_22314_, _22293_, _22271_);
  and (_22315_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_22325_, _22129_, _21226_);
  nor (_22336_, _22325_, _22140_);
  and (_22347_, _22336_, _22315_);
  nor (_22358_, _22336_, _22315_);
  nor (_22369_, _22358_, _22347_);
  not (_22380_, _22369_);
  and (_22391_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_22402_, _22107_, _22085_);
  nor (_22412_, _22402_, _22118_);
  and (_22423_, _22412_, _22391_);
  nor (_22434_, _22412_, _22391_);
  nor (_22445_, _22434_, _22423_);
  and (_22456_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_22467_, _22075_, _22053_);
  nor (_22478_, _22467_, _22085_);
  and (_22489_, _22478_, _22456_);
  nor (_22499_, _22478_, _22456_);
  nor (_22510_, _22499_, _22489_);
  not (_22521_, _22510_);
  and (_22532_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_22543_, _22042_, _22020_);
  nor (_22554_, _22543_, _22053_);
  and (_22565_, _22554_, _22532_);
  and (_22576_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_22586_, _22009_, _21988_);
  nor (_22607_, _22586_, _22020_);
  and (_22608_, _22607_, _22576_);
  and (_22619_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_22630_, _21977_, _21955_);
  nor (_22641_, _22630_, _21988_);
  and (_22652_, _22641_, _22619_);
  nor (_22662_, _22607_, _22576_);
  nor (_22673_, _22662_, _22608_);
  and (_22684_, _22673_, _22652_);
  nor (_22695_, _22684_, _22608_);
  not (_22716_, _22695_);
  nor (_22717_, _22554_, _22532_);
  nor (_22728_, _22717_, _22565_);
  and (_22739_, _22728_, _22716_);
  nor (_22749_, _22739_, _22565_);
  nor (_22760_, _22749_, _22521_);
  nor (_22771_, _22760_, _22489_);
  not (_22782_, _22771_);
  and (_22793_, _22782_, _22445_);
  nor (_22804_, _22793_, _22423_);
  nor (_22815_, _22804_, _22380_);
  nor (_22826_, _22815_, _22347_);
  nor (_22836_, _22293_, _22271_);
  nor (_22847_, _22836_, _22314_);
  not (_22858_, _22847_);
  nor (_22869_, _22858_, _22826_);
  nor (_22880_, _22869_, _22314_);
  nor (_22891_, _22880_, _22260_);
  nor (_22902_, _22891_, _22228_);
  not (_22913_, _22902_);
  and (_22933_, _22913_, _18407_);
  and (_22934_, _22933_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_22945_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_22956_, _22945_, _22934_);
  and (_22967_, _22956_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_22978_, _22967_, _18396_);
  not (_22989_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_23000_, _18374_, _22989_);
  or (_23011_, _23000_, _22978_);
  nand (_23022_, _22978_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  and (_23033_, _23022_, _23011_);
  and (_24374_, _23033_, _42882_);
  nor (_23053_, _18265_, _18298_);
  and (_23064_, _18265_, _18298_);
  or (_23075_, _23064_, _23053_);
  and (_02356_, _23075_, _42882_);
  and (_23096_, _21933_, _19185_);
  and (_02542_, _23096_, _42882_);
  nor (_23117_, _21944_, _21596_);
  nor (_23128_, _23117_, _21955_);
  and (_02695_, _23128_, _42882_);
  nor (_23149_, _22641_, _22619_);
  nor (_23159_, _23149_, _22652_);
  and (_02877_, _23159_, _42882_);
  nor (_23190_, _22673_, _22652_);
  nor (_23191_, _23190_, _22684_);
  and (_03117_, _23191_, _42882_);
  nor (_23212_, _22728_, _22716_);
  nor (_23223_, _23212_, _22739_);
  and (_03361_, _23223_, _42882_);
  and (_23244_, _22749_, _22521_);
  nor (_23255_, _23244_, _22760_);
  and (_03562_, _23255_, _42882_);
  nor (_23275_, _22782_, _22445_);
  nor (_23286_, _23275_, _22793_);
  and (_03757_, _23286_, _42882_);
  and (_23307_, _22804_, _22380_);
  nor (_23318_, _23307_, _22815_);
  and (_03954_, _23318_, _42882_);
  and (_23339_, _22858_, _22826_);
  nor (_23350_, _23339_, _22869_);
  and (_04054_, _23350_, _42882_);
  and (_23370_, _22880_, _22260_);
  nor (_23381_, _23370_, _22891_);
  and (_04147_, _23381_, _42882_);
  nor (_23402_, _22913_, _18407_);
  nor (_23413_, _23402_, _22933_);
  and (_04246_, _23413_, _42882_);
  and (_23434_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_23445_, _23434_, _22933_);
  nor (_23466_, _23445_, _22934_);
  and (_04345_, _23466_, _42882_);
  nor (_23476_, _22945_, _22934_);
  nor (_23487_, _23476_, _22956_);
  and (_04444_, _23487_, _42882_);
  and (_23508_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_23519_, _23508_, _22956_);
  nor (_23530_, _23519_, _22967_);
  and (_04542_, _23530_, _42882_);
  nor (_23551_, _22967_, _18396_);
  nor (_23562_, _23551_, _22978_);
  and (_04641_, _23562_, _42882_);
  and (_23582_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _18199_);
  nor (_23593_, _23582_, _18210_);
  not (_23604_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_23615_, _18232_, _23604_);
  and (_23626_, _23615_, _23593_);
  and (_23637_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_23648_, _23637_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_23658_, _23637_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_23669_, _23658_, _23648_);
  and (_00925_, _23669_, _42882_);
  and (_00956_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _42882_);
  not (_23700_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_23711_, _19975_, _23700_);
  and (_23722_, _19653_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23733_, _23722_, _23711_);
  nor (_23743_, _23733_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_23754_, _19805_, _23700_);
  and (_23765_, _20149_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_23776_, _23765_, _23754_);
  and (_23787_, _23776_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_23798_, _23787_, _23743_);
  nor (_23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_23820_, _23809_, _20323_);
  nor (_23830_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor (_23841_, _23830_, _23820_);
  not (_23852_, _23841_);
  and (_23863_, _18988_, _23700_);
  and (_23874_, _18669_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23895_, _23874_, _23863_);
  nor (_23896_, _23895_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_23907_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_23917_, _18834_, _23700_);
  and (_23928_, _19164_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23939_, _23928_, _23917_);
  nor (_23950_, _23939_, _23907_);
  nor (_23961_, _23950_, _23896_);
  nor (_23972_, _23961_, _23852_);
  and (_23983_, _23961_, _23852_);
  nor (_23994_, _23983_, _23972_);
  and (_24004_, _23809_, _19479_);
  nor (_24015_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor (_24026_, _24015_, _24004_);
  not (_24037_, _24026_);
  nor (_24048_, _19975_, _23700_);
  nor (_24059_, _24048_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24079_, _19653_, _23700_);
  and (_24080_, _19805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24091_, _24080_, _24079_);
  nor (_24102_, _24091_, _23907_);
  nor (_24113_, _24102_, _24059_);
  nor (_24124_, _24113_, _24037_);
  and (_24135_, _24113_, _24037_);
  nor (_24146_, _24135_, _24124_);
  not (_24157_, _24146_);
  and (_24167_, _23809_, _20519_);
  nor (_24178_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  nor (_24189_, _24178_, _24167_);
  not (_24200_, _24189_);
  nor (_24211_, _18988_, _23700_);
  nor (_24222_, _24211_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24233_, _18669_, _23700_);
  and (_24243_, _18834_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24254_, _24243_, _24233_);
  nor (_24265_, _24254_, _23907_);
  nor (_24276_, _24265_, _24222_);
  nor (_24287_, _24276_, _24200_);
  and (_24298_, _24276_, _24200_);
  and (_24309_, _23733_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24320_, _24309_);
  nor (_24330_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_24341_, _23809_, _20693_);
  nor (_24352_, _24341_, _24330_);
  and (_24363_, _24352_, _24320_);
  and (_24375_, _23895_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24386_, _24375_);
  and (_24397_, _23809_, _21052_);
  nor (_24408_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_24418_, _24408_, _24397_);
  and (_24429_, _24418_, _24386_);
  nor (_24440_, _24418_, _24386_);
  nor (_24451_, _24440_, _24429_);
  not (_24462_, _24451_);
  and (_24473_, _24048_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24484_, _24473_);
  and (_24495_, _23809_, _21553_);
  nor (_24505_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_24516_, _24505_, _24495_);
  and (_24527_, _24516_, _24484_);
  and (_24538_, _24211_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24549_, _24538_);
  nor (_24560_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and (_24571_, _23809_, _21379_);
  nor (_24581_, _24571_, _24560_);
  nor (_24592_, _24581_, _24549_);
  not (_24613_, _24592_);
  nor (_24614_, _24516_, _24484_);
  nor (_24625_, _24614_, _24527_);
  and (_24636_, _24625_, _24613_);
  nor (_24647_, _24636_, _24527_);
  nor (_24658_, _24647_, _24462_);
  nor (_24668_, _24658_, _24429_);
  nor (_24679_, _24352_, _24320_);
  nor (_24690_, _24679_, _24363_);
  not (_24701_, _24690_);
  nor (_24712_, _24701_, _24668_);
  nor (_24723_, _24712_, _24363_);
  nor (_24734_, _24723_, _24298_);
  nor (_24745_, _24734_, _24287_);
  nor (_24755_, _24745_, _24157_);
  nor (_24766_, _24755_, _24124_);
  not (_24777_, _24766_);
  and (_24788_, _24777_, _23994_);
  or (_24799_, _24788_, _23972_);
  and (_24810_, _20149_, _19164_);
  or (_24821_, _24810_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_24832_, _23939_);
  and (_24843_, _23776_, _24832_);
  nor (_24854_, _24254_, _24091_);
  and (_24865_, _24854_, _24843_);
  or (_24876_, _24865_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24887_, _24876_, _24821_);
  and (_24898_, _24887_, _24799_);
  and (_24909_, _24898_, _23798_);
  nor (_24920_, _24777_, _23994_);
  or (_24931_, _24920_, _24788_);
  and (_24942_, _24931_, _24909_);
  nor (_24953_, _24909_, _23841_);
  nor (_24964_, _24953_, _24942_);
  not (_24975_, _24964_);
  and (_24986_, _24964_, _23798_);
  not (_24997_, _23961_);
  nor (_25008_, _24909_, _24037_);
  and (_25018_, _24745_, _24157_);
  nor (_25029_, _25018_, _24755_);
  and (_25040_, _25029_, _24909_);
  or (_25051_, _25040_, _25008_);
  and (_25062_, _25051_, _24997_);
  nor (_25073_, _25051_, _24997_);
  nor (_25084_, _25073_, _25062_);
  not (_25095_, _25084_);
  not (_25106_, _24113_);
  nor (_25117_, _24909_, _24200_);
  nor (_25128_, _24298_, _24287_);
  nor (_25139_, _25128_, _24723_);
  and (_25160_, _25128_, _24723_);
  or (_25161_, _25160_, _25139_);
  and (_25172_, _25161_, _24909_);
  or (_25183_, _25172_, _25117_);
  and (_25194_, _25183_, _25106_);
  nor (_25205_, _25183_, _25106_);
  not (_25216_, _24276_);
  and (_25227_, _24701_, _24668_);
  or (_25238_, _25227_, _24712_);
  and (_25249_, _25238_, _24909_);
  nor (_25260_, _24909_, _24352_);
  nor (_25271_, _25260_, _25249_);
  and (_25282_, _25271_, _25216_);
  and (_25293_, _24647_, _24462_);
  nor (_25304_, _25293_, _24658_);
  not (_25315_, _25304_);
  and (_25326_, _25315_, _24909_);
  nor (_25337_, _24909_, _24418_);
  nor (_25348_, _25337_, _25326_);
  and (_25359_, _25348_, _24320_);
  nor (_25370_, _25348_, _24320_);
  nor (_25381_, _25370_, _25359_);
  not (_25391_, _25381_);
  nor (_25402_, _24625_, _24613_);
  nor (_25423_, _25402_, _24636_);
  not (_25424_, _25423_);
  and (_25435_, _25424_, _24909_);
  nor (_25446_, _24909_, _24516_);
  nor (_25457_, _25446_, _25435_);
  and (_25468_, _25457_, _24386_);
  not (_25479_, _24581_);
  and (_25490_, _24909_, _24538_);
  or (_25501_, _25490_, _25479_);
  nand (_25512_, _24909_, _24538_);
  or (_25523_, _25512_, _24581_);
  and (_25534_, _25523_, _25501_);
  nor (_25545_, _25534_, _24473_);
  and (_25556_, _25534_, _24473_);
  nor (_25567_, _25556_, _25545_);
  and (_25578_, _23809_, _21922_);
  nor (_25589_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_25600_, _25589_, _25578_);
  nor (_25611_, _25600_, _24549_);
  not (_25622_, _25611_);
  and (_25633_, _25622_, _25567_);
  nor (_25644_, _25633_, _25545_);
  nor (_25655_, _25457_, _24386_);
  nor (_25666_, _25655_, _25468_);
  not (_25677_, _25666_);
  nor (_25688_, _25677_, _25644_);
  nor (_25699_, _25688_, _25468_);
  nor (_25710_, _25699_, _25391_);
  nor (_25731_, _25710_, _25359_);
  nor (_25732_, _25271_, _25216_);
  nor (_25742_, _25732_, _25282_);
  not (_25753_, _25742_);
  nor (_25764_, _25753_, _25731_);
  nor (_25775_, _25764_, _25282_);
  nor (_25786_, _25775_, _25205_);
  nor (_25797_, _25786_, _25194_);
  nor (_25808_, _25797_, _25095_);
  or (_25819_, _25808_, _25062_);
  or (_25830_, _25819_, _24986_);
  and (_25841_, _25830_, _24887_);
  nor (_25852_, _25841_, _24975_);
  and (_25863_, _24986_, _24887_);
  and (_25874_, _25863_, _25819_);
  or (_25885_, _25874_, _25852_);
  and (_00976_, _25885_, _42882_);
  or (_25906_, _24964_, _23798_);
  and (_25917_, _25906_, _25841_);
  and (_02832_, _25917_, _42882_);
  and (_02844_, _24909_, _42882_);
  and (_02866_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _42882_);
  and (_02890_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _42882_);
  and (_02914_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _42882_);
  or (_25978_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_25989_, _23637_, rst);
  and (_02924_, _25989_, _25978_);
  not (_26010_, _25600_);
  and (_26021_, _25917_, _24538_);
  nor (_26032_, _26021_, _26010_);
  and (_26053_, _26021_, _26010_);
  or (_26054_, _26053_, _26032_);
  and (_02936_, _26054_, _42882_);
  nor (_26074_, _25917_, _25534_);
  nor (_26085_, _25622_, _25567_);
  nor (_26096_, _26085_, _25633_);
  and (_26107_, _26096_, _25917_);
  or (_26118_, _26107_, _26074_);
  and (_02948_, _26118_, _42882_);
  and (_26139_, _25677_, _25644_);
  or (_26150_, _26139_, _25688_);
  nand (_26161_, _26150_, _25917_);
  or (_26172_, _25917_, _25457_);
  and (_26183_, _26172_, _26161_);
  and (_02960_, _26183_, _42882_);
  and (_26204_, _25699_, _25391_);
  or (_26215_, _26204_, _25710_);
  nand (_26226_, _26215_, _25917_);
  or (_26237_, _25917_, _25348_);
  and (_26248_, _26237_, _26226_);
  and (_02971_, _26248_, _42882_);
  and (_26269_, _25753_, _25731_);
  or (_26280_, _26269_, _25764_);
  nand (_26291_, _26280_, _25917_);
  or (_26302_, _25917_, _25271_);
  and (_26313_, _26302_, _26291_);
  and (_02984_, _26313_, _42882_);
  or (_26334_, _25205_, _25194_);
  and (_26345_, _26334_, _25775_);
  nor (_26356_, _26334_, _25775_);
  or (_26367_, _26356_, _26345_);
  nand (_26378_, _26367_, _25917_);
  or (_26389_, _25917_, _25183_);
  and (_26400_, _26389_, _26378_);
  and (_02997_, _26400_, _42882_);
  and (_26420_, _25797_, _25095_);
  or (_26431_, _26420_, _25808_);
  nand (_26442_, _26431_, _25917_);
  or (_26453_, _25917_, _25051_);
  and (_26464_, _26453_, _26442_);
  and (_03011_, _26464_, _42882_);
  not (_26485_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_26496_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _18199_);
  and (_26507_, _26496_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_26528_, _26507_, _26485_);
  and (_26529_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_26540_, _26529_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_26551_, _26529_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_26562_, _26551_, _26540_);
  and (_26573_, _26562_, _26528_);
  not (_26584_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_26595_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _18199_);
  and (_26606_, _26595_, _26485_);
  and (_26617_, _26606_, _26584_);
  and (_26628_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_26639_, _26628_, _26573_);
  not (_26650_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_26661_, _26496_, _26650_);
  and (_26672_, _26661_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_26683_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_26694_, _26661_, _26485_);
  and (_26705_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or (_26716_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_26727_, _26716_, _18199_);
  nor (_26738_, _26727_, _26496_);
  and (_26759_, _26738_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_26760_, _26759_, _26705_);
  nor (_26771_, _26760_, _26683_);
  and (_26781_, _26771_, _26639_);
  and (_26792_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor (_26803_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_26814_, _26803_, _26529_);
  and (_26825_, _26814_, _26528_);
  nor (_26836_, _26825_, _26792_);
  and (_26847_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_26858_, _26738_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_26869_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_26880_, _26869_, _26858_);
  nor (_26891_, _26880_, _26847_);
  and (_26902_, _26891_, _26836_);
  and (_26913_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_26924_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_26935_, _26924_, _26913_);
  and (_26946_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not (_26957_, _26946_);
  not (_26968_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_26979_, _26528_, _26968_);
  and (_26990_, _26738_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_27001_, _26990_, _26979_);
  and (_27012_, _27001_, _26957_);
  and (_27023_, _27012_, _26935_);
  and (_27034_, _27023_, _26902_);
  and (_27045_, _27034_, _26781_);
  and (_27056_, _26540_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_27067_, _27056_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_27078_, _27067_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_27089_, _27078_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_27100_, _27089_);
  not (_27111_, _26528_);
  nor (_27122_, _27078_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_27132_, _27122_, _27111_);
  and (_27143_, _27132_, _27100_);
  not (_27154_, _27143_);
  and (_27165_, _26507_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27176_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_27187_, _27176_, _27165_);
  and (_27198_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_27209_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_27220_, _27209_, _27198_);
  and (_27231_, _27220_, _27187_);
  and (_27242_, _27231_, _27154_);
  nor (_27253_, _27067_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_27264_, _27253_);
  nor (_27275_, _27078_, _27111_);
  and (_27286_, _27275_, _27264_);
  not (_27297_, _27286_);
  and (_27308_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_27319_, _27308_, _27165_);
  and (_27340_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_27341_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_27352_, _27341_, _27340_);
  and (_27363_, _27352_, _27319_);
  and (_27374_, _27363_, _27297_);
  nor (_27385_, _27374_, _27242_);
  not (_27396_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_27407_, _27089_, _27396_);
  and (_27418_, _27089_, _27396_);
  nor (_27429_, _27418_, _27407_);
  nor (_27440_, _27429_, _27111_);
  not (_27451_, _27440_);
  and (_27462_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_27473_, _27462_);
  not (_27483_, _27165_);
  and (_27494_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_27505_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_27516_, _27505_, _27494_);
  and (_27527_, _27516_, _27483_);
  and (_27538_, _27527_, _27473_);
  and (_27549_, _27538_, _27451_);
  not (_27560_, _27549_);
  and (_27571_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_27582_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_27593_, _27582_, _27571_);
  not (_27604_, _27056_);
  nor (_27615_, _26540_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_27626_, _27615_, _27111_);
  and (_27637_, _27626_, _27604_);
  and (_27648_, _26738_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_27659_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_27670_, _27659_, _27648_);
  not (_27681_, _27670_);
  nor (_27692_, _27681_, _27637_);
  and (_27703_, _27692_, _27593_);
  not (_27714_, _27703_);
  and (_27725_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_27736_, _27725_, _27165_);
  nor (_27747_, _27056_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_27758_, _27747_, _27111_);
  nor (_27769_, _27758_, _27067_);
  and (_27780_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_27791_, _27780_, _27769_);
  and (_27801_, _27791_, _27736_);
  and (_27812_, _26738_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_27823_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_27834_, _27823_, _27812_);
  and (_27845_, _27834_, _27801_);
  nor (_27856_, _27845_, _27714_);
  and (_27867_, _27856_, _27560_);
  and (_27878_, _27867_, _27385_);
  nand (_27889_, _27878_, _27045_);
  and (_27900_, _25885_, _23626_);
  not (_27911_, _27900_);
  and (_27922_, _23033_, _18265_);
  not (_27933_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_27944_, _18210_, _27933_);
  and (_27955_, _27944_, _18254_);
  not (_27976_, _27955_);
  nor (_27977_, _20323_, _20149_);
  and (_27988_, _20323_, _20149_);
  nor (_27999_, _27988_, _27977_);
  not (_28010_, _19164_);
  nor (_28021_, _19479_, _28010_);
  nor (_28032_, _19479_, _19164_);
  and (_28043_, _19479_, _19164_);
  nor (_28054_, _28043_, _28032_);
  not (_28065_, _19805_);
  nor (_28076_, _20519_, _28065_);
  nor (_28087_, _20519_, _19805_);
  and (_28098_, _20519_, _19805_);
  nor (_28109_, _28098_, _28087_);
  not (_28120_, _18834_);
  and (_28130_, _20693_, _28120_);
  nor (_28141_, _28130_, _28109_);
  nor (_28152_, _28141_, _28076_);
  nor (_28163_, _28152_, _28054_);
  nor (_28174_, _28163_, _28021_);
  and (_28185_, _28152_, _28054_);
  nor (_28196_, _28185_, _28163_);
  not (_28207_, _28196_);
  and (_28218_, _28130_, _28109_);
  nor (_28229_, _28218_, _28141_);
  not (_28240_, _28229_);
  nor (_28251_, _20693_, _18834_);
  and (_28262_, _20693_, _18834_);
  nor (_28283_, _28262_, _28251_);
  not (_28284_, _28283_);
  and (_28295_, _21052_, _19653_);
  nor (_28306_, _21052_, _19653_);
  nor (_28317_, _28306_, _28295_);
  not (_28328_, _28317_);
  nor (_28339_, _21553_, _18669_);
  and (_28350_, _21553_, _18669_);
  nor (_28361_, _28350_, _28339_);
  nor (_28372_, _21379_, _19975_);
  and (_28383_, _21379_, _19975_);
  nor (_28394_, _28383_, _28372_);
  not (_28405_, _18988_);
  and (_28416_, _21922_, _28405_);
  nor (_28427_, _28416_, _28394_);
  not (_28437_, _19975_);
  nor (_28448_, _21379_, _28437_);
  nor (_28459_, _28448_, _28427_);
  nor (_28470_, _28459_, _28361_);
  not (_28481_, _18669_);
  nor (_28492_, _21553_, _28481_);
  nor (_28503_, _28492_, _28470_);
  nor (_28514_, _28503_, _28328_);
  and (_28525_, _28503_, _28328_);
  nor (_28536_, _28525_, _28514_);
  and (_28547_, _28459_, _28361_);
  nor (_28558_, _28547_, _28470_);
  not (_28569_, _28558_);
  nor (_28580_, _21922_, _18988_);
  and (_28591_, _21922_, _18988_);
  nor (_28602_, _28591_, _28580_);
  not (_28613_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_28634_, _18473_, _28613_);
  not (_28635_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_28646_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28657_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _28646_);
  and (_28668_, _28657_, _19696_);
  nor (_28679_, _28668_, _28635_);
  nor (_28690_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28701_, _28690_, _18714_);
  not (_28712_, _28701_);
  and (_28723_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28733_, _28723_, _20040_);
  not (_28744_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_28755_, _28744_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28766_, _28755_, _19054_);
  nor (_28777_, _28766_, _28733_);
  and (_28788_, _28777_, _28712_);
  and (_28799_, _28788_, _28679_);
  and (_28810_, _28657_, _19871_);
  nor (_28821_, _28810_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_28832_, _28755_, _18516_);
  not (_28843_, _28832_);
  and (_28854_, _28723_, _19544_);
  and (_28865_, _28690_, _18878_);
  nor (_28876_, _28865_, _28854_);
  and (_28887_, _28876_, _28843_);
  and (_28898_, _28887_, _28821_);
  nor (_28909_, _28898_, _28799_);
  nor (_28920_, _28909_, _18473_);
  nor (_28931_, _28920_, _28634_);
  and (_28942_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_28953_, _28942_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_28964_, _28953_);
  and (_28975_, _28964_, _28931_);
  and (_28986_, _28964_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_29007_, _28986_, _28975_);
  nor (_29008_, _29007_, _28602_);
  and (_29019_, _28416_, _28394_);
  nor (_29030_, _29019_, _28427_);
  not (_29040_, _29030_);
  and (_29051_, _29040_, _29008_);
  and (_29062_, _29051_, _28569_);
  and (_29073_, _29062_, _28536_);
  not (_29084_, _19653_);
  or (_29095_, _21052_, _29084_);
  and (_29106_, _21052_, _29084_);
  or (_29117_, _28503_, _29106_);
  and (_29128_, _29117_, _29095_);
  or (_29139_, _29128_, _29073_);
  and (_29150_, _29139_, _28284_);
  and (_29161_, _29150_, _28240_);
  and (_29172_, _29161_, _28207_);
  nor (_29183_, _29172_, _28174_);
  nor (_29194_, _29183_, _27999_);
  and (_29205_, _29183_, _27999_);
  nor (_29216_, _29205_, _29194_);
  nor (_29227_, _29216_, _27976_);
  not (_29238_, _29227_);
  not (_29249_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_29260_, _23582_, _29249_);
  and (_29271_, _29260_, _18254_);
  not (_29282_, _27999_);
  not (_29293_, _28054_);
  and (_29304_, _28251_, _28109_);
  nor (_29315_, _29304_, _28087_);
  nor (_29326_, _29315_, _29293_);
  not (_29337_, _28361_);
  and (_29347_, _28580_, _28394_);
  nor (_29358_, _29347_, _28372_);
  nor (_29369_, _29358_, _29337_);
  nor (_29380_, _29369_, _28339_);
  nor (_29391_, _29380_, _28317_);
  and (_29402_, _29380_, _28317_);
  nor (_29413_, _29402_, _29391_);
  not (_29424_, _28602_);
  nor (_29435_, _29007_, _29424_);
  and (_29446_, _29435_, _28394_);
  and (_29457_, _29358_, _29337_);
  nor (_29468_, _29457_, _29369_);
  and (_29479_, _29468_, _29446_);
  not (_29490_, _29479_);
  nor (_29501_, _29490_, _29413_);
  nor (_29512_, _29380_, _28295_);
  or (_29533_, _29512_, _28306_);
  or (_29534_, _29533_, _29501_);
  and (_29545_, _29534_, _28283_);
  nor (_29556_, _28251_, _28109_);
  nor (_29567_, _29556_, _29304_);
  and (_29578_, _29567_, _29545_);
  and (_29589_, _29315_, _29293_);
  nor (_29600_, _29589_, _29326_);
  and (_29611_, _29600_, _29578_);
  or (_29622_, _29611_, _29326_);
  nor (_29633_, _29622_, _28032_);
  nor (_29644_, _29633_, _29282_);
  and (_29654_, _29633_, _29282_);
  nor (_29665_, _29654_, _29644_);
  and (_29676_, _29665_, _29271_);
  and (_29687_, _18243_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_29698_, _29687_, _27944_);
  nor (_29709_, _21922_, _21379_);
  and (_29720_, _29709_, _21564_);
  and (_29731_, _29720_, _21063_);
  and (_29742_, _29731_, _20704_);
  and (_29753_, _29742_, _20530_);
  and (_29763_, _29753_, _19490_);
  and (_29774_, _29763_, _29007_);
  not (_29785_, _29007_);
  and (_29806_, _19479_, _20519_);
  and (_29807_, _21553_, _21379_);
  and (_29818_, _29807_, _21922_);
  and (_29829_, _29818_, _21052_);
  and (_29840_, _29829_, _20693_);
  and (_29851_, _29840_, _29806_);
  and (_29862_, _29851_, _29785_);
  nor (_29872_, _29862_, _29774_);
  and (_29883_, _29872_, _20323_);
  nor (_29894_, _29872_, _20323_);
  nor (_29905_, _29894_, _29883_);
  and (_29916_, _29905_, _29698_);
  not (_29927_, _20149_);
  nor (_29938_, _29007_, _29927_);
  not (_29949_, _29938_);
  and (_29960_, _29007_, _20323_);
  and (_29971_, _29687_, _18221_);
  not (_29981_, _29971_);
  nor (_29992_, _29981_, _29960_);
  and (_30003_, _29992_, _29949_);
  nor (_30014_, _30003_, _29916_);
  and (_30025_, _29260_, _23615_);
  not (_30036_, _30025_);
  nor (_30047_, _29807_, _21052_);
  and (_30058_, _30047_, _30025_);
  and (_30069_, _30058_, _20704_);
  not (_30080_, _30069_);
  and (_30090_, _30080_, _29806_);
  nor (_30101_, _29806_, _20323_);
  nor (_30112_, _30101_, _30058_);
  and (_30123_, _30112_, _29007_);
  nor (_30134_, _30123_, _30090_);
  and (_30145_, _30134_, _20323_);
  nor (_30156_, _30134_, _20323_);
  nor (_30167_, _30156_, _30145_);
  nor (_30178_, _30167_, _30036_);
  and (_30189_, _29687_, _29260_);
  not (_30199_, _30189_);
  nor (_30210_, _30199_, _29007_);
  not (_30221_, _30210_);
  not (_30232_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_30243_, _18243_, _30232_);
  and (_30254_, _30243_, _29260_);
  not (_30265_, _30254_);
  nor (_30276_, _30265_, _27988_);
  and (_30287_, _30243_, _23593_);
  and (_30298_, _30287_, _27999_);
  nor (_30308_, _30298_, _30276_);
  and (_30319_, _23615_, _18221_);
  and (_30330_, _30319_, _27977_);
  and (_30341_, _27944_, _23615_);
  and (_30352_, _30341_, _20323_);
  nor (_30363_, _30352_, _30330_);
  and (_30374_, _23593_, _18254_);
  not (_30385_, _30374_);
  nor (_30396_, _30385_, _20323_);
  and (_30407_, _29687_, _23593_);
  and (_30427_, _30407_, _21933_);
  and (_30428_, _30243_, _18210_);
  not (_30439_, _30428_);
  nor (_30450_, _30439_, _19479_);
  or (_30461_, _30450_, _30427_);
  nor (_30472_, _30461_, _30396_);
  and (_30483_, _30472_, _30363_);
  and (_30494_, _30483_, _30308_);
  and (_30505_, _30494_, _30221_);
  not (_30516_, _30505_);
  nor (_30526_, _30516_, _30178_);
  and (_30537_, _30526_, _30014_);
  not (_30548_, _30537_);
  nor (_30559_, _30548_, _29676_);
  and (_30570_, _30559_, _29238_);
  not (_30581_, _30570_);
  nor (_30592_, _30581_, _27922_);
  and (_30603_, _30592_, _27911_);
  not (_30614_, _30603_);
  or (_30625_, _30614_, _27889_);
  not (_30635_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_30646_, \oc8051_top_1.oc8051_decoder1.wr , _18199_);
  not (_30657_, _30646_);
  nor (_30668_, _30657_, _26606_);
  and (_30679_, _30668_, _30635_);
  not (_30690_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_30701_, _27889_, _30690_);
  and (_30712_, _30701_, _30679_);
  and (_30723_, _30712_, _30625_);
  nor (_30734_, _30668_, _30690_);
  not (_30744_, _29271_);
  nor (_30755_, _29644_, _27977_);
  nor (_30766_, _30755_, _30744_);
  not (_30777_, _30766_);
  and (_30788_, _20323_, _29927_);
  nor (_30799_, _30788_, _29194_);
  nor (_30810_, _30799_, _27976_);
  nor (_30821_, _30069_, _20530_);
  and (_30832_, _29007_, _19479_);
  and (_30843_, _30832_, _30821_);
  nor (_30853_, _30843_, _29960_);
  nor (_30864_, _29007_, _20323_);
  not (_30875_, _30864_);
  nor (_30886_, _30875_, _30090_);
  nor (_30897_, _30886_, _30036_);
  and (_30908_, _30897_, _30853_);
  or (_30919_, _30908_, _30058_);
  nor (_30930_, _28986_, _28931_);
  not (_30941_, _30287_);
  nor (_30952_, _30941_, _28975_);
  nor (_30962_, _30952_, _30254_);
  nor (_30973_, _30962_, _30930_);
  not (_30984_, _30973_);
  and (_30995_, _28953_, _28931_);
  and (_31006_, _30243_, _27944_);
  and (_31017_, _30319_, _28931_);
  nor (_31028_, _31017_, _31006_);
  nor (_31039_, _31028_, _30995_);
  nand (_31050_, _30407_, _28986_);
  nor (_31061_, _31050_, _28931_);
  nor (_31071_, _30199_, _21922_);
  and (_31082_, _30243_, _18221_);
  not (_31093_, _31082_);
  nor (_31104_, _31093_, _20323_);
  nor (_31115_, _31104_, _31071_);
  not (_31137_, _31115_);
  nor (_31138_, _31137_, _31061_);
  not (_31160_, _31138_);
  nor (_31161_, _31160_, _31039_);
  nor (_31183_, _30385_, _29007_);
  and (_31184_, _30341_, _29007_);
  nor (_31205_, _31184_, _31183_);
  and (_31206_, _31205_, _31161_);
  and (_31217_, _31206_, _30984_);
  not (_31228_, _31217_);
  nor (_31239_, _31228_, _30919_);
  not (_31260_, _31239_);
  nor (_31261_, _31260_, _30810_);
  and (_31282_, _31261_, _30777_);
  not (_31283_, _26781_);
  nor (_31303_, _27023_, _26902_);
  and (_31304_, _31303_, _31283_);
  and (_31325_, _31304_, _27878_);
  nand (_31326_, _31325_, _31282_);
  or (_31347_, _31325_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_31348_, _30668_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_31369_, _31348_, _31347_);
  and (_31370_, _31369_, _31326_);
  or (_31391_, _31370_, _30734_);
  or (_31392_, _31391_, _30723_);
  and (_06662_, _31392_, _42882_);
  and (_31412_, _26054_, _23626_);
  not (_31433_, _31412_);
  and (_31434_, _29007_, _29424_);
  nor (_31455_, _31434_, _29435_);
  nand (_31456_, _29271_, _31455_);
  nor (_31477_, _31093_, _29007_);
  and (_31478_, _30319_, _28580_);
  and (_31499_, _30341_, _21922_);
  nor (_31500_, _31499_, _31478_);
  nor (_31520_, _29981_, _18988_);
  and (_31521_, _29698_, _21922_);
  nor (_31542_, _31521_, _31520_);
  nor (_31543_, _30374_, _30025_);
  nor (_31564_, _31543_, _21922_);
  not (_31565_, _31564_);
  and (_31586_, _31565_, _31542_);
  nand (_31587_, _31586_, _31500_);
  nor (_31608_, _31587_, _31477_);
  and (_31609_, _23350_, _18265_);
  and (_31629_, _31455_, _27955_);
  nor (_31630_, _30941_, _28580_);
  nor (_31651_, _31630_, _30254_);
  or (_31652_, _31651_, _28591_);
  and (_31673_, _29687_, _29249_);
  not (_31674_, _31673_);
  nor (_31695_, _31674_, _21379_);
  and (_31696_, _31006_, _20334_);
  nor (_31717_, _31696_, _31695_);
  nand (_31718_, _31717_, _31652_);
  or (_31738_, _31718_, _31629_);
  nor (_31739_, _31738_, _31609_);
  and (_31760_, _31739_, _31608_);
  and (_31761_, _31760_, _31456_);
  and (_31782_, _31761_, _31433_);
  not (_31783_, _31782_);
  or (_31804_, _31783_, _27889_);
  not (_31805_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_31826_, _27889_, _31805_);
  and (_31827_, _31826_, _30679_);
  and (_31847_, _31827_, _31804_);
  nor (_31848_, _30668_, _31805_);
  not (_31859_, _31282_);
  or (_31870_, _31859_, _27889_);
  and (_31881_, _31826_, _31348_);
  and (_31892_, _31881_, _31870_);
  or (_31903_, _31892_, _31848_);
  or (_31914_, _31903_, _31847_);
  and (_08903_, _31914_, _42882_);
  and (_31935_, _23381_, _18265_);
  not (_31946_, _31935_);
  and (_31956_, _26118_, _23626_);
  nor (_31967_, _29981_, _19975_);
  and (_31978_, _21922_, _21379_);
  nor (_31989_, _31978_, _29709_);
  not (_32000_, _31989_);
  nor (_32011_, _32000_, _29007_);
  and (_32022_, _32000_, _29007_);
  nor (_32033_, _32022_, _32011_);
  and (_32044_, _32033_, _29698_);
  nor (_32054_, _32044_, _31967_);
  nor (_32065_, _30047_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_32076_, _32065_, _21389_);
  nor (_32087_, _32065_, _21389_);
  nor (_32098_, _32087_, _32076_);
  nor (_32109_, _32098_, _30036_);
  not (_32120_, _32109_);
  and (_32131_, _30287_, _28394_);
  nor (_32142_, _30265_, _28383_);
  not (_32153_, _32142_);
  and (_32164_, _30319_, _28372_);
  and (_32174_, _30341_, _21379_);
  nor (_32185_, _32174_, _32164_);
  nand (_32196_, _32185_, _32153_);
  nor (_32207_, _32196_, _32131_);
  nor (_32218_, _30439_, _21922_);
  not (_32229_, _32218_);
  nor (_32240_, _30385_, _21379_);
  nor (_32251_, _31674_, _21553_);
  nor (_32262_, _32251_, _32240_);
  and (_32273_, _32262_, _32229_);
  and (_32283_, _32273_, _32207_);
  and (_32294_, _32283_, _32120_);
  and (_32305_, _32294_, _32054_);
  nor (_32316_, _28580_, _28394_);
  or (_32327_, _32316_, _29347_);
  and (_32338_, _32327_, _29435_);
  nor (_32349_, _32327_, _29435_);
  or (_32360_, _32349_, _32338_);
  and (_32371_, _32360_, _29271_);
  nor (_32382_, _29040_, _29008_);
  nor (_32392_, _32382_, _29051_);
  nor (_32403_, _32392_, _27976_);
  nor (_32414_, _32403_, _32371_);
  and (_32425_, _32414_, _32305_);
  not (_32436_, _32425_);
  nor (_32447_, _32436_, _31956_);
  and (_32458_, _32447_, _31946_);
  not (_32469_, _32458_);
  or (_32480_, _32469_, _27889_);
  not (_32491_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_32501_, _27889_, _32491_);
  and (_32512_, _32501_, _30679_);
  and (_32523_, _32512_, _32480_);
  nor (_32534_, _30668_, _32491_);
  not (_32545_, _27023_);
  and (_32556_, _32545_, _26902_);
  and (_32567_, _32556_, _26781_);
  and (_32578_, _32567_, _27878_);
  nand (_32589_, _32578_, _31282_);
  or (_32600_, _32578_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_32610_, _32600_, _31348_);
  and (_32621_, _32610_, _32589_);
  or (_32632_, _32621_, _32534_);
  or (_32643_, _32632_, _32523_);
  and (_08914_, _32643_, _42882_);
  and (_32664_, _23413_, _18265_);
  not (_32675_, _32664_);
  and (_32686_, _26183_, _23626_);
  nor (_32697_, _29981_, _18669_);
  nor (_32708_, _31978_, _29007_);
  nor (_32718_, _29709_, _29785_);
  nor (_32729_, _32718_, _32708_);
  nor (_32740_, _32729_, _21564_);
  and (_32751_, _32729_, _21564_);
  nor (_32762_, _32751_, _32740_);
  and (_32773_, _32762_, _29698_);
  nor (_32784_, _32773_, _32697_);
  nor (_32795_, _29051_, _28569_);
  nor (_32806_, _32795_, _29062_);
  nor (_32817_, _32806_, _27976_);
  and (_32827_, _30287_, _28361_);
  not (_32838_, _32827_);
  nor (_32849_, _30265_, _28350_);
  not (_32860_, _32849_);
  and (_32871_, _30319_, _28339_);
  and (_32882_, _30341_, _21553_);
  nor (_32893_, _32882_, _32871_);
  and (_32904_, _32893_, _32860_);
  and (_32915_, _32904_, _32838_);
  nor (_32926_, _30439_, _21379_);
  not (_32936_, _32926_);
  nor (_32947_, _30385_, _21553_);
  nor (_32958_, _31674_, _21052_);
  nor (_32969_, _32958_, _32947_);
  and (_32980_, _32969_, _32936_);
  and (_32991_, _32980_, _32915_);
  not (_33002_, _32991_);
  nor (_33013_, _33002_, _32817_);
  nor (_33024_, _29468_, _29446_);
  nor (_33035_, _33024_, _30744_);
  and (_33045_, _33035_, _29490_);
  nor (_33056_, _32087_, _21553_);
  and (_33067_, _29807_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_33078_, _33067_, _33056_);
  nor (_33089_, _33078_, _30036_);
  nor (_33100_, _33089_, _33045_);
  and (_33111_, _33100_, _33013_);
  and (_33122_, _33111_, _32784_);
  not (_33133_, _33122_);
  nor (_33144_, _33133_, _32686_);
  and (_33154_, _33144_, _32675_);
  not (_33165_, _33154_);
  or (_33176_, _33165_, _27889_);
  not (_33187_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_33198_, _27889_, _33187_);
  and (_33209_, _33198_, _30679_);
  and (_33220_, _33209_, _33176_);
  nor (_33231_, _30668_, _33187_);
  nand (_33242_, _27878_, _26781_);
  or (_33253_, _31303_, _33242_);
  and (_33263_, _33253_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_33274_, _26902_);
  and (_33285_, _26781_, _27023_);
  and (_33296_, _33285_, _33274_);
  not (_33307_, _33296_);
  nor (_33318_, _33307_, _31282_);
  and (_33329_, _26781_, _26902_);
  and (_33340_, _33329_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_33351_, _33340_, _33318_);
  and (_33362_, _33351_, _27878_);
  or (_33372_, _33362_, _33263_);
  and (_33383_, _33372_, _31348_);
  or (_33394_, _33383_, _33231_);
  or (_33405_, _33394_, _33220_);
  and (_08925_, _33405_, _42882_);
  and (_33426_, _26248_, _23626_);
  not (_33437_, _33426_);
  and (_33448_, _23466_, _18265_);
  and (_33459_, _29490_, _29413_);
  or (_33470_, _33459_, _30744_);
  nor (_33480_, _33470_, _29501_);
  not (_33491_, _33480_);
  nor (_33502_, _29062_, _28536_);
  nor (_33513_, _33502_, _29073_);
  nor (_33524_, _33513_, _27976_);
  nor (_33535_, _29981_, _19653_);
  and (_33546_, _29720_, _29007_);
  and (_33557_, _29818_, _29785_);
  nor (_33568_, _33557_, _33546_);
  nor (_33579_, _33568_, _21052_);
  not (_33589_, _29698_);
  and (_33600_, _33568_, _21052_);
  or (_33611_, _33600_, _33589_);
  nor (_33622_, _33611_, _33579_);
  nor (_33633_, _33622_, _33535_);
  not (_33644_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_33655_, _29807_, _33644_);
  nor (_33666_, _33655_, _21063_);
  nor (_33677_, _30385_, _21052_);
  nor (_33688_, _30047_, _30036_);
  nor (_33698_, _33688_, _33677_);
  or (_33709_, _33698_, _33666_);
  nor (_33720_, _30265_, _28295_);
  and (_33731_, _30287_, _28317_);
  nor (_33742_, _33731_, _33720_);
  and (_33753_, _30319_, _28306_);
  and (_33764_, _30341_, _21052_);
  nor (_33775_, _33764_, _33753_);
  nor (_33786_, _31674_, _20693_);
  nor (_33797_, _30439_, _21553_);
  nor (_33807_, _33797_, _33786_);
  and (_33818_, _33807_, _33775_);
  and (_33829_, _33818_, _33742_);
  and (_33840_, _33829_, _33709_);
  nand (_33851_, _33840_, _33633_);
  nor (_33862_, _33851_, _33524_);
  and (_33873_, _33862_, _33491_);
  not (_33884_, _33873_);
  nor (_33895_, _33884_, _33448_);
  and (_33906_, _33895_, _33437_);
  not (_33916_, _33906_);
  or (_33927_, _33916_, _27889_);
  not (_33938_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_33949_, _27889_, _33938_);
  and (_33960_, _33949_, _30679_);
  and (_33971_, _33960_, _33927_);
  nor (_33982_, _30668_, _33938_);
  and (_33993_, _33242_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_34004_, _31303_, _26781_);
  and (_34015_, _34004_, _31859_);
  or (_34026_, _31303_, _31283_);
  nor (_34036_, _34026_, _33938_);
  or (_34047_, _34036_, _34015_);
  and (_34058_, _34047_, _27878_);
  or (_34069_, _34058_, _33993_);
  and (_34080_, _34069_, _31348_);
  or (_34091_, _34080_, _33982_);
  or (_34102_, _34091_, _33971_);
  and (_08936_, _34102_, _42882_);
  and (_34123_, _26313_, _23626_);
  not (_34134_, _34123_);
  and (_34144_, _23487_, _18265_);
  nor (_34155_, _29534_, _28283_);
  not (_34166_, _34155_);
  nor (_34177_, _30744_, _29545_);
  and (_34188_, _34177_, _34166_);
  not (_34199_, _34188_);
  nor (_34210_, _29139_, _28283_);
  and (_34221_, _29139_, _28283_);
  nor (_34232_, _34221_, _34210_);
  and (_34243_, _34232_, _27955_);
  and (_34253_, _29731_, _29007_);
  and (_34264_, _29829_, _29785_);
  nor (_34277_, _34264_, _34253_);
  and (_34296_, _34277_, _20693_);
  nor (_34307_, _34277_, _20693_);
  nor (_34318_, _34307_, _34296_);
  and (_34329_, _34318_, _29698_);
  nor (_34340_, _29007_, _18834_);
  and (_34351_, _29007_, _20704_);
  nor (_34361_, _34351_, _34340_);
  nor (_34372_, _34361_, _29981_);
  and (_34383_, _30319_, _28251_);
  and (_34394_, _30341_, _20693_);
  nor (_34405_, _34394_, _34383_);
  and (_34416_, _30287_, _28283_);
  nor (_34427_, _30265_, _28262_);
  or (_34438_, _34427_, _34416_);
  not (_34449_, _34438_);
  and (_34460_, _34449_, _34405_);
  not (_34470_, _34460_);
  or (_34481_, _34470_, _34372_);
  nor (_34492_, _34481_, _34329_);
  nor (_34503_, _30058_, _20704_);
  nor (_34514_, _30385_, _20693_);
  nor (_34525_, _30069_, _30036_);
  nor (_34536_, _34525_, _34514_);
  or (_34547_, _34536_, _34503_);
  nor (_34558_, _31674_, _20519_);
  nor (_34569_, _30439_, _21052_);
  nor (_34580_, _34569_, _34558_);
  and (_34590_, _34580_, _34547_);
  and (_34601_, _34590_, _34492_);
  not (_34612_, _34601_);
  nor (_34623_, _34612_, _34243_);
  and (_34634_, _34623_, _34199_);
  not (_34645_, _34634_);
  nor (_34656_, _34645_, _34144_);
  and (_34667_, _34656_, _34134_);
  not (_34678_, _34667_);
  or (_34689_, _34678_, _27889_);
  not (_34699_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_34710_, _27889_, _34699_);
  and (_34721_, _34710_, _30679_);
  and (_34732_, _34721_, _34689_);
  nor (_34743_, _30668_, _34699_);
  not (_34754_, _27878_);
  and (_34765_, _27034_, _31283_);
  nor (_34776_, _27034_, _31283_);
  nor (_34787_, _34776_, _34765_);
  or (_34798_, _34787_, _34754_);
  and (_34808_, _34798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_34819_, _34765_, _31859_);
  and (_34830_, _34776_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_34841_, _34830_, _34819_);
  and (_34852_, _34841_, _27878_);
  or (_34863_, _34852_, _34808_);
  and (_34874_, _34863_, _31348_);
  or (_34885_, _34874_, _34743_);
  or (_34896_, _34885_, _34732_);
  and (_08947_, _34896_, _42882_);
  and (_34916_, _23530_, _18265_);
  not (_34927_, _34916_);
  and (_34938_, _26400_, _23626_);
  nor (_34949_, _29150_, _28240_);
  nor (_34960_, _34949_, _29161_);
  nor (_34971_, _34960_, _27976_);
  not (_34982_, _34971_);
  nor (_34993_, _30265_, _28098_);
  and (_35004_, _30287_, _28109_);
  nor (_35015_, _35004_, _34993_);
  and (_35025_, _30319_, _28087_);
  and (_35036_, _30341_, _20519_);
  nor (_35047_, _35036_, _35025_);
  nor (_35058_, _31674_, _19479_);
  not (_35069_, _35058_);
  nor (_35080_, _30385_, _20519_);
  nor (_35091_, _30439_, _20693_);
  nor (_35101_, _35091_, _35080_);
  and (_35112_, _35101_, _35069_);
  and (_35123_, _35112_, _35047_);
  and (_35134_, _35123_, _35015_);
  nor (_35145_, _29567_, _29545_);
  not (_35156_, _35145_);
  nor (_35167_, _30744_, _29578_);
  and (_35178_, _35167_, _35156_);
  nor (_35189_, _29007_, _19805_);
  and (_35200_, _29007_, _20530_);
  nor (_35211_, _35200_, _35189_);
  nor (_35221_, _35211_, _29981_);
  and (_35232_, _29742_, _29007_);
  and (_35243_, _29840_, _29785_);
  nor (_35254_, _35243_, _35232_);
  and (_35265_, _35254_, _20519_);
  nor (_35276_, _35254_, _20519_);
  or (_35287_, _35276_, _33589_);
  nor (_35298_, _35287_, _35265_);
  nor (_35309_, _35298_, _35221_);
  not (_35320_, _30123_);
  and (_35331_, _35320_, _30821_);
  nor (_35341_, _30123_, _30069_);
  nor (_35352_, _35341_, _20519_);
  nor (_35363_, _35352_, _35331_);
  nor (_35374_, _35363_, _30036_);
  not (_35385_, _35374_);
  nand (_35396_, _35385_, _35309_);
  nor (_35407_, _35396_, _35178_);
  and (_35418_, _35407_, _35134_);
  and (_35429_, _35418_, _34982_);
  not (_35440_, _35429_);
  nor (_35451_, _35440_, _34938_);
  and (_35461_, _35451_, _34927_);
  not (_35472_, _35461_);
  or (_35483_, _35472_, _27889_);
  not (_35494_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_35505_, _27889_, _35494_);
  and (_35516_, _35505_, _30679_);
  and (_35527_, _35516_, _35483_);
  nor (_35538_, _30668_, _35494_);
  and (_35549_, _32556_, _31283_);
  and (_35560_, _35549_, _27878_);
  nand (_35571_, _35560_, _31282_);
  or (_35582_, _35560_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_35592_, _35582_, _31348_);
  and (_35603_, _35592_, _35571_);
  or (_35614_, _35603_, _35538_);
  or (_35625_, _35614_, _35527_);
  and (_08958_, _35625_, _42882_);
  and (_35646_, _26464_, _23626_);
  not (_35657_, _35646_);
  and (_35668_, _23562_, _18265_);
  nor (_35679_, _29600_, _29578_);
  not (_35690_, _35679_);
  nor (_35701_, _30744_, _29611_);
  and (_35712_, _35701_, _35690_);
  not (_35722_, _35712_);
  nor (_35733_, _29161_, _28207_);
  nor (_35744_, _35733_, _29172_);
  nor (_35755_, _35744_, _27976_);
  nor (_35766_, _29007_, _28010_);
  or (_35777_, _35766_, _29981_);
  nor (_35788_, _35777_, _30832_);
  or (_35799_, _29007_, _20519_);
  or (_35810_, _35243_, _29753_);
  and (_35821_, _35810_, _35799_);
  and (_35832_, _35821_, _19490_);
  nor (_35842_, _35821_, _19490_);
  or (_35853_, _35842_, _33589_);
  nor (_35864_, _35853_, _35832_);
  nor (_35875_, _35864_, _35788_);
  nor (_35886_, _35331_, _19479_);
  and (_35897_, _35331_, _19479_);
  nor (_35908_, _35897_, _35886_);
  nor (_35919_, _35908_, _30036_);
  and (_35929_, _30287_, _28054_);
  nor (_35940_, _30265_, _28043_);
  not (_35951_, _35940_);
  and (_35962_, _30319_, _28032_);
  and (_35973_, _30341_, _19479_);
  nor (_35984_, _35973_, _35962_);
  nand (_35995_, _35984_, _35951_);
  nor (_36006_, _35995_, _35929_);
  nor (_36016_, _30439_, _20519_);
  not (_36027_, _36016_);
  nor (_36038_, _30385_, _19479_);
  nor (_36049_, _31674_, _20323_);
  nor (_36060_, _36049_, _36038_);
  and (_36071_, _36060_, _36027_);
  and (_36082_, _36071_, _36006_);
  not (_36092_, _36082_);
  nor (_36103_, _36092_, _35919_);
  and (_36114_, _36103_, _35875_);
  not (_36125_, _36114_);
  nor (_36136_, _36125_, _35755_);
  and (_36147_, _36136_, _35722_);
  not (_36158_, _36147_);
  nor (_36169_, _36158_, _35668_);
  and (_36179_, _36169_, _35657_);
  not (_36190_, _36179_);
  or (_36201_, _36190_, _27889_);
  not (_36212_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_36223_, _27889_, _36212_);
  and (_36234_, _36223_, _30679_);
  and (_36245_, _36234_, _36201_);
  nor (_36256_, _30668_, _36212_);
  nor (_36266_, _26781_, _26902_);
  and (_36277_, _36266_, _27023_);
  and (_36288_, _36277_, _27878_);
  nand (_36299_, _36288_, _31282_);
  or (_36310_, _36288_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_36321_, _36310_, _31348_);
  and (_36332_, _36321_, _36299_);
  or (_36343_, _36332_, _36256_);
  or (_36353_, _36343_, _36245_);
  and (_08969_, _36353_, _42882_);
  and (_36374_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36385_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_36396_, _36385_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_36407_, _36396_);
  not (_36418_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_36428_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_36439_, _36428_, _36418_);
  and (_36450_, _36385_, _18199_);
  and (_36461_, _36450_, _36439_);
  not (_36472_, _36461_);
  not (_36483_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_36494_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_36505_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_36516_, _36505_, _36494_);
  and (_36527_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_36537_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_36548_, _36537_, _36494_);
  and (_36559_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  not (_36570_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_36581_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _36570_);
  and (_36592_, _36581_, _36494_);
  and (_36603_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_36614_, _36603_, _36559_);
  or (_36625_, _36614_, _36527_);
  and (_36636_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_36646_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_36657_, _36646_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_36668_, _36657_, _36494_);
  and (_36679_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_36690_, _36679_, _36636_);
  nor (_36701_, _36505_, _36494_);
  and (_36712_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_36723_, _36505_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_36734_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_36745_, _36734_, _36712_);
  or (_36756_, _36745_, _36690_);
  nor (_36767_, _36756_, _36625_);
  and (_36778_, _36767_, _36483_);
  nor (_36789_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _36483_);
  nor (_36800_, _36789_, _36778_);
  nor (_36811_, _36800_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_36822_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_36833_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _36822_);
  nor (_36844_, _36833_, _36811_);
  nor (_36855_, _36844_, _36472_);
  not (_36866_, _36855_);
  not (_36877_, _36439_);
  nor (_36888_, _36450_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_36898_, _36888_, _36877_);
  and (_36909_, _36898_, _36866_);
  not (_36920_, _36909_);
  and (_36931_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_36942_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_36953_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_36964_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_36975_, _36964_, _36953_);
  and (_36986_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_36997_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_37007_, _36997_, _36986_);
  and (_37018_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_37029_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_37040_, _37029_, _37018_);
  and (_37051_, _37040_, _37007_);
  and (_37062_, _37051_, _36975_);
  or (_37073_, _36636_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_37084_, _37073_, _37062_);
  nor (_37095_, _37084_, _36942_);
  nor (_37106_, _37095_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37117_, _37106_, _36931_);
  and (_37127_, _37117_, _36461_);
  not (_37138_, _37127_);
  nor (_37149_, _36450_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_37160_, _37149_, _36877_);
  and (_37171_, _37160_, _37138_);
  and (_37182_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37193_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37204_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_37215_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_37226_, _37215_, _37204_);
  and (_37236_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_37247_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_37258_, _37247_, _37236_);
  and (_37269_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_37280_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_37291_, _37280_, _37269_);
  and (_37302_, _37291_, _37258_);
  and (_37313_, _37302_, _37226_);
  nor (_37324_, _37313_, _37073_);
  or (_37335_, _37324_, _37193_);
  and (_37346_, _37335_, _36822_);
  nor (_37357_, _37346_, _37182_);
  and (_37368_, _37357_, _36461_);
  not (_37379_, _37368_);
  nor (_37390_, _36450_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_37401_, _37390_, _36877_);
  and (_37410_, _37401_, _37379_);
  not (_37421_, _37410_);
  and (_37432_, _37421_, _37171_);
  and (_37443_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37454_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37465_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_37476_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_37487_, _37476_, _37465_);
  and (_37498_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_37509_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_37520_, _37509_, _37498_);
  and (_37531_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_37542_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_37553_, _37542_, _37531_);
  and (_37564_, _37553_, _37520_);
  and (_37575_, _37564_, _37487_);
  nor (_37586_, _37575_, _36636_);
  and (_37597_, _37586_, _36483_);
  or (_37608_, _37597_, _37454_);
  and (_37619_, _37608_, _36822_);
  nor (_37630_, _37619_, _37443_);
  and (_37641_, _37630_, _36461_);
  not (_37652_, _37641_);
  nor (_37663_, _36450_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_37674_, _37663_, _36877_);
  and (_37685_, _37674_, _37652_);
  and (_37696_, _37685_, _37432_);
  and (_37707_, _37696_, _36920_);
  and (_37718_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37729_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37740_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_37751_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_37762_, _37751_, _37740_);
  and (_37773_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_37784_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_37795_, _37784_, _37773_);
  and (_37806_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_37817_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_37828_, _37817_, _37806_);
  and (_37839_, _37828_, _37795_);
  and (_37850_, _37839_, _37762_);
  nor (_37861_, _37850_, _36636_);
  and (_37872_, _37861_, _36483_);
  or (_37883_, _37872_, _37729_);
  and (_37894_, _37883_, _36822_);
  nor (_37905_, _37894_, _37718_);
  and (_37916_, _37905_, _36461_);
  not (_37927_, _37916_);
  nor (_37938_, _36450_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_37949_, _37938_, _36877_);
  and (_37960_, _37949_, _37927_);
  and (_37971_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37982_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37993_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_38004_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_38015_, _38004_, _37993_);
  and (_38026_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_38037_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_38048_, _38037_, _38026_);
  and (_38059_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_38069_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_38080_, _38069_, _38059_);
  and (_38091_, _38080_, _38048_);
  and (_38101_, _38091_, _38015_);
  nor (_38112_, _38101_, _37073_);
  nor (_38123_, _38112_, _37982_);
  nor (_38134_, _38123_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_38145_, _38134_, _37971_);
  nor (_38156_, _38145_, _36472_);
  and (_38165_, _36472_, \oc8051_top_1.oc8051_decoder1.op [2]);
  or (_38166_, _38165_, _38156_);
  and (_38167_, _38166_, _36439_);
  and (_38168_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_38169_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_38170_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_38171_, _38170_, _38169_);
  or (_38172_, _38171_, _38168_);
  and (_38173_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_38174_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_38175_, _38174_, _38173_);
  and (_38176_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_38177_, _38176_, _36636_);
  nand (_38178_, _38177_, _38175_);
  nor (_38179_, _38178_, _38172_);
  and (_38180_, _38179_, _36483_);
  nor (_38181_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _36483_);
  nor (_38182_, _38181_, _38180_);
  nor (_38183_, _38182_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_38184_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _36822_);
  nor (_38185_, _38184_, _38183_);
  nor (_38186_, _38185_, _36472_);
  not (_38187_, _38186_);
  nor (_38188_, _36450_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_38189_, _38188_, _36877_);
  and (_38190_, _38189_, _38187_);
  not (_38191_, _38190_);
  nor (_38192_, _38191_, _38167_);
  and (_38193_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_38194_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_38195_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_38196_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_38197_, _38196_, _38195_);
  and (_38198_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_38199_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_38200_, _38199_, _38198_);
  and (_38201_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_38202_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_38203_, _38202_, _38201_);
  and (_38204_, _38203_, _38200_);
  and (_38205_, _38204_, _38197_);
  nor (_38206_, _38205_, _36636_);
  and (_38207_, _38206_, _36483_);
  or (_38208_, _38207_, _38194_);
  and (_38209_, _38208_, _36822_);
  nor (_38210_, _38209_, _38193_);
  and (_38211_, _38210_, _36461_);
  not (_38212_, _38211_);
  nor (_38213_, _36450_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_38214_, _38213_, _36877_);
  and (_38215_, _38214_, _38212_);
  not (_38216_, _38215_);
  and (_38217_, _38216_, _38192_);
  and (_38218_, _38217_, _37960_);
  and (_38219_, _38218_, _37707_);
  not (_38220_, _37171_);
  and (_38221_, _37685_, _37410_);
  and (_38222_, _38221_, _38220_);
  and (_38223_, _38222_, _36909_);
  and (_38224_, _38218_, _38223_);
  nor (_38225_, _37685_, _37410_);
  and (_38226_, _38225_, _37171_);
  and (_38227_, _38226_, _36909_);
  and (_38228_, _38218_, _38227_);
  nor (_38229_, _38228_, _38224_);
  not (_38230_, _38229_);
  nor (_38231_, _38230_, _38219_);
  and (_38232_, _38226_, _36920_);
  and (_38233_, _38216_, _38167_);
  nor (_38234_, _37960_, _38190_);
  and (_38235_, _38234_, _38233_);
  and (_38236_, _38235_, _38232_);
  and (_38237_, _38235_, _37707_);
  nor (_38238_, _38237_, _38236_);
  and (_38239_, _38238_, _38231_);
  nor (_38240_, _38239_, _36407_);
  not (_38241_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_38242_, _18199_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_38243_, _38242_, _38241_);
  and (_38244_, _37410_, _38220_);
  nor (_38245_, _38215_, _38167_);
  and (_38246_, _38234_, _38245_);
  and (_38247_, _38246_, _38244_);
  and (_38248_, _38247_, _38243_);
  and (_38249_, _38237_, _18199_);
  and (_38250_, _38236_, _18199_);
  nor (_38251_, _38250_, _38249_);
  nor (_38252_, _38251_, _36385_);
  nor (_38253_, _38252_, _38248_);
  not (_38254_, _38253_);
  nor (_38255_, _38254_, _38240_);
  nor (_38256_, _38255_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38257_, _38256_, _36374_);
  and (_38258_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38259_, _37960_, _38215_);
  and (_38260_, _38259_, _38192_);
  and (_38261_, _38260_, _37707_);
  not (_38262_, _37960_);
  nor (_38263_, _37685_, _37421_);
  and (_38264_, _38263_, _37171_);
  and (_38265_, _38264_, _36909_);
  and (_38266_, _38265_, _38217_);
  and (_38267_, _38266_, _38262_);
  nor (_38268_, _38267_, _38261_);
  and (_38269_, _38190_, _38167_);
  nor (_38270_, _38215_, _36909_);
  and (_38271_, _38270_, _38269_);
  and (_38272_, _38271_, _37696_);
  and (_38273_, _38227_, _38260_);
  and (_38274_, _37960_, _38191_);
  and (_38275_, _38274_, _38233_);
  and (_38276_, _38275_, _38232_);
  nor (_38277_, _38276_, _38273_);
  not (_38278_, _38277_);
  nor (_38279_, _38278_, _38272_);
  and (_38280_, _38221_, _37171_);
  and (_38281_, _38280_, _36920_);
  and (_38282_, _38281_, _38275_);
  and (_38283_, _37432_, _36909_);
  and (_38284_, _38283_, _38275_);
  nor (_38285_, _38284_, _38282_);
  and (_38286_, _38285_, _38279_);
  and (_38287_, _38222_, _36920_);
  and (_38288_, _38287_, _38275_);
  and (_38289_, _38264_, _36920_);
  and (_38290_, _38289_, _38275_);
  nor (_38291_, _38290_, _38288_);
  and (_38292_, _38215_, _37707_);
  not (_38293_, _38292_);
  nor (_38294_, _37410_, _37171_);
  and (_38295_, _38294_, _37685_);
  and (_38296_, _38295_, _38260_);
  not (_38297_, _37685_);
  and (_38298_, _38294_, _38297_);
  and (_38299_, _38298_, _36920_);
  and (_38300_, _38299_, _38275_);
  nor (_38301_, _38300_, _38296_);
  and (_38302_, _38301_, _38293_);
  and (_38303_, _38302_, _38291_);
  and (_38304_, _38303_, _38286_);
  and (_38305_, _38304_, _38268_);
  and (_38306_, _38275_, _38265_);
  and (_38307_, _38298_, _36909_);
  and (_38308_, _38307_, _38275_);
  nor (_38309_, _38308_, _38306_);
  and (_38310_, _38246_, _37696_);
  and (_38311_, _38244_, _38297_);
  and (_38312_, _38311_, _36920_);
  and (_38313_, _38312_, _38275_);
  nor (_38314_, _38313_, _38310_);
  and (_38315_, _38314_, _38309_);
  and (_38316_, _38289_, _38260_);
  and (_38317_, _37696_, _36909_);
  and (_38318_, _38317_, _38260_);
  nor (_38319_, _38318_, _38316_);
  and (_38320_, _38223_, _38260_);
  and (_38321_, _38312_, _38217_);
  nor (_38322_, _38321_, _38320_);
  and (_38323_, _38322_, _38319_);
  and (_38324_, _38323_, _38315_);
  and (_38325_, _38232_, _38260_);
  and (_38326_, _38311_, _36909_);
  and (_38327_, _38326_, _38217_);
  nor (_38328_, _38327_, _38325_);
  not (_38329_, _38328_);
  nor (_38330_, _38326_, _38295_);
  not (_38331_, _38330_);
  and (_38332_, _38331_, _38275_);
  nor (_38333_, _38332_, _38329_);
  and (_38334_, _38295_, _36909_);
  and (_38335_, _38334_, _38246_);
  not (_38336_, _38335_);
  and (_38337_, _38295_, _36920_);
  and (_38338_, _38337_, _38246_);
  and (_38339_, _38246_, _38307_);
  nor (_38340_, _38339_, _38338_);
  and (_38341_, _38340_, _38336_);
  and (_38342_, _38246_, _38264_);
  and (_38343_, _38287_, _38217_);
  nor (_38344_, _38343_, _38342_);
  and (_38345_, _38344_, _38341_);
  and (_38346_, _38345_, _38333_);
  and (_38347_, _38346_, _38324_);
  and (_38348_, _38347_, _38305_);
  nor (_38349_, _38348_, _36407_);
  and (_38350_, \oc8051_top_1.oc8051_decoder1.state [0], _18199_);
  and (_38351_, _38350_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_38352_, _38351_, _38296_);
  nor (_38353_, _38352_, _38248_);
  not (_38354_, _38353_);
  nor (_38355_, _38354_, _38349_);
  nor (_38356_, _38355_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38357_, _38356_, _38258_);
  and (_38358_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_38359_, _38269_, _38216_);
  and (_38360_, _38359_, _38264_);
  nor (_38361_, _38215_, _36920_);
  and (_38362_, _38361_, _38269_);
  and (_38363_, _38362_, _38226_);
  nor (_38364_, _38363_, _38360_);
  and (_38365_, _38362_, _37696_);
  and (_38366_, _38298_, _38359_);
  nor (_38367_, _38366_, _38365_);
  not (_38368_, _38367_);
  and (_38369_, _38362_, _38311_);
  and (_38370_, _38295_, _38359_);
  or (_38371_, _38370_, _38369_);
  nor (_38372_, _38371_, _38368_);
  and (_38373_, _38372_, _38364_);
  and (_38374_, _37960_, _38216_);
  and (_38375_, _38374_, _38192_);
  and (_38376_, _38375_, _37707_);
  or (_38377_, _38223_, _38227_);
  and (_38378_, _38377_, _38375_);
  nor (_38379_, _38378_, _38376_);
  and (_38380_, _38246_, _38265_);
  and (_38381_, _38226_, _38271_);
  nor (_38382_, _38381_, _38380_);
  and (_38383_, _38311_, _38271_);
  and (_38384_, _38280_, _38271_);
  nor (_38385_, _38384_, _38383_);
  and (_38386_, _38222_, _38271_);
  nor (_38387_, _38386_, _38296_);
  and (_38388_, _38387_, _38385_);
  and (_38389_, _38388_, _38382_);
  and (_38390_, _38389_, _38379_);
  and (_38391_, _38390_, _38373_);
  nor (_38392_, _38391_, _36407_);
  and (_38393_, _38243_, _38222_);
  and (_38394_, _38393_, _38246_);
  or (_38395_, _38394_, _38352_);
  nor (_38396_, _38395_, _38392_);
  nor (_38397_, _38396_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38398_, _38397_, _38358_);
  nor (_38399_, _38398_, _38357_);
  and (_38400_, _38399_, _38257_);
  and (_09519_, _38400_, _42882_);
  and (_38401_, _30679_, _27703_);
  and (_38402_, _38401_, _26781_);
  and (_38403_, _27845_, _27374_);
  and (_38404_, _27242_, _27560_);
  and (_38405_, _38404_, _38403_);
  and (_38406_, _38405_, _32556_);
  and (_38407_, _38406_, _38402_);
  nor (_38408_, _38407_, _27396_);
  not (_38409_, _38407_);
  and (_38410_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_38411_, _23626_, _18265_);
  and (_38412_, _29260_, _23604_);
  nor (_38413_, _30374_, _38412_);
  and (_38414_, _38413_, _38411_);
  nor (_38415_, _30428_, _31673_);
  and (_38416_, _38415_, _38414_);
  nor (_38417_, _38416_, _19479_);
  not (_38418_, _38417_);
  and (_38419_, _38418_, _36006_);
  and (_38420_, _38419_, _35875_);
  nor (_38421_, _38420_, _38409_);
  nor (_38422_, _38421_, _38410_);
  and (_38423_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_38424_, _38416_, _20519_);
  not (_38425_, _38424_);
  and (_38426_, _38425_, _35047_);
  and (_38427_, _38426_, _35015_);
  and (_38428_, _38427_, _35309_);
  nor (_38429_, _38428_, _38409_);
  nor (_38430_, _38429_, _38423_);
  and (_38431_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_38432_, _38416_, _20693_);
  not (_38433_, _38432_);
  and (_38434_, _38433_, _34492_);
  nor (_38435_, _38434_, _38409_);
  nor (_38436_, _38435_, _38431_);
  and (_38437_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_38438_, _38416_, _21052_);
  not (_38439_, _38438_);
  and (_38440_, _38439_, _33775_);
  and (_38441_, _38440_, _33742_);
  and (_38442_, _38441_, _33633_);
  nor (_38443_, _38442_, _38409_);
  nor (_38444_, _38443_, _38437_);
  and (_38445_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_38446_, _38416_, _21553_);
  not (_38447_, _38446_);
  and (_38448_, _38447_, _32915_);
  and (_38449_, _38448_, _32784_);
  nor (_38450_, _38449_, _38409_);
  nor (_38451_, _38450_, _38445_);
  and (_38452_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_38453_, _38416_, _21379_);
  not (_38454_, _38453_);
  and (_38455_, _38454_, _32207_);
  and (_38456_, _38455_, _32054_);
  nor (_38457_, _38456_, _38409_);
  nor (_38458_, _38457_, _38452_);
  nor (_38459_, _38407_, _26968_);
  nor (_38460_, _38416_, _21922_);
  not (_38461_, _38460_);
  and (_38462_, _38461_, _31542_);
  and (_38463_, _38462_, _31500_);
  and (_38464_, _38463_, _31652_);
  not (_38465_, _38464_);
  and (_38466_, _38465_, _38407_);
  nor (_38467_, _38466_, _38459_);
  and (_38468_, _38467_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38469_, _38468_, _38458_);
  and (_38470_, _38469_, _38451_);
  and (_38471_, _38470_, _38444_);
  and (_38472_, _38471_, _38436_);
  and (_38473_, _38472_, _38430_);
  and (_38474_, _38473_, _38422_);
  and (_38475_, _38474_, _38408_);
  nor (_38476_, _38474_, _38408_);
  nor (_38477_, _38476_, _38475_);
  and (_38478_, _38477_, _27111_);
  nor (_38479_, _38407_, _27440_);
  not (_38480_, _38479_);
  nor (_38481_, _38480_, _38478_);
  or (_38482_, _38416_, _20323_);
  and (_38483_, _38482_, _30363_);
  and (_38484_, _38483_, _30308_);
  and (_38485_, _38484_, _30014_);
  and (_38486_, _38485_, _38407_);
  or (_38487_, _38486_, _38481_);
  nor (_09540_, _38487_, rst);
  not (_38488_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38489_, _38467_, _38488_);
  nor (_38490_, _38467_, _38488_);
  nor (_38491_, _38490_, _38489_);
  and (_38492_, _38491_, _27111_);
  nor (_38493_, _38492_, _26979_);
  nor (_38494_, _38493_, _38407_);
  nor (_38495_, _38494_, _38466_);
  nand (_10696_, _38495_, _42882_);
  nor (_38496_, _38468_, _38458_);
  nor (_38497_, _38496_, _38469_);
  nor (_38498_, _38497_, _26528_);
  nor (_38499_, _38498_, _26825_);
  nor (_38500_, _38499_, _38407_);
  nor (_38501_, _38500_, _38457_);
  nand (_10707_, _38501_, _42882_);
  nor (_38502_, _38469_, _38451_);
  nor (_38503_, _38502_, _38470_);
  nor (_38504_, _38503_, _26528_);
  nor (_38505_, _38504_, _26573_);
  nor (_38506_, _38505_, _38407_);
  nor (_38507_, _38506_, _38450_);
  nand (_10718_, _38507_, _42882_);
  nor (_38508_, _38470_, _38444_);
  nor (_38509_, _38508_, _38471_);
  nor (_38510_, _38509_, _26528_);
  nor (_38511_, _38510_, _27637_);
  nor (_38512_, _38511_, _38407_);
  nor (_38513_, _38512_, _38443_);
  nor (_10729_, _38513_, rst);
  nor (_38514_, _38471_, _38436_);
  nor (_38515_, _38514_, _38472_);
  nor (_38516_, _38515_, _26528_);
  nor (_38517_, _38516_, _27769_);
  nor (_38518_, _38517_, _38407_);
  nor (_38519_, _38518_, _38435_);
  nor (_10740_, _38519_, rst);
  nor (_38520_, _38472_, _38430_);
  nor (_38521_, _38520_, _38473_);
  nor (_38522_, _38521_, _26528_);
  nor (_38523_, _38522_, _27286_);
  nor (_38524_, _38523_, _38407_);
  nor (_38525_, _38524_, _38429_);
  nor (_10751_, _38525_, rst);
  nor (_38526_, _38473_, _38422_);
  nor (_38527_, _38526_, _38474_);
  nor (_38528_, _38527_, _26528_);
  nor (_38529_, _38528_, _27143_);
  nor (_38530_, _38529_, _38407_);
  nor (_38531_, _38530_, _38421_);
  nor (_10762_, _38531_, rst);
  and (_38532_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18199_);
  and (_38533_, _38532_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not (_38534_, _38533_);
  nor (_38535_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38536_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38537_, _38536_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38538_, _38537_, _38535_);
  nor (_38539_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38540_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38541_, _38540_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38542_, _38541_, _38539_);
  nor (_38543_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38544_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38545_, _38544_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38546_, _38545_, _38543_);
  nor (_38547_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38548_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38549_, _38548_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38550_, _38549_, _38547_);
  nor (_38551_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38552_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38553_, _38552_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38554_, _38553_, _38551_);
  not (_38555_, _38554_);
  nor (_38556_, _38555_, _30755_);
  nor (_38557_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38558_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38559_, _38558_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38560_, _38559_, _38557_);
  and (_38561_, _38560_, _38556_);
  nor (_38562_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38563_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38564_, _38563_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38565_, _38564_, _38562_);
  and (_38566_, _38565_, _38561_);
  and (_38567_, _38566_, _38550_);
  nor (_38568_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38569_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38570_, _38569_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38571_, _38570_, _38568_);
  and (_38572_, _38571_, _38567_);
  and (_38573_, _38572_, _38546_);
  and (_38574_, _38573_, _38542_);
  nand (_38575_, _38574_, _38538_);
  or (_38576_, _38574_, _38538_);
  and (_38577_, _38576_, _38575_);
  and (_38578_, _38577_, _29271_);
  not (_38579_, _38578_);
  and (_38580_, _23318_, _18265_);
  and (_38581_, _29763_, _20334_);
  and (_38582_, _38581_, _28405_);
  and (_38583_, _38582_, _28437_);
  and (_38584_, _38583_, _28481_);
  and (_38585_, _38584_, _29084_);
  nor (_38586_, _38585_, _29785_);
  and (_38587_, _29007_, _18834_);
  nor (_38588_, _38587_, _38586_);
  and (_38589_, _29851_, _20323_);
  and (_38590_, _19653_, _18669_);
  and (_38591_, _19975_, _18988_);
  and (_38592_, _38591_, _38590_);
  and (_38593_, _38592_, _38589_);
  and (_38594_, _19805_, _18834_);
  and (_38595_, _38594_, _38593_);
  nor (_38596_, _38595_, _29007_);
  and (_38597_, _29007_, _19805_);
  nor (_38598_, _38597_, _38596_);
  and (_38599_, _38598_, _38588_);
  nor (_38600_, _29007_, _19164_);
  and (_38601_, _29007_, _19164_);
  nor (_38602_, _38601_, _38600_);
  and (_38603_, _38602_, _38599_);
  and (_38604_, _38603_, _29927_);
  nor (_38605_, _38603_, _29927_);
  nor (_38606_, _38605_, _38604_);
  and (_38607_, _38606_, _29698_);
  and (_38608_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_38609_, _29007_, _29927_);
  nor (_38610_, _38609_, _30864_);
  nor (_38611_, _38610_, _29981_);
  nor (_38612_, _31093_, _21052_);
  nor (_38613_, _30385_, _20149_);
  or (_38614_, _38613_, _38612_);
  or (_38615_, _38614_, _38611_);
  nor (_38616_, _38615_, _38608_);
  not (_38617_, _38616_);
  nor (_38618_, _38617_, _38607_);
  not (_38619_, _38618_);
  nor (_38620_, _38619_, _38580_);
  and (_38621_, _38620_, _38579_);
  nor (_38622_, _38621_, _38534_);
  and (_38623_, _38405_, _34004_);
  and (_38624_, _38623_, _38401_);
  or (_38625_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_38626_, _38625_, _38534_);
  nand (_38627_, _38624_, _30603_);
  and (_38628_, _38627_, _38626_);
  or (_38629_, _38628_, _38622_);
  and (_12713_, _38629_, _42882_);
  and (_38630_, _38405_, _33296_);
  and (_38631_, _38630_, _38401_);
  nor (_38632_, _38631_, _38533_);
  not (_38633_, _38632_);
  nand (_38634_, _38633_, _30603_);
  or (_38635_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38636_, _38635_, _42882_);
  and (_12734_, _38636_, _38634_);
  and (_38637_, _25917_, _23626_);
  not (_38638_, _38637_);
  and (_38639_, _38555_, _30755_);
  nor (_38640_, _38639_, _38556_);
  and (_38641_, _38640_, _29271_);
  nor (_38642_, _30864_, _29960_);
  not (_38643_, _38642_);
  nor (_38644_, _38643_, _29872_);
  nor (_38645_, _38644_, _28405_);
  and (_38646_, _38644_, _28405_);
  nor (_38647_, _38646_, _38645_);
  and (_38648_, _38647_, _29698_);
  nor (_38649_, _30385_, _18988_);
  and (_38650_, _23096_, _18265_);
  nor (_38651_, _31093_, _20693_);
  nor (_38652_, _29981_, _21922_);
  or (_38653_, _38652_, _38651_);
  or (_38654_, _38653_, _38650_);
  nor (_38655_, _38654_, _38649_);
  not (_38656_, _38655_);
  nor (_38657_, _38656_, _38648_);
  not (_38658_, _38657_);
  nor (_38659_, _38658_, _38641_);
  and (_38660_, _38659_, _38638_);
  nor (_38661_, _38660_, _38534_);
  or (_38662_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_38663_, _38662_, _38534_);
  nand (_38664_, _38624_, _31782_);
  and (_38665_, _38664_, _38663_);
  or (_38666_, _38665_, _38661_);
  and (_13647_, _38666_, _42882_);
  nor (_38667_, _38560_, _38556_);
  nor (_38668_, _38667_, _38561_);
  and (_38669_, _38668_, _29271_);
  not (_38670_, _38669_);
  and (_38671_, _24909_, _23626_);
  nor (_38672_, _20323_, _18988_);
  and (_38673_, _38672_, _29763_);
  and (_38674_, _38673_, _29007_);
  and (_38675_, _38589_, _18988_);
  and (_38676_, _38675_, _29785_);
  nor (_38677_, _38676_, _38674_);
  nor (_38678_, _38677_, _28437_);
  and (_38679_, _38677_, _28437_);
  nor (_38680_, _38679_, _38678_);
  nor (_38681_, _38680_, _33589_);
  nor (_38682_, _30385_, _19975_);
  and (_38683_, _23128_, _18265_);
  nor (_38684_, _31093_, _20519_);
  nor (_38685_, _29981_, _21379_);
  or (_38686_, _38685_, _38684_);
  or (_38687_, _38686_, _38683_);
  nor (_38688_, _38687_, _38682_);
  not (_38689_, _38688_);
  nor (_38690_, _38689_, _38681_);
  not (_38691_, _38690_);
  nor (_38692_, _38691_, _38671_);
  and (_38693_, _38692_, _38670_);
  nor (_38694_, _38693_, _38534_);
  or (_38695_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_38696_, _38695_, _38534_);
  nand (_38697_, _38624_, _32458_);
  and (_38698_, _38697_, _38696_);
  or (_38699_, _38698_, _38694_);
  and (_13657_, _38699_, _42882_);
  nor (_38700_, _38565_, _38561_);
  nor (_38701_, _38700_, _38566_);
  and (_38702_, _38701_, _29271_);
  not (_38703_, _38702_);
  and (_38704_, _38675_, _19975_);
  and (_38705_, _38704_, _29785_);
  and (_38706_, _38673_, _28437_);
  and (_38707_, _38706_, _29007_);
  nor (_38708_, _38707_, _38705_);
  and (_38709_, _38708_, _18669_);
  nor (_38710_, _38708_, _18669_);
  nor (_38711_, _38710_, _38709_);
  and (_38712_, _38711_, _29698_);
  not (_38713_, _38712_);
  nor (_38714_, _29981_, _21553_);
  and (_38715_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38716_, _38715_, _38714_);
  and (_38717_, _23159_, _18265_);
  nor (_38718_, _31093_, _19479_);
  nor (_38719_, _30385_, _18669_);
  or (_38720_, _38719_, _38718_);
  nor (_38721_, _38720_, _38717_);
  and (_38722_, _38721_, _38716_);
  and (_38723_, _38722_, _38713_);
  and (_38724_, _38723_, _38703_);
  nor (_38725_, _38724_, _38534_);
  or (_38726_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_38727_, _38726_, _38534_);
  nand (_38728_, _38624_, _33154_);
  and (_38729_, _38728_, _38727_);
  or (_38730_, _38729_, _38725_);
  and (_13668_, _38730_, _42882_);
  nor (_38731_, _38566_, _38550_);
  not (_38732_, _38731_);
  nor (_38733_, _38567_, _30744_);
  and (_38734_, _38733_, _38732_);
  not (_38735_, _38734_);
  and (_38736_, _23191_, _18265_);
  not (_38737_, _38736_);
  nor (_38738_, _38584_, _29084_);
  not (_38739_, _38738_);
  and (_38740_, _38739_, _38586_);
  and (_38741_, _38704_, _18669_);
  nor (_38742_, _38741_, _19653_);
  nor (_38743_, _38742_, _38593_);
  nor (_38744_, _38743_, _29007_);
  nor (_38745_, _38744_, _38740_);
  nor (_38746_, _38745_, _33589_);
  nor (_38747_, _30385_, _19653_);
  nor (_38748_, _29981_, _21052_);
  and (_38749_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_38750_, _38749_, _38748_);
  or (_38751_, _38750_, _31104_);
  nor (_38752_, _38751_, _38747_);
  not (_38753_, _38752_);
  nor (_38754_, _38753_, _38746_);
  and (_38755_, _38754_, _38737_);
  and (_38756_, _38755_, _38735_);
  nor (_38757_, _38756_, _38534_);
  or (_38758_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_38759_, _38758_, _38534_);
  nand (_38760_, _38624_, _33906_);
  and (_38761_, _38760_, _38759_);
  or (_38762_, _38761_, _38757_);
  and (_13679_, _38762_, _42882_);
  nor (_38763_, _38571_, _38567_);
  nor (_38764_, _38763_, _38572_);
  and (_38765_, _38764_, _29271_);
  not (_38766_, _38765_);
  and (_38767_, _23223_, _18265_);
  nor (_38768_, _38593_, _29007_);
  nor (_38769_, _38768_, _38586_);
  nor (_38770_, _38769_, _28120_);
  and (_38771_, _38769_, _28120_);
  nor (_38772_, _38771_, _38770_);
  and (_38773_, _38772_, _29698_);
  and (_38774_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_38775_, _29007_, _20704_);
  or (_38776_, _38775_, _29981_);
  nor (_38777_, _38776_, _38587_);
  nor (_38778_, _31093_, _21922_);
  nor (_38779_, _30385_, _18834_);
  or (_38780_, _38779_, _38778_);
  or (_38781_, _38780_, _38777_);
  nor (_38782_, _38781_, _38774_);
  not (_38783_, _38782_);
  nor (_38784_, _38783_, _38773_);
  not (_38785_, _38784_);
  nor (_38786_, _38785_, _38767_);
  and (_38787_, _38786_, _38766_);
  nor (_38788_, _38787_, _38534_);
  or (_38789_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_38790_, _38789_, _38534_);
  nand (_38791_, _38624_, _34667_);
  and (_38792_, _38791_, _38790_);
  or (_38793_, _38792_, _38788_);
  and (_13690_, _38793_, _42882_);
  nor (_38794_, _38572_, _38546_);
  not (_38795_, _38794_);
  nor (_38796_, _38573_, _30744_);
  and (_38797_, _38796_, _38795_);
  not (_38798_, _38797_);
  and (_38799_, _23255_, _18265_);
  and (_38800_, _38593_, _18834_);
  nor (_38801_, _38800_, _29007_);
  not (_38802_, _38801_);
  and (_38803_, _38802_, _38588_);
  and (_38804_, _38803_, _19805_);
  nor (_38805_, _38803_, _19805_);
  nor (_38806_, _38805_, _38804_);
  nor (_38807_, _38806_, _33589_);
  and (_38808_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_38809_, _29007_, _20530_);
  or (_38810_, _38809_, _29981_);
  nor (_38811_, _38810_, _38597_);
  nor (_38812_, _31093_, _21379_);
  nor (_38813_, _30385_, _19805_);
  or (_38814_, _38813_, _38812_);
  or (_38815_, _38814_, _38811_);
  nor (_38816_, _38815_, _38808_);
  not (_38817_, _38816_);
  nor (_38818_, _38817_, _38807_);
  not (_38819_, _38818_);
  nor (_38820_, _38819_, _38799_);
  and (_38821_, _38820_, _38798_);
  nor (_38822_, _38821_, _38534_);
  or (_38823_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_38824_, _38823_, _38534_);
  nand (_38825_, _38624_, _35461_);
  and (_38826_, _38825_, _38824_);
  or (_38827_, _38826_, _38822_);
  and (_13701_, _38827_, _42882_);
  nor (_38828_, _38573_, _38542_);
  nor (_38829_, _38828_, _38574_);
  and (_38830_, _38829_, _29271_);
  and (_38831_, _23286_, _18265_);
  and (_38832_, _38599_, _19164_);
  nor (_38833_, _38599_, _19164_);
  or (_38834_, _38833_, _38832_);
  and (_38835_, _38834_, _29698_);
  or (_38836_, _29007_, _19490_);
  nor (_38837_, _38601_, _29981_);
  and (_38838_, _38837_, _38836_);
  nor (_38839_, _31093_, _21553_);
  nor (_38840_, _30385_, _19164_);
  and (_38841_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or (_38842_, _38841_, _38840_);
  or (_38843_, _38842_, _38839_);
  or (_38844_, _38843_, _38838_);
  or (_38845_, _38844_, _38835_);
  or (_38846_, _38845_, _38831_);
  or (_38847_, _38846_, _38830_);
  and (_38848_, _38847_, _38533_);
  or (_38849_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_38850_, _38849_, _38534_);
  nand (_38851_, _38624_, _36179_);
  and (_38852_, _38851_, _38850_);
  or (_38853_, _38852_, _38848_);
  and (_13712_, _38853_, _42882_);
  nand (_38854_, _38633_, _31782_);
  or (_38855_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_38856_, _38855_, _42882_);
  and (_13723_, _38856_, _38854_);
  nand (_38857_, _38633_, _32458_);
  or (_38858_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38859_, _38858_, _42882_);
  and (_13733_, _38859_, _38857_);
  nand (_38860_, _38633_, _33154_);
  or (_38861_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38862_, _38861_, _42882_);
  and (_13744_, _38862_, _38860_);
  nand (_38863_, _38633_, _33906_);
  or (_38864_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38865_, _38864_, _42882_);
  and (_13755_, _38865_, _38863_);
  nand (_38866_, _38633_, _34667_);
  or (_38867_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38868_, _38867_, _42882_);
  and (_13766_, _38868_, _38866_);
  nand (_38869_, _38633_, _35461_);
  or (_38870_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38871_, _38870_, _42882_);
  and (_13777_, _38871_, _38869_);
  nand (_38872_, _38633_, _36179_);
  or (_38873_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38874_, _38873_, _42882_);
  and (_13788_, _38874_, _38872_);
  nor (_38875_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_38876_, _38875_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_38877_, _38875_, _31282_);
  or (_38878_, _38877_, _38876_);
  not (_38879_, _27374_);
  nor (_38880_, _38879_, _27242_);
  and (_38881_, _38880_, _31348_);
  and (_38882_, _38881_, _27867_);
  not (_38883_, _38882_);
  and (_38884_, _38883_, _38878_);
  and (_38885_, _38880_, _27867_);
  and (_38886_, _38885_, _31348_);
  not (_38887_, _31304_);
  nor (_38888_, _38887_, _31282_);
  not (_38889_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_38890_, _31304_, _38889_);
  or (_38891_, _38890_, _38888_);
  and (_38892_, _38891_, _38886_);
  or (_38893_, _38892_, _38884_);
  and (_38894_, _38401_, _27045_);
  nor (_38895_, _27242_, _27549_);
  nor (_38896_, _27845_, _38879_);
  and (_38897_, _38896_, _38895_);
  and (_38898_, _38897_, _38894_);
  or (_38899_, _38898_, _38893_);
  and (_38900_, _38894_, _38895_);
  and (_38901_, _38900_, _38896_);
  nand (_38902_, _38901_, _38485_);
  and (_38903_, _38902_, _42882_);
  and (_15193_, _38903_, _38899_);
  not (_38904_, _38901_);
  not (_38905_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_38906_, _38886_, _32567_);
  nand (_38907_, _38906_, _38905_);
  and (_38908_, _38907_, _38904_);
  or (_38909_, _38906_, _31859_);
  and (_38910_, _38909_, _38908_);
  nor (_38911_, _38904_, _38456_);
  or (_38912_, _38911_, _38910_);
  and (_17374_, _38912_, _42882_);
  or (_38913_, _30799_, _29183_);
  not (_38914_, _30788_);
  nand (_38915_, _38914_, _29183_);
  and (_38916_, _38915_, _27955_);
  and (_38917_, _38916_, _38913_);
  not (_38918_, _27977_);
  nand (_38919_, _29633_, _38918_);
  or (_38920_, _29633_, _27988_);
  and (_38921_, _29271_, _38920_);
  and (_38922_, _38921_, _38919_);
  and (_38923_, _38594_, _24810_);
  and (_38924_, _38592_, _23626_);
  nand (_38925_, _38924_, _38923_);
  nand (_38926_, _38925_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_38927_, _38926_, _38922_);
  or (_38928_, _38927_, _38917_);
  or (_38929_, _23381_, _23350_);
  or (_38930_, _38929_, _23413_);
  or (_38931_, _38930_, _23466_);
  or (_38932_, _38931_, _23487_);
  or (_38933_, _38932_, _23530_);
  or (_38934_, _38933_, _23562_);
  and (_38935_, _38934_, _18265_);
  or (_38936_, _38935_, _38928_);
  or (_38937_, _38936_, _27922_);
  nor (_38938_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_38939_, _38938_, _38882_);
  and (_38940_, _38939_, _38937_);
  and (_38941_, _33307_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_38942_, _38941_, _33318_);
  and (_38943_, _38942_, _38886_);
  or (_38944_, _38943_, _38898_);
  or (_38945_, _38944_, _38940_);
  nand (_38946_, _38901_, _38449_);
  and (_38947_, _38946_, _42882_);
  and (_17385_, _38947_, _38945_);
  not (_38948_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_38949_, _38886_, _34004_);
  nand (_38950_, _38949_, _38948_);
  and (_38951_, _38950_, _38904_);
  or (_38952_, _38949_, _31859_);
  and (_38953_, _38952_, _38951_);
  nor (_38954_, _38904_, _38442_);
  or (_38957_, _38954_, _38953_);
  and (_17396_, _38957_, _42882_);
  or (_38959_, _38883_, _34787_);
  and (_38960_, _38959_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_38961_, _34776_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_38962_, _38961_, _34819_);
  and (_38963_, _38962_, _38886_);
  or (_38964_, _38963_, _38960_);
  and (_38965_, _38964_, _38904_);
  nor (_38966_, _38904_, _38434_);
  or (_38967_, _38966_, _38965_);
  and (_17407_, _38967_, _42882_);
  not (_38977_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand (_38983_, _38886_, _35549_);
  nand (_38989_, _38983_, _38977_);
  and (_38992_, _38989_, _38904_);
  or (_38993_, _38983_, _31859_);
  and (_38994_, _38993_, _38992_);
  nor (_38995_, _38904_, _38428_);
  or (_38996_, _38995_, _38994_);
  and (_17418_, _38996_, _42882_);
  nand (_38997_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_38998_, _29271_, _29534_);
  and (_38999_, _29139_, _27955_);
  nor (_39000_, _38999_, _38998_);
  nor (_39001_, _39000_, _38997_);
  or (_39002_, _38997_, _30374_);
  and (_39003_, _39002_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_39004_, _39003_, _38882_);
  or (_39005_, _39004_, _39001_);
  not (_39006_, _36277_);
  nor (_39007_, _39006_, _31282_);
  or (_39008_, _36277_, _33644_);
  nand (_39009_, _39008_, _38882_);
  or (_39010_, _39009_, _39007_);
  and (_39011_, _39010_, _39005_);
  or (_39012_, _39011_, _38901_);
  nand (_39013_, _38901_, _38420_);
  and (_39014_, _39013_, _42882_);
  and (_17429_, _39014_, _39012_);
  not (_39017_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39018_, _38532_, _39017_);
  not (_39019_, _39018_);
  nor (_39020_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_39021_, _39020_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39022_, _27045_, _27703_);
  and (_39023_, _27845_, _38879_);
  and (_39024_, _39023_, _38895_);
  and (_39025_, _39024_, _39022_);
  and (_39026_, _39025_, _30679_);
  nor (_39027_, _39026_, _39021_);
  nor (_39028_, _39027_, _30603_);
  and (_39029_, _27845_, _27703_);
  not (_39030_, _31348_);
  nor (_39031_, _39030_, _27549_);
  and (_39032_, _39031_, _27385_);
  and (_39033_, _39032_, _39029_);
  and (_39034_, _39033_, _31304_);
  and (_39035_, _39034_, _31282_);
  nor (_39036_, _39034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_39037_, _39036_);
  and (_39038_, _39027_, _39019_);
  and (_39039_, _39038_, _39037_);
  not (_39040_, _39039_);
  nor (_39041_, _39040_, _39035_);
  or (_39042_, _39041_, _39028_);
  and (_39043_, _39042_, _39019_);
  nor (_39044_, _39019_, _38621_);
  or (_39045_, _39044_, _39043_);
  and (_17998_, _39045_, _42882_);
  nor (_39046_, _39019_, _38660_);
  nor (_39047_, _39027_, _31783_);
  not (_39048_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_39049_, _39029_, _27560_);
  and (_39050_, _31348_, _27385_);
  and (_39051_, _39050_, _39049_);
  nor (_39052_, _39051_, _39048_);
  not (_39053_, _39052_);
  and (_39055_, _39053_, _39027_);
  not (_39059_, _39055_);
  not (_39065_, _27045_);
  nor (_39070_, _31282_, _39065_);
  nor (_39077_, _27045_, _39048_);
  nor (_39085_, _39077_, _39070_);
  and (_39093_, _39038_, _39051_);
  not (_39094_, _39093_);
  nor (_39095_, _39094_, _39085_);
  nor (_39096_, _39095_, _39059_);
  nor (_39097_, _39096_, _39018_);
  not (_39098_, _39097_);
  nor (_39099_, _39098_, _39047_);
  nor (_39100_, _39099_, _39046_);
  nor (_19849_, _39100_, rst);
  and (_39101_, _39018_, _38693_);
  nor (_39102_, _39027_, _32458_);
  and (_39103_, _39033_, _32567_);
  and (_39104_, _39103_, _31282_);
  nor (_39105_, _39103_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not (_39106_, _39105_);
  and (_39107_, _39106_, _39038_);
  not (_39108_, _39107_);
  nor (_39109_, _39108_, _39104_);
  nor (_39110_, _39109_, _39018_);
  not (_39111_, _39110_);
  nor (_39112_, _39111_, _39102_);
  nor (_39113_, _39112_, _39101_);
  and (_19860_, _39113_, _42882_);
  nor (_39114_, _39027_, _33154_);
  and (_39115_, _39033_, _33296_);
  and (_39116_, _39115_, _31282_);
  nor (_39117_, _39115_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_39118_, _39117_);
  and (_39119_, _39118_, _39038_);
  not (_39120_, _39119_);
  nor (_39121_, _39120_, _39116_);
  or (_39122_, _39121_, _39114_);
  and (_39123_, _39122_, _39019_);
  nor (_39124_, _39019_, _38724_);
  or (_39125_, _39124_, _39123_);
  and (_19872_, _39125_, _42882_);
  nor (_39126_, _39027_, _33906_);
  not (_39127_, _39033_);
  and (_39133_, _39038_, _39127_);
  and (_39144_, _39133_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  not (_39145_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_39146_, _34004_, _39145_);
  nor (_39147_, _39146_, _34015_);
  nor (_39158_, _39147_, _39094_);
  nor (_39164_, _39158_, _39144_);
  and (_39165_, _39164_, _39019_);
  not (_39166_, _39165_);
  nor (_39167_, _39166_, _39126_);
  and (_39168_, _39018_, _38756_);
  or (_39169_, _39168_, _39167_);
  nor (_19884_, _39169_, rst);
  nor (_39170_, _39027_, _34667_);
  and (_39171_, _39033_, _34765_);
  and (_39172_, _39171_, _31282_);
  nor (_39173_, _39171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_39174_, _39173_);
  and (_39175_, _39174_, _39038_);
  not (_39176_, _39175_);
  nor (_39177_, _39176_, _39172_);
  or (_39178_, _39177_, _39170_);
  and (_39179_, _39178_, _39019_);
  nor (_39180_, _39019_, _38787_);
  or (_39181_, _39180_, _39179_);
  and (_19896_, _39181_, _42882_);
  nor (_39182_, _39027_, _35461_);
  and (_39183_, _39033_, _35549_);
  and (_39184_, _39183_, _31282_);
  nor (_39185_, _39183_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not (_39186_, _39185_);
  and (_39187_, _39186_, _39038_);
  not (_39188_, _39187_);
  nor (_39189_, _39188_, _39184_);
  or (_39190_, _39189_, _39182_);
  and (_39191_, _39190_, _39019_);
  nor (_39192_, _39019_, _38821_);
  or (_39193_, _39192_, _39191_);
  and (_19908_, _39193_, _42882_);
  nor (_39194_, _39027_, _36179_);
  and (_39195_, _39133_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_39196_, _39006_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_39197_, _39196_, _39007_);
  nor (_39198_, _39197_, _39094_);
  nor (_39199_, _39198_, _39195_);
  and (_39200_, _39199_, _39019_);
  not (_39201_, _39200_);
  nor (_39202_, _39201_, _39194_);
  nor (_39203_, _39019_, _38847_);
  or (_39204_, _39203_, _39202_);
  nor (_19920_, _39204_, rst);
  and (_39205_, _27374_, _27242_);
  and (_39206_, _39049_, _39205_);
  and (_39207_, _39206_, _31304_);
  nand (_39208_, _39207_, _31282_);
  or (_39209_, _39207_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39210_, _39209_, _31348_);
  and (_39211_, _39210_, _39208_);
  and (_39212_, _38405_, _39022_);
  nand (_39213_, _39212_, _38485_);
  or (_39214_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39215_, _39214_, _30679_);
  and (_39216_, _39215_, _39213_);
  not (_39217_, _30668_);
  and (_39218_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_39219_, _39218_, rst);
  or (_39220_, _39219_, _39216_);
  or (_31126_, _39220_, _39211_);
  and (_39221_, _39205_, _27867_);
  and (_39222_, _39221_, _31304_);
  nand (_39223_, _39222_, _31282_);
  or (_39224_, _39222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39225_, _39224_, _31348_);
  and (_39226_, _39225_, _39223_);
  and (_39227_, _38896_, _38404_);
  and (_39228_, _39227_, _39022_);
  nand (_39229_, _39228_, _38485_);
  or (_39230_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39231_, _39230_, _30679_);
  and (_39232_, _39231_, _39229_);
  and (_39233_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_39234_, _39233_, rst);
  or (_39235_, _39234_, _39232_);
  or (_31149_, _39235_, _39226_);
  and (_39236_, _38879_, _27242_);
  and (_39237_, _39236_, _39049_);
  and (_39238_, _39237_, _31304_);
  nand (_39239_, _39238_, _31282_);
  or (_39240_, _39238_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_39241_, _39240_, _31348_);
  and (_39242_, _39241_, _39239_);
  and (_39243_, _39023_, _38404_);
  and (_39244_, _39243_, _39022_);
  not (_39245_, _39244_);
  nor (_39246_, _39245_, _38485_);
  and (_39247_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_39248_, _39247_, _39246_);
  and (_39249_, _39248_, _30679_);
  and (_39250_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_39251_, _39250_, rst);
  or (_39252_, _39251_, _39249_);
  or (_31172_, _39252_, _39242_);
  and (_39253_, _39236_, _27867_);
  and (_39254_, _39253_, _31304_);
  nand (_39255_, _39254_, _31282_);
  or (_39256_, _39254_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_39257_, _39256_, _31348_);
  and (_39258_, _39257_, _39255_);
  nor (_39259_, _27845_, _27374_);
  and (_39260_, _38404_, _39259_);
  and (_39261_, _39260_, _39022_);
  not (_39262_, _39261_);
  nor (_39263_, _39262_, _38485_);
  and (_39264_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_39265_, _39264_, _39263_);
  and (_39266_, _39265_, _30679_);
  and (_39267_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_39268_, _39267_, rst);
  or (_39269_, _39268_, _39266_);
  or (_31194_, _39269_, _39258_);
  or (_39270_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_39271_, _39270_, _31348_);
  nand (_39272_, _39212_, _31282_);
  and (_39273_, _39272_, _39271_);
  nand (_39274_, _39212_, _38464_);
  and (_39275_, _39274_, _30679_);
  and (_39276_, _39275_, _39270_);
  and (_39277_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_39278_, _39277_, rst);
  or (_39279_, _39278_, _39276_);
  or (_40589_, _39279_, _39273_);
  and (_39280_, _32567_, _27703_);
  and (_39281_, _39280_, _38405_);
  nand (_39282_, _39281_, _31282_);
  or (_39283_, _39281_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39284_, _39283_, _31348_);
  and (_39285_, _39284_, _39282_);
  nand (_39286_, _39212_, _38456_);
  or (_39287_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39288_, _39287_, _30679_);
  and (_39289_, _39288_, _39286_);
  and (_39290_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_39291_, _39290_, rst);
  or (_39292_, _39291_, _39289_);
  or (_40591_, _39292_, _39285_);
  not (_39293_, _34026_);
  nand (_39294_, _39206_, _39293_);
  and (_39295_, _39294_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39296_, _33329_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39297_, _39296_, _33318_);
  and (_39298_, _39297_, _39206_);
  or (_39299_, _39298_, _39295_);
  and (_39300_, _39299_, _31348_);
  nand (_39301_, _39212_, _38449_);
  or (_39302_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39303_, _39302_, _30679_);
  and (_39304_, _39303_, _39301_);
  and (_39305_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39306_, _39305_, rst);
  or (_39307_, _39306_, _39304_);
  or (_40593_, _39307_, _39300_);
  nand (_39308_, _39206_, _26781_);
  and (_39309_, _39308_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39310_, _39293_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_39311_, _39310_, _34015_);
  and (_39312_, _39311_, _39206_);
  or (_39313_, _39312_, _39309_);
  and (_39314_, _39313_, _31348_);
  nand (_39315_, _39212_, _38442_);
  or (_39316_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39317_, _39316_, _30679_);
  and (_39318_, _39317_, _39315_);
  and (_39319_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_39320_, _39319_, rst);
  or (_39321_, _39320_, _39318_);
  or (_40595_, _39321_, _39314_);
  not (_39322_, _39206_);
  or (_39323_, _39322_, _34787_);
  and (_39324_, _39323_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39325_, _34776_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39326_, _39325_, _34819_);
  and (_39327_, _39326_, _39206_);
  or (_39328_, _39327_, _39324_);
  and (_39329_, _39328_, _31348_);
  nand (_39330_, _39212_, _38434_);
  or (_39331_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39332_, _39331_, _30679_);
  and (_39333_, _39332_, _39330_);
  and (_39334_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39335_, _39334_, rst);
  or (_39336_, _39335_, _39333_);
  or (_40597_, _39336_, _39329_);
  and (_39337_, _39206_, _35549_);
  nand (_39338_, _39337_, _31282_);
  or (_39347_, _39337_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39358_, _39347_, _31348_);
  and (_39369_, _39358_, _39338_);
  nand (_39378_, _39212_, _38428_);
  or (_39384_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39395_, _39384_, _30679_);
  and (_39406_, _39395_, _39378_);
  and (_39417_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39428_, _39417_, rst);
  or (_39439_, _39428_, _39406_);
  or (_40599_, _39439_, _39369_);
  and (_39460_, _39206_, _36277_);
  nand (_39471_, _39460_, _31282_);
  or (_39482_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39493_, _39482_, _31348_);
  and (_39504_, _39493_, _39471_);
  nand (_39515_, _39212_, _38420_);
  or (_39526_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39537_, _39526_, _30679_);
  and (_39548_, _39537_, _39515_);
  and (_39552_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_39553_, _39552_, rst);
  or (_39554_, _39553_, _39548_);
  or (_40601_, _39554_, _39504_);
  and (_39555_, _39221_, _27045_);
  nand (_39556_, _39555_, _31282_);
  or (_39557_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39558_, _39557_, _31348_);
  and (_39559_, _39558_, _39556_);
  nand (_39560_, _39228_, _38464_);
  and (_39561_, _39560_, _30679_);
  and (_39562_, _39561_, _39557_);
  and (_39563_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_39564_, _39563_, rst);
  or (_39565_, _39564_, _39562_);
  or (_40603_, _39565_, _39559_);
  and (_39566_, _39221_, _32567_);
  nand (_39567_, _39566_, _31282_);
  or (_39568_, _39566_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39569_, _39568_, _31348_);
  and (_39570_, _39569_, _39567_);
  nand (_39571_, _39228_, _38456_);
  or (_39572_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39573_, _39572_, _30679_);
  and (_39574_, _39573_, _39571_);
  and (_39575_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39576_, _39575_, rst);
  or (_39577_, _39576_, _39574_);
  or (_40605_, _39577_, _39570_);
  and (_39578_, _39221_, _33296_);
  nand (_39579_, _39578_, _31282_);
  or (_39580_, _39578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39581_, _39580_, _31348_);
  and (_39582_, _39581_, _39579_);
  nand (_39583_, _39228_, _38449_);
  or (_39584_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39585_, _39584_, _30679_);
  and (_39586_, _39585_, _39583_);
  and (_39587_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_39588_, _39587_, rst);
  or (_39589_, _39588_, _39586_);
  or (_40607_, _39589_, _39582_);
  and (_39590_, _39221_, _34004_);
  nand (_39591_, _39590_, _31282_);
  or (_39592_, _39590_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39593_, _39592_, _31348_);
  and (_39594_, _39593_, _39591_);
  nand (_39595_, _39228_, _38442_);
  or (_39596_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39597_, _39596_, _30679_);
  and (_39598_, _39597_, _39595_);
  and (_39599_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39600_, _39599_, rst);
  or (_39601_, _39600_, _39598_);
  or (_40609_, _39601_, _39594_);
  and (_39602_, _39221_, _34765_);
  nand (_39603_, _39602_, _31282_);
  or (_39604_, _39602_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39605_, _39604_, _31348_);
  and (_39606_, _39605_, _39603_);
  nand (_39607_, _39228_, _38434_);
  or (_39608_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39609_, _39608_, _30679_);
  and (_39610_, _39609_, _39607_);
  and (_39611_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39612_, _39611_, rst);
  or (_39613_, _39612_, _39610_);
  or (_40611_, _39613_, _39606_);
  and (_39614_, _39221_, _35549_);
  nand (_39615_, _39614_, _31282_);
  or (_39616_, _39614_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39617_, _39616_, _31348_);
  and (_39618_, _39617_, _39615_);
  nand (_39619_, _39228_, _38428_);
  or (_39620_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39621_, _39620_, _30679_);
  and (_39622_, _39621_, _39619_);
  and (_39623_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39624_, _39623_, rst);
  or (_39625_, _39624_, _39622_);
  or (_40612_, _39625_, _39618_);
  and (_39626_, _39221_, _36277_);
  nand (_39627_, _39626_, _31282_);
  or (_39628_, _39626_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39629_, _39628_, _31348_);
  and (_39630_, _39629_, _39627_);
  nand (_39631_, _39228_, _38420_);
  or (_39632_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39633_, _39632_, _30679_);
  and (_39634_, _39633_, _39631_);
  and (_39635_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39636_, _39635_, rst);
  or (_39637_, _39636_, _39634_);
  or (_40614_, _39637_, _39630_);
  nand (_39638_, _39244_, _31282_);
  or (_39639_, _39244_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39640_, _39639_, _31348_);
  and (_39641_, _39640_, _39638_);
  and (_39642_, _39244_, _38465_);
  and (_39643_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_39644_, _39643_, _39642_);
  and (_39645_, _39644_, _30679_);
  and (_39646_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_39647_, _39646_, rst);
  or (_39648_, _39647_, _39645_);
  or (_40616_, _39648_, _39641_);
  and (_39649_, _39237_, _32567_);
  nand (_39650_, _39649_, _31282_);
  or (_39651_, _39649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39652_, _39651_, _31348_);
  and (_39653_, _39652_, _39650_);
  nor (_39654_, _39245_, _38456_);
  and (_39655_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39656_, _39655_, _39654_);
  and (_39657_, _39656_, _30679_);
  and (_39658_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39659_, _39658_, rst);
  or (_39660_, _39659_, _39657_);
  or (_40618_, _39660_, _39653_);
  and (_39661_, _39237_, _33296_);
  nand (_39662_, _39661_, _31282_);
  or (_39663_, _39661_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39664_, _39663_, _31348_);
  and (_39665_, _39664_, _39662_);
  nor (_39666_, _39245_, _38449_);
  and (_39667_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39668_, _39667_, _39666_);
  and (_39669_, _39668_, _30679_);
  and (_39670_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39671_, _39670_, rst);
  or (_39672_, _39671_, _39669_);
  or (_40620_, _39672_, _39665_);
  and (_39673_, _39237_, _34004_);
  nand (_39674_, _39673_, _31282_);
  or (_39675_, _39673_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39676_, _39675_, _31348_);
  and (_39677_, _39676_, _39674_);
  nor (_39678_, _39245_, _38442_);
  and (_39679_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39680_, _39679_, _39678_);
  and (_39681_, _39680_, _30679_);
  and (_39682_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39683_, _39682_, rst);
  or (_39684_, _39683_, _39681_);
  or (_40622_, _39684_, _39677_);
  and (_39685_, _39237_, _34765_);
  nand (_39686_, _39685_, _31282_);
  or (_39687_, _39685_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39688_, _39687_, _31348_);
  and (_39689_, _39688_, _39686_);
  nor (_39690_, _39245_, _38434_);
  and (_39691_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39692_, _39691_, _39690_);
  and (_39693_, _39692_, _30679_);
  and (_39694_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39695_, _39694_, rst);
  or (_39696_, _39695_, _39693_);
  or (_40624_, _39696_, _39689_);
  and (_39697_, _39237_, _35549_);
  nand (_39698_, _39697_, _31282_);
  or (_39699_, _39697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39700_, _39699_, _31348_);
  and (_39701_, _39700_, _39698_);
  nor (_39702_, _39245_, _38428_);
  and (_39703_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39704_, _39703_, _39702_);
  and (_39705_, _39704_, _30679_);
  and (_39706_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39707_, _39706_, rst);
  or (_39708_, _39707_, _39705_);
  or (_40626_, _39708_, _39701_);
  and (_39709_, _39237_, _36277_);
  nand (_39710_, _39709_, _31282_);
  or (_39711_, _39709_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39712_, _39711_, _31348_);
  and (_39713_, _39712_, _39710_);
  nor (_39714_, _39245_, _38420_);
  and (_39715_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39716_, _39715_, _39714_);
  and (_39717_, _39716_, _30679_);
  and (_39718_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39719_, _39718_, rst);
  or (_39720_, _39719_, _39717_);
  or (_40628_, _39720_, _39713_);
  and (_39721_, _39253_, _27045_);
  nand (_39722_, _39721_, _31282_);
  or (_39723_, _39721_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39724_, _39723_, _31348_);
  and (_39725_, _39724_, _39722_);
  and (_39726_, _39261_, _38465_);
  and (_39727_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_39728_, _39727_, _39726_);
  and (_39729_, _39728_, _30679_);
  and (_39730_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_39731_, _39730_, rst);
  or (_39732_, _39731_, _39729_);
  or (_40630_, _39732_, _39725_);
  and (_39733_, _39253_, _32567_);
  nand (_39734_, _39733_, _31282_);
  or (_39735_, _39733_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39736_, _39735_, _31348_);
  and (_39737_, _39736_, _39734_);
  nor (_39738_, _39262_, _38456_);
  and (_39739_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39740_, _39739_, _39738_);
  and (_39741_, _39740_, _30679_);
  and (_39742_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39743_, _39742_, rst);
  or (_39744_, _39743_, _39741_);
  or (_40632_, _39744_, _39737_);
  and (_39745_, _39253_, _33296_);
  nand (_39746_, _39745_, _31282_);
  or (_39747_, _39745_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_39748_, _39747_, _31348_);
  and (_39749_, _39748_, _39746_);
  nor (_39750_, _39262_, _38449_);
  and (_39751_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39752_, _39751_, _39750_);
  and (_39753_, _39752_, _30679_);
  and (_39754_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39755_, _39754_, rst);
  or (_39756_, _39755_, _39753_);
  or (_40634_, _39756_, _39749_);
  and (_39757_, _39253_, _34004_);
  nand (_39758_, _39757_, _31282_);
  or (_39759_, _39757_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_39761_, _39759_, _31348_);
  and (_39766_, _39761_, _39758_);
  nor (_39767_, _39262_, _38442_);
  and (_39768_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39769_, _39768_, _39767_);
  and (_39770_, _39769_, _30679_);
  and (_39771_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39772_, _39771_, rst);
  or (_39773_, _39772_, _39770_);
  or (_40636_, _39773_, _39766_);
  and (_39774_, _39253_, _34765_);
  nand (_39775_, _39774_, _31282_);
  or (_39776_, _39774_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_39777_, _39776_, _31348_);
  and (_39778_, _39777_, _39775_);
  nor (_39779_, _39262_, _38434_);
  and (_39780_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39781_, _39780_, _39779_);
  and (_39782_, _39781_, _30679_);
  and (_39783_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39784_, _39783_, rst);
  or (_39785_, _39784_, _39782_);
  or (_40638_, _39785_, _39778_);
  and (_39786_, _39253_, _35549_);
  nand (_39787_, _39786_, _31282_);
  or (_39788_, _39786_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_39789_, _39788_, _31348_);
  and (_39790_, _39789_, _39787_);
  nor (_39791_, _39262_, _38428_);
  and (_39802_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39813_, _39802_, _39791_);
  and (_39822_, _39813_, _30679_);
  and (_39823_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39824_, _39823_, rst);
  or (_39825_, _39824_, _39822_);
  or (_40640_, _39825_, _39790_);
  and (_39826_, _39253_, _36277_);
  nand (_39827_, _39826_, _31282_);
  or (_39828_, _39826_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_39829_, _39828_, _31348_);
  and (_39830_, _39829_, _39827_);
  nor (_39831_, _39262_, _38420_);
  and (_39832_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39833_, _39832_, _39831_);
  and (_39834_, _39833_, _30679_);
  and (_39835_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39836_, _39835_, rst);
  or (_39837_, _39836_, _39834_);
  or (_40642_, _39837_, _39830_);
  and (_41092_, t0_i, _42882_);
  and (_41095_, t1_i, _42882_);
  not (_39838_, _30679_);
  nor (_39839_, _39838_, _27703_);
  and (_39840_, _39839_, _34004_);
  and (_39841_, _39840_, _38405_);
  nand (_39842_, _39841_, _38485_);
  nor (_39843_, _26781_, _27703_);
  and (_39844_, _39843_, _38406_);
  and (_39845_, _39844_, _30679_);
  not (_39846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_39847_, _39846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_39848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_39852_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _39848_);
  nor (_39856_, _39852_, _39847_);
  nor (_39857_, _39856_, _39845_);
  not (_39858_, _39857_);
  and (_39859_, _39858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_39860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_39861_, t1_i);
  and (_39862_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _39861_);
  nor (_39863_, _39862_, _39860_);
  not (_39864_, _39863_);
  not (_39865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_39866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _39865_);
  nor (_39867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_39868_, _39867_);
  and (_39869_, _39868_, _39866_);
  and (_39870_, _39869_, _39864_);
  not (_39871_, _39870_);
  nand (_39872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_39873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or (_39874_, _39873_, _39872_);
  nor (_39875_, _39874_, _39871_);
  and (_39876_, _39875_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_39877_, _39876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_39878_, _39877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_39879_, _39878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_39880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_39881_, _39874_, _39880_);
  and (_39882_, _39881_, _39870_);
  and (_39883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_39884_, _39883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_39885_, _39884_, _39882_);
  nor (_39886_, _39885_, _39856_);
  and (_39887_, _39886_, _39879_);
  and (_39888_, _39885_, _39847_);
  and (_39889_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39890_, _39889_, _39887_);
  nor (_39891_, _39890_, _39845_);
  or (_39892_, _39891_, _39859_);
  or (_39893_, _39841_, _39892_);
  and (_39894_, _39893_, _42882_);
  and (_41098_, _39894_, _39842_);
  nand (_39895_, _39845_, _38485_);
  and (_39896_, _39839_, _38623_);
  not (_39897_, _39896_);
  and (_39898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_39899_, _39898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_39900_, _39884_, _39881_);
  and (_39901_, _39900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_39902_, _39901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_39903_, _39902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_39904_, _39903_, _39870_);
  and (_39905_, _39904_, _39899_);
  and (_39906_, _39905_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_39907_, _39906_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39908_, _39906_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39909_, _39908_, _39907_);
  and (_39910_, _39909_, _39852_);
  and (_39911_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_39912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_39913_, _39912_, _39881_);
  and (_39914_, _39913_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_39915_, _39914_, _39870_);
  and (_39916_, _39915_, _39899_);
  and (_39917_, _39916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_39918_, _39917_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_39920_, _39917_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_39921_, _39920_, _39919_);
  nor (_39922_, _39921_, _39918_);
  or (_39923_, _39922_, _39911_);
  or (_39924_, _39923_, _39910_);
  or (_39925_, _39924_, _39845_);
  and (_39926_, _39925_, _39897_);
  and (_39927_, _39926_, _39895_);
  and (_39928_, _39896_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_39929_, _39928_, _39927_);
  and (_41101_, _39929_, _42882_);
  not (_39930_, _39845_);
  and (_39931_, _39871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or (_39932_, _39931_, _39907_);
  and (_39933_, _39932_, _39852_);
  or (_39934_, _39931_, _39918_);
  and (_39942_, _39934_, _39919_);
  nand (_39946_, _39870_, _39846_);
  and (_39947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_39948_, _39947_, _39946_);
  or (_39949_, _39948_, _39888_);
  or (_39950_, _39949_, _39942_);
  or (_39951_, _39950_, _39933_);
  nor (_39952_, _39896_, rst);
  and (_39953_, _39952_, _39951_);
  and (_41104_, _39953_, _39930_);
  and (_39954_, _39839_, _34765_);
  and (_39955_, _39954_, _38405_);
  nor (_39956_, _39955_, rst);
  and (_39957_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_39958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_39959_, _39958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_39960_, _39959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_39961_, _39960_, _39957_);
  and (_39962_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_39963_, _39962_, _39961_);
  or (_39964_, _39963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_39965_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_39966_, _39965_);
  and (_39967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_39968_, _39967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_39969_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_39970_, t0_i);
  and (_39971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _39970_);
  nor (_39972_, _39971_, _39969_);
  not (_39973_, _39972_);
  not (_39974_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_39975_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_39976_, _39975_, _39974_);
  and (_39977_, _39976_, _39973_);
  and (_39978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_39979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_39980_, _39979_, _39978_);
  and (_39981_, _39980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_39982_, _39981_, _39977_);
  and (_39983_, _39982_, _39968_);
  and (_39984_, _39983_, _39966_);
  and (_39985_, _39984_, _39964_);
  not (_39986_, _39977_);
  and (_39987_, _39986_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and (_39988_, _39982_, _39961_);
  and (_39989_, _39988_, _39962_);
  and (_39990_, _39989_, _39965_);
  or (_39991_, _39990_, _39987_);
  nor (_39992_, _39991_, _39985_);
  and (_39993_, _39839_, _33296_);
  and (_39994_, _39993_, _38405_);
  nor (_39995_, _39994_, _39992_);
  and (_41107_, _39995_, _39956_);
  and (_39996_, _39839_, _38630_);
  nand (_39997_, _39996_, _38485_);
  not (_39998_, _39955_);
  or (_39999_, _39998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_40000_, _39965_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_40001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_40002_, _40001_, _39982_);
  or (_40003_, _40002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_40004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_40005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _40004_);
  nand (_40006_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_40007_, _40006_, _39983_);
  and (_40008_, _40007_, _39966_);
  or (_40009_, _40008_, _39955_);
  and (_40010_, _40009_, _40003_);
  or (_40011_, _40010_, _40000_);
  and (_40012_, _40011_, _39999_);
  or (_40013_, _40012_, _39996_);
  and (_40014_, _40013_, _42882_);
  and (_41110_, _40014_, _39997_);
  nand (_40017_, _39955_, _38485_);
  not (_40020_, _39994_);
  and (_40021_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _40004_);
  or (_40022_, _40005_, _40021_);
  not (_40023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_40024_, _39981_, _39968_);
  and (_40025_, _39977_, _40004_);
  and (_40026_, _40025_, _40024_);
  and (_40027_, _40026_, _39961_);
  and (_40028_, _40027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_40029_, _40028_, _40023_);
  and (_40030_, _40028_, _40023_);
  or (_40031_, _40030_, _40029_);
  and (_40032_, _40031_, _40022_);
  and (_40033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_40035_, _40034_, _39960_);
  and (_40038_, _40035_, _39957_);
  and (_40046_, _40038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40047_, _40046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_40048_, _40034_, _39963_);
  and (_40049_, _40048_, _40047_);
  and (_40050_, _40049_, _40033_);
  and (_40051_, _39988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40052_, _40051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_40053_, _39989_, _39966_);
  and (_40054_, _40053_, _40052_);
  or (_40055_, _40054_, _40050_);
  or (_40056_, _40055_, _40032_);
  or (_40057_, _40056_, _39955_);
  and (_40058_, _40057_, _40020_);
  and (_40059_, _40058_, _40017_);
  and (_40060_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_40061_, _40060_, _40059_);
  and (_41113_, _40061_, _42882_);
  and (_40062_, _27023_, _33274_);
  nor (_40063_, _31283_, _27703_);
  and (_40064_, _40063_, _40062_);
  nand (_40065_, _40064_, _38405_);
  or (_40066_, _40065_, _39838_);
  not (_40067_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  or (_40068_, _40034_, _40067_);
  nand (_40069_, _40068_, _40048_);
  nand (_40070_, _40069_, _40033_);
  nor (_40071_, _40070_, _39955_);
  and (_40072_, _40071_, _40066_);
  and (_41116_, _40072_, _42882_);
  and (_40073_, _40063_, _38406_);
  and (_40074_, _40073_, _30679_);
  or (_40075_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_40076_, _40075_, _42882_);
  nand (_40077_, _40074_, _38485_);
  and (_41119_, _40077_, _40076_);
  not (_40078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_40079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_40080_, _40079_, _39845_);
  and (_40081_, _40080_, _39870_);
  nor (_40082_, _40081_, _40078_);
  and (_40083_, _40081_, _40078_);
  or (_40084_, _40083_, _40082_);
  nand (_40085_, _39901_, _39847_);
  nor (_40086_, _40085_, _39845_);
  or (_40087_, _40086_, _39841_);
  or (_40088_, _40087_, _40084_);
  nand (_40089_, _39841_, _38464_);
  and (_40090_, _40089_, _42882_);
  and (_41601_, _40090_, _40088_);
  and (_40091_, _39870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_40092_, _40091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_40093_, _40091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_40094_, _40093_, _40092_);
  nand (_40095_, _40094_, _40080_);
  or (_40096_, _40080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_40097_, _40096_, _40095_);
  nand (_40098_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_40099_, _40098_, _39845_);
  or (_40100_, _40099_, _39896_);
  or (_40101_, _40100_, _40097_);
  nand (_40102_, _39896_, _38456_);
  and (_40103_, _40102_, _42882_);
  and (_41603_, _40103_, _40101_);
  not (_40104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_40105_, _40080_, _40104_);
  nand (_40106_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_40107_, _40106_, _39845_);
  or (_40108_, _40107_, _40105_);
  nor (_40109_, _40092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_40110_, _40092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_40111_, _40110_, _40109_);
  and (_40112_, _40111_, _40080_);
  or (_40113_, _40112_, _39841_);
  or (_40114_, _40113_, _40108_);
  nand (_40115_, _39841_, _38449_);
  and (_40116_, _40115_, _42882_);
  and (_41605_, _40116_, _40114_);
  not (_40117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_40118_, _40080_, _40117_);
  or (_40119_, _40110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_40120_, _40079_, _39875_);
  and (_40121_, _40120_, _40119_);
  and (_40122_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_40123_, _40122_, _40121_);
  nor (_40124_, _40123_, _39845_);
  or (_40125_, _40124_, _40118_);
  and (_40126_, _40125_, _39897_);
  nor (_40127_, _39897_, _38442_);
  or (_40128_, _40127_, _40126_);
  and (_41606_, _40128_, _42882_);
  nor (_40129_, _39875_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_40130_, _40129_, _39882_);
  and (_40131_, _40130_, _40080_);
  nor (_40132_, _40080_, _39880_);
  nand (_40133_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_40134_, _40133_, _39845_);
  or (_40135_, _40134_, _40132_);
  or (_40136_, _40135_, _40131_);
  or (_40137_, _40136_, _39841_);
  nand (_40138_, _39841_, _38434_);
  and (_40139_, _40138_, _42882_);
  and (_41608_, _40139_, _40137_);
  nand (_40140_, _39841_, _38428_);
  and (_40141_, _39882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_40142_, _39882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_40143_, _40142_, _40141_);
  and (_40144_, _40143_, _39857_);
  and (_40145_, _39858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand (_40146_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_40147_, _40146_, _39845_);
  or (_40148_, _40147_, _40145_);
  or (_40149_, _40148_, _40144_);
  or (_40150_, _40149_, _39841_);
  and (_40151_, _40150_, _42882_);
  and (_41610_, _40151_, _40140_);
  nand (_40152_, _39841_, _38420_);
  and (_40153_, _39858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_40154_, _39847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40155_, _40154_, _39870_);
  and (_40156_, _40155_, _39900_);
  nor (_40157_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_40158_, _40157_, _39856_);
  nor (_40159_, _40158_, _39878_);
  nor (_40160_, _40159_, _40156_);
  nor (_40161_, _40160_, _39845_);
  or (_40162_, _40161_, _40153_);
  or (_40163_, _40162_, _39841_);
  and (_40164_, _40163_, _42882_);
  and (_41612_, _40164_, _40152_);
  nand (_40165_, _39845_, _38464_);
  not (_40166_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_40167_, _39882_, _39848_);
  nor (_40168_, _39884_, _39846_);
  not (_40169_, _40168_);
  and (_40170_, _40169_, _40167_);
  nor (_40171_, _40170_, _40166_);
  and (_40172_, _40170_, _40166_);
  or (_40173_, _40172_, _40171_);
  or (_40174_, _40173_, _39845_);
  and (_40175_, _40174_, _40165_);
  or (_40176_, _40175_, _39896_);
  nand (_40177_, _39896_, _40166_);
  and (_40178_, _40177_, _42882_);
  and (_41614_, _40178_, _40176_);
  not (_40179_, _39852_);
  nor (_40180_, _39885_, _40179_);
  not (_40181_, _40180_);
  nor (_40182_, _40167_, _39852_);
  nor (_40183_, _40182_, _40166_);
  and (_40184_, _40183_, _40181_);
  or (_40185_, _40184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_40186_, _40184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_40187_, _40186_, _40185_);
  or (_40188_, _40187_, _39845_);
  nand (_40189_, _39845_, _38456_);
  and (_40190_, _40189_, _40188_);
  or (_40191_, _40190_, _39896_);
  or (_40192_, _39897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_40193_, _40192_, _42882_);
  and (_41616_, _40193_, _40191_);
  nand (_40194_, _39845_, _38449_);
  and (_40195_, _39912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_40196_, _40195_, _39882_);
  and (_40197_, _40196_, _39848_);
  nand (_40198_, _40197_, _40169_);
  and (_40199_, _40198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_40200_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_40201_, _40200_);
  not (_40202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_40203_, _39912_, _40202_);
  and (_40204_, _40203_, _39882_);
  and (_40205_, _40204_, _40201_);
  or (_40206_, _40205_, _40199_);
  or (_40207_, _40206_, _39845_);
  and (_40208_, _40207_, _40194_);
  or (_40209_, _40208_, _39896_);
  nand (_40210_, _39896_, _40202_);
  and (_40211_, _40210_, _42882_);
  and (_41618_, _40211_, _40209_);
  nand (_40212_, _39845_, _38442_);
  nor (_40213_, _39904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_40214_, _40196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_40215_, _40214_, _39884_);
  nor (_40216_, _40215_, _40213_);
  or (_40217_, _40216_, _40179_);
  not (_40218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_40219_, _40197_, _40218_);
  nor (_40220_, _40197_, _40218_);
  or (_40221_, _40220_, _39852_);
  or (_40222_, _40221_, _40219_);
  and (_40223_, _40222_, _40217_);
  or (_40224_, _40223_, _39845_);
  and (_40225_, _40224_, _40212_);
  or (_40226_, _40225_, _39896_);
  nand (_40227_, _39896_, _40218_);
  and (_40228_, _40227_, _42882_);
  and (_41620_, _40228_, _40226_);
  nand (_40229_, _39845_, _38434_);
  and (_40230_, _39904_, _39898_);
  or (_40231_, _40215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_40232_, _40231_, _39852_);
  nor (_40233_, _40232_, _40230_);
  and (_40234_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_40235_, _40234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not (_40237_, _39919_);
  and (_40238_, _40214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_40239_, _40238_, _40237_);
  or (_40240_, _40239_, _40236_);
  and (_40241_, _40240_, _40235_);
  or (_40242_, _40241_, _40233_);
  nor (_40243_, _40242_, _39845_);
  nor (_40244_, _40243_, _39841_);
  and (_40245_, _40244_, _40229_);
  and (_40246_, _39896_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_40247_, _40246_, _40245_);
  and (_41622_, _40247_, _42882_);
  nand (_40248_, _39845_, _38428_);
  and (_40249_, _40230_, _39848_);
  nor (_40250_, _40249_, _39919_);
  nor (_40251_, _40250_, _40239_);
  nand (_40252_, _40251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_40253_, _40251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_40254_, _40253_, _40252_);
  or (_40255_, _40254_, _39845_);
  and (_40256_, _40255_, _40248_);
  or (_40257_, _40256_, _39896_);
  or (_40258_, _39897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_40259_, _40258_, _42882_);
  and (_41623_, _40259_, _40257_);
  nand (_40260_, _39845_, _38420_);
  and (_40261_, _40238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_40262_, _40201_, _40261_);
  or (_40263_, _40262_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_40264_, _40262_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40265_, _40264_, _40263_);
  nor (_40266_, _40265_, _39845_);
  nor (_40267_, _40266_, _39841_);
  and (_40268_, _40267_, _40260_);
  and (_40269_, _39896_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_40270_, _40269_, _40268_);
  and (_41625_, _40270_, _42882_);
  nor (_40271_, _39986_, _39955_);
  or (_40272_, _40271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_40273_, _39977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_40274_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40275_, _40274_, _40024_);
  nand (_40276_, _40275_, _40273_);
  or (_40277_, _40276_, _39955_);
  and (_40278_, _40277_, _40272_);
  or (_40279_, _40278_, _39994_);
  nand (_40280_, _39994_, _38464_);
  and (_40281_, _40280_, _42882_);
  and (_41627_, _40281_, _40279_);
  nand (_40282_, _39994_, _38456_);
  and (_40283_, _39955_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_40284_, _40273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_40285_, _40273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_40286_, _40285_, _40284_);
  and (_40287_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40288_, _40287_, _39983_);
  nor (_40289_, _40288_, _40286_);
  nor (_40290_, _40289_, _39955_);
  or (_40291_, _40290_, _40283_);
  or (_40292_, _40291_, _39994_);
  and (_40293_, _40292_, _42882_);
  and (_41629_, _40293_, _40282_);
  not (_40294_, _39996_);
  nor (_40295_, _40285_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_40296_, _40273_, _39978_);
  nor (_40297_, _40296_, _40295_);
  and (_40298_, _40005_, _39983_);
  and (_40299_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_40300_, _40299_, _40297_);
  nor (_40301_, _40300_, _39955_);
  and (_40302_, _39955_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_40303_, _40302_, _40301_);
  and (_40304_, _40303_, _40294_);
  nor (_40305_, _40020_, _38449_);
  or (_40306_, _40305_, _40304_);
  and (_41631_, _40306_, _42882_);
  and (_40307_, _39980_, _39977_);
  nor (_40308_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_40309_, _40308_, _40307_);
  and (_40310_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_40311_, _40310_, _40309_);
  nor (_40312_, _40311_, _39955_);
  and (_40313_, _39955_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_40314_, _40313_, _40312_);
  and (_40315_, _40314_, _40294_);
  nor (_40316_, _40020_, _38442_);
  or (_40317_, _40316_, _40315_);
  and (_41633_, _40317_, _42882_);
  nand (_40318_, _39994_, _38434_);
  or (_40319_, _39998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_40320_, _40307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_40321_, _40320_, _39982_);
  and (_40322_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_40323_, _40322_, _40321_);
  or (_40324_, _40323_, _39955_);
  and (_40325_, _40324_, _40319_);
  or (_40326_, _40325_, _39994_);
  and (_40327_, _40326_, _42882_);
  and (_41635_, _40327_, _40318_);
  nand (_40328_, _39994_, _38428_);
  not (_40329_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_40330_, _39982_, _39966_);
  and (_40331_, _40330_, _40329_);
  and (_40332_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_40333_, _40332_, _40331_);
  nor (_40334_, _40333_, _39955_);
  and (_40335_, _40330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_40336_, _40335_);
  or (_40337_, _40336_, _39955_);
  and (_40338_, _40337_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_40339_, _40338_, _40334_);
  or (_40340_, _40339_, _39994_);
  and (_40341_, _40340_, _42882_);
  and (_41637_, _40341_, _40328_);
  and (_40342_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_40343_, _40342_, _39977_);
  and (_40344_, _40343_, _40024_);
  nor (_40345_, _40336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_40346_, _40345_, _40344_);
  nor (_40347_, _40346_, _39955_);
  and (_40348_, _40337_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_40349_, _40348_, _40347_);
  and (_40350_, _40349_, _40294_);
  nor (_40351_, _40020_, _38420_);
  or (_40352_, _40351_, _40350_);
  and (_41638_, _40352_, _42882_);
  or (_40353_, _40026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40354_, _40353_, _40022_);
  and (_40355_, _40026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_40356_, _40355_, _40354_);
  and (_40357_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_40358_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40359_, _40358_, _40033_);
  nor (_40360_, _40359_, _40357_);
  and (_40361_, _39982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_40362_, _39982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40363_, _40362_, _39965_);
  nor (_40364_, _40363_, _40361_);
  or (_40365_, _40364_, _40360_);
  or (_40366_, _40365_, _40356_);
  or (_40367_, _40366_, _39955_);
  nand (_40368_, _39955_, _38464_);
  and (_40369_, _40368_, _40367_);
  and (_40370_, _40369_, _40066_);
  and (_40371_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_40372_, _40371_, _40370_);
  and (_41640_, _40372_, _42882_);
  nand (_40373_, _39955_, _38456_);
  or (_40374_, _40355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40375_, _40024_, _39977_);
  and (_40376_, _40375_, _39958_);
  not (_40377_, _40376_);
  or (_40378_, _40377_, _40005_);
  and (_40379_, _40378_, _40022_);
  and (_40380_, _40379_, _40374_);
  and (_40381_, _40034_, _39958_);
  or (_40382_, _40357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_40383_, _40382_, _40033_);
  nor (_40384_, _40383_, _40381_);
  and (_40385_, _40361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_40386_, _40361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_40387_, _40386_, _39965_);
  nor (_40388_, _40387_, _40385_);
  or (_40389_, _40388_, _40384_);
  or (_40390_, _40389_, _40380_);
  or (_40391_, _40390_, _39955_);
  and (_40392_, _40391_, _40020_);
  and (_40393_, _40392_, _40373_);
  and (_40394_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_40395_, _40394_, _40393_);
  and (_41642_, _40395_, _42882_);
  nor (_40396_, _39998_, _38449_);
  or (_40397_, _40376_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40398_, _40375_, _39959_);
  not (_40399_, _40398_);
  and (_40400_, _40399_, _40021_);
  and (_40401_, _40400_, _40397_);
  and (_40402_, _39977_, _39958_);
  and (_40403_, _40402_, _39981_);
  or (_40404_, _40403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40405_, _39982_, _39959_);
  nor (_40406_, _40405_, _39966_);
  and (_40407_, _40406_, _40404_);
  and (_40408_, _40381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_40409_, _40408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40410_, _40034_, _39959_);
  nand (_40411_, _40410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40412_, _40411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40413_, _40412_, _40409_);
  or (_40414_, _40413_, _40407_);
  nor (_40415_, _40414_, _40401_);
  nor (_40416_, _40415_, _39955_);
  or (_40417_, _40416_, _39996_);
  or (_40418_, _40417_, _40396_);
  or (_40419_, _40294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40420_, _40419_, _42882_);
  and (_41644_, _40420_, _40418_);
  nor (_40421_, _39998_, _38442_);
  not (_40422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40423_, _40398_, _40004_);
  nor (_40424_, _40423_, _40422_);
  and (_40425_, _40423_, _40422_);
  or (_40426_, _40425_, _40424_);
  and (_40427_, _40426_, _40022_);
  or (_40428_, _40410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_40429_, _40035_);
  and (_40430_, _40429_, _40033_);
  and (_40431_, _40430_, _40428_);
  or (_40432_, _40405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40433_, _39982_, _39960_);
  nor (_40434_, _40433_, _39966_);
  and (_40435_, _40434_, _40432_);
  or (_40436_, _40435_, _40431_);
  nor (_40437_, _40436_, _40427_);
  nor (_40438_, _40437_, _39955_);
  or (_40439_, _40438_, _39996_);
  or (_40440_, _40439_, _40421_);
  nand (_40441_, _39996_, _40422_);
  and (_40442_, _40441_, _42882_);
  and (_41646_, _40442_, _40440_);
  nand (_40443_, _39955_, _38434_);
  or (_40444_, _40433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40445_, _40403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40446_, _40445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40447_, _40446_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_40448_, _40447_, _39966_);
  and (_40449_, _40448_, _40444_);
  and (_40450_, _40375_, _39960_);
  nand (_40451_, _40450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_40452_, _40450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40453_, _40452_, _40021_);
  and (_40454_, _40453_, _40451_);
  and (_40455_, _40035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_40456_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40457_, _40456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40458_, _40035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_40459_, _40458_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40460_, _40459_, _40457_);
  or (_40461_, _40460_, _40454_);
  or (_40462_, _40461_, _40449_);
  or (_40463_, _40462_, _39955_);
  and (_40464_, _40463_, _40020_);
  and (_40465_, _40464_, _40443_);
  and (_40466_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_40467_, _40466_, _40465_);
  and (_41648_, _40467_, _42882_);
  nor (_40468_, _39998_, _38428_);
  not (_40469_, _40447_);
  nor (_40470_, _40469_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40471_, _40469_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_40472_, _40471_, _40470_);
  and (_40473_, _40472_, _39965_);
  nor (_40474_, _40451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_40475_, _40474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_40476_, _40474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40477_, _40476_, _40022_);
  and (_40478_, _40477_, _40475_);
  not (_40479_, _40038_);
  and (_40480_, _40479_, _40033_);
  or (_40481_, _40458_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40482_, _40481_, _40480_);
  or (_40483_, _40482_, _40478_);
  nor (_40484_, _40483_, _40473_);
  nor (_40485_, _40484_, _39955_);
  or (_40486_, _40485_, _39996_);
  or (_40487_, _40486_, _40468_);
  or (_40488_, _40294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40489_, _40488_, _42882_);
  and (_41650_, _40489_, _40487_);
  nand (_40490_, _39955_, _38420_);
  or (_40491_, _40027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_40492_, _40491_, _40022_);
  nor (_40493_, _40492_, _40028_);
  or (_40494_, _40038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_40495_, _40046_);
  and (_40496_, _40495_, _40033_);
  and (_40497_, _40496_, _40494_);
  or (_40498_, _39988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_40499_, _40051_, _39966_);
  and (_40500_, _40499_, _40498_);
  or (_40501_, _40500_, _40497_);
  or (_40502_, _40501_, _40493_);
  or (_40503_, _40502_, _39955_);
  and (_40504_, _40503_, _40020_);
  and (_40505_, _40504_, _40490_);
  and (_40506_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40507_, _40506_, _40505_);
  and (_41652_, _40507_, _42882_);
  nand (_40508_, _40074_, _38464_);
  or (_40509_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40510_, _40509_, _42882_);
  and (_41653_, _40510_, _40508_);
  or (_40511_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40512_, _40511_, _42882_);
  nand (_40513_, _40074_, _38456_);
  and (_41655_, _40513_, _40512_);
  or (_40514_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_40515_, _40514_, _42882_);
  nand (_40516_, _40074_, _38449_);
  and (_41657_, _40516_, _40515_);
  or (_40517_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_40518_, _40517_, _42882_);
  nand (_40519_, _40074_, _38442_);
  and (_41659_, _40519_, _40518_);
  or (_40520_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_40521_, _40520_, _42882_);
  nand (_40522_, _40074_, _38434_);
  and (_41660_, _40522_, _40521_);
  or (_40523_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_40524_, _40523_, _42882_);
  nand (_40525_, _40074_, _38428_);
  and (_41662_, _40525_, _40524_);
  or (_40526_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_40527_, _40526_, _42882_);
  nand (_40528_, _40074_, _38420_);
  and (_41664_, _40528_, _40527_);
  nor (_40529_, _27845_, _27703_);
  and (_40530_, _40529_, _39031_);
  and (_40531_, _40530_, _39236_);
  and (_40532_, _40531_, _31304_);
  nand (_40533_, _40532_, _31282_);
  and (_40534_, _38401_, _31304_);
  and (_40535_, _40534_, _39260_);
  not (_40536_, _40535_);
  or (_40537_, _40532_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_40538_, _40537_, _40536_);
  and (_40539_, _40538_, _40533_);
  nor (_40540_, _40536_, _38485_);
  or (_40541_, _40540_, _40539_);
  and (_42827_, _40541_, _42882_);
  and (_40542_, _39839_, _27045_);
  and (_40543_, _40542_, _39243_);
  not (_40544_, _40543_);
  and (_40545_, _27845_, _27714_);
  and (_40546_, _40545_, _39031_);
  and (_40547_, _40546_, _39236_);
  and (_40548_, _40547_, _31304_);
  or (_40549_, _40548_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_40550_, _40549_, _40544_);
  nand (_40551_, _40548_, _31282_);
  and (_40552_, _40551_, _40550_);
  nor (_40553_, _40544_, _38485_);
  or (_40554_, _40553_, _40552_);
  and (_42830_, _40554_, _42882_);
  and (_40555_, _40542_, _38405_);
  nor (_40556_, _39030_, _27703_);
  and (_40557_, _40556_, _27845_);
  and (_40558_, _40557_, _27560_);
  and (_40559_, _40558_, _39205_);
  nand (_40560_, _40559_, _27023_);
  and (_40561_, _40560_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40562_, _40561_, _40555_);
  or (_40563_, _27034_, _33285_);
  and (_40564_, _40563_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40565_, _40564_, _39007_);
  and (_40566_, _40565_, _40559_);
  or (_40567_, _40566_, _40562_);
  nand (_40568_, _40555_, _38420_);
  and (_40569_, _40568_, _42882_);
  and (_42832_, _40569_, _40567_);
  not (_40570_, _40555_);
  nor (_40571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_40572_, _40571_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not (_40573_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_40574_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_40575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40576_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40575_);
  and (_40577_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40578_, _40577_, _40576_);
  nor (_40579_, _40578_, _40574_);
  or (_40580_, _40579_, _40573_);
  and (_40581_, _40575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_40582_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_40583_, _40582_, _40581_);
  nor (_40584_, _40583_, _40574_);
  and (_40585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40575_);
  and (_40586_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40587_, _40586_, _40585_);
  nand (_40588_, _40587_, _40584_);
  or (_40590_, _40588_, _40580_);
  and (_40592_, _40590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_40594_, _40592_, _40572_);
  and (_40596_, _38405_, _31304_);
  and (_40598_, _40596_, _40556_);
  or (_40600_, _40598_, _40594_);
  and (_40602_, _40600_, _40570_);
  nand (_40604_, _40598_, _31282_);
  and (_40606_, _40604_, _40602_);
  nor (_40608_, _40570_, _38485_);
  or (_40610_, _40608_, _40606_);
  and (_42834_, _40610_, _42882_);
  and (_40613_, _39844_, _31348_);
  nand (_40615_, _40613_, _31282_);
  not (_40617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_40619_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_40621_, _40587_, _40574_);
  not (_40623_, _40621_);
  or (_40625_, _40623_, _40584_);
  or (_40627_, _40625_, _40580_);
  and (_40629_, _40627_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_40631_, _40629_, _40619_);
  or (_40633_, _40631_, _40613_);
  and (_40635_, _40633_, _40570_);
  and (_40637_, _40635_, _40615_);
  nor (_40639_, _40570_, _38428_);
  or (_40641_, _40639_, _40637_);
  and (_42836_, _40641_, _42882_);
  not (_40643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_40644_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _40643_);
  nand (_40645_, _40579_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_40646_, _40621_, _40584_);
  or (_40647_, _40646_, _40645_);
  and (_40648_, _40647_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_40649_, _40648_, _40644_);
  and (_40650_, _40073_, _31348_);
  or (_40651_, _40650_, _40649_);
  and (_40652_, _40651_, _40570_);
  nand (_40653_, _40650_, _31282_);
  and (_40654_, _40653_, _40652_);
  nor (_40655_, _40570_, _38456_);
  or (_40656_, _40655_, _40654_);
  and (_42838_, _40656_, _42882_);
  and (_40657_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_40658_, _40645_, _40625_);
  and (_40659_, _40658_, _40657_);
  and (_40660_, _40556_, _38623_);
  or (_40661_, _40660_, _40659_);
  and (_40662_, _40661_, _40570_);
  nand (_40663_, _40660_, _31282_);
  and (_40664_, _40663_, _40662_);
  nor (_40665_, _40570_, _38442_);
  or (_40666_, _40665_, _40664_);
  and (_42840_, _40666_, _42882_);
  and (_40667_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40668_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40575_);
  nor (_40669_, _40668_, _40667_);
  and (_40670_, _40669_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_40671_, _40670_, _40574_);
  and (_40672_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40673_, _40672_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_40674_, _40673_);
  and (_40675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40676_, _40675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_40677_, _40676_);
  and (_40678_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40679_, _40678_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40680_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_40681_, _40680_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_40682_, _40681_, _40679_);
  and (_40683_, _40682_, _40677_);
  and (_40684_, _40683_, _40674_);
  not (_40685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_40686_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_40687_, _40686_, _40685_);
  nand (_40688_, _40687_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_40689_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_40690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_40691_, _40690_, _40689_);
  and (_40692_, _40691_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_40693_, _40692_);
  and (_40694_, _40693_, _40688_);
  and (_40695_, _40694_, _40684_);
  nor (_40696_, _40695_, _40671_);
  and (_40697_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_40698_, _40697_, _40575_);
  and (_40699_, _40698_, _40696_);
  not (_40700_, _40699_);
  not (_40701_, _40698_);
  and (_40702_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _40574_);
  not (_40703_, _40702_);
  not (_40704_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40705_, _40675_, _40704_);
  not (_40706_, _40705_);
  not (_40707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40708_, _40678_, _40707_);
  not (_40709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_40710_, _40680_, _40709_);
  nor (_40711_, _40710_, _40708_);
  and (_40712_, _40711_, _40706_);
  nor (_40713_, _40712_, _40703_);
  not (_40714_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40715_, _40687_, _40714_);
  not (_40716_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40717_, _40691_, _40716_);
  nor (_40718_, _40717_, _40715_);
  not (_40719_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40720_, _40672_, _40719_);
  not (_40721_, _40720_);
  and (_40722_, _40721_, _40718_);
  nor (_40723_, _40722_, _40703_);
  nor (_40724_, _40723_, _40713_);
  or (_40725_, _40724_, _40701_);
  and (_40726_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42882_);
  and (_40727_, _40726_, _40725_);
  and (_42870_, _40727_, _40700_);
  nor (_40728_, _40697_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40729_, _40728_);
  not (_40730_, _40696_);
  and (_40731_, _40724_, _40730_);
  nor (_40732_, _40731_, _40729_);
  nand (_40733_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42882_);
  nor (_42872_, _40733_, _40732_);
  and (_40734_, _40694_, _40674_);
  nand (_40735_, _40734_, _40696_);
  or (_40736_, _40723_, _40696_);
  and (_40737_, _40736_, _40698_);
  and (_40738_, _40737_, _40735_);
  or (_40739_, _40738_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_40740_, _40700_, _40683_);
  nor (_40741_, _40701_, _40696_);
  nand (_40742_, _40741_, _40713_);
  and (_40743_, _40742_, _42882_);
  and (_40744_, _40743_, _40740_);
  and (_42873_, _40744_, _40739_);
  and (_40745_, _40735_, _40728_);
  or (_40746_, _40745_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40747_, _40728_, _40696_);
  not (_40748_, _40747_);
  or (_40749_, _40748_, _40683_);
  or (_40750_, _40723_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand (_40754_, _40728_, _40713_);
  and (_40755_, _40754_, _40750_);
  or (_40761_, _40755_, _40696_);
  and (_40767_, _40761_, _42882_);
  and (_40773_, _40767_, _40749_);
  and (_42875_, _40773_, _40746_);
  nand (_40779_, _40731_, _40574_);
  nor (_40780_, _40575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_40781_, _40780_, _40697_);
  and (_40782_, _40781_, _42882_);
  and (_42877_, _40782_, _40779_);
  and (_40783_, _40731_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_40784_, _40575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_40785_, _40784_, _40780_);
  nor (_40786_, _40785_, _40730_);
  or (_40787_, _40786_, _40697_);
  or (_40788_, _40787_, _40783_);
  not (_40789_, _40697_);
  or (_40790_, _40785_, _40789_);
  and (_40791_, _40790_, _42882_);
  and (_42879_, _40791_, _40788_);
  and (_40796_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42882_);
  and (_42880_, _40796_, _40697_);
  nor (_42885_, _40571_, rst);
  and (_42886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _42882_);
  nor (_40804_, _40731_, _40697_);
  and (_40810_, _40697_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_40811_, _40810_, _40804_);
  and (_00130_, _40811_, _42882_);
  and (_40812_, _40697_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_40817_, _40812_, _40804_);
  and (_00132_, _40817_, _42882_);
  and (_40822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42882_);
  and (_00134_, _40822_, _40697_);
  not (_40826_, _40710_);
  nor (_40832_, _40717_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_40833_, _40832_, _40715_);
  or (_40834_, _40833_, _40720_);
  and (_40839_, _40834_, _40826_);
  or (_40840_, _40839_, _40708_);
  nor (_40845_, _40724_, _40696_);
  and (_40846_, _40845_, _40706_);
  and (_40847_, _40846_, _40840_);
  not (_40852_, _40681_);
  or (_40857_, _40692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40858_, _40857_, _40688_);
  or (_40859_, _40858_, _40673_);
  and (_40868_, _40859_, _40852_);
  or (_40869_, _40868_, _40679_);
  and (_40870_, _40696_, _40677_);
  and (_40871_, _40870_, _40869_);
  or (_40875_, _40871_, _40697_);
  or (_40881_, _40875_, _40847_);
  or (_40882_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40883_, _40882_, _42882_);
  and (_00136_, _40883_, _40881_);
  not (_40888_, _40679_);
  or (_40893_, _40681_, _40673_);
  and (_40894_, _40694_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_40895_, _40894_, _40893_);
  and (_40900_, _40895_, _40888_);
  and (_40905_, _40900_, _40870_);
  nor (_40906_, _40708_, _40705_);
  or (_40907_, _40720_, _40710_);
  and (_40911_, _40718_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_40917_, _40911_, _40907_);
  and (_40918_, _40917_, _40906_);
  and (_40922_, _40918_, _40845_);
  or (_40923_, _40922_, _40697_);
  or (_40929_, _40923_, _40905_);
  or (_40930_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_40931_, _40930_, _42882_);
  and (_00138_, _40931_, _40929_);
  and (_40938_, _40721_, _40702_);
  nand (_40941_, _40938_, _40712_);
  nor (_40942_, _40941_, _40718_);
  nor (_40944_, _40694_, _40671_);
  or (_40950_, _40944_, _40942_);
  or (_40953_, _40684_, _40671_);
  and (_40954_, _40953_, _40950_);
  or (_40955_, _40954_, _40697_);
  or (_40961_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_40965_, _40961_, _42882_);
  and (_00140_, _40965_, _40955_);
  and (_40966_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42882_);
  and (_00141_, _40966_, _40697_);
  and (_40974_, _40697_, _40575_);
  or (_40975_, _40974_, _40732_);
  or (_40976_, _40975_, _40741_);
  and (_00143_, _40976_, _42882_);
  not (_40977_, _40804_);
  and (_40978_, _40977_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_40979_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_40980_, _40692_, _40575_);
  or (_40981_, _40980_, _40979_);
  nor (_40982_, _40688_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40983_, _40982_, _40673_);
  nand (_40984_, _40983_, _40981_);
  or (_40985_, _40674_, _40577_);
  and (_40986_, _40985_, _40984_);
  or (_40987_, _40986_, _40681_);
  or (_40988_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40575_);
  or (_40989_, _40988_, _40852_);
  and (_40990_, _40989_, _40888_);
  and (_40991_, _40990_, _40987_);
  and (_40992_, _40679_, _40577_);
  or (_40993_, _40992_, _40676_);
  or (_40994_, _40993_, _40991_);
  or (_40995_, _40988_, _40677_);
  and (_40996_, _40995_, _40696_);
  and (_40997_, _40996_, _40994_);
  and (_40998_, _40717_, _40575_);
  or (_40999_, _40998_, _40979_);
  and (_41000_, _40715_, _40575_);
  nor (_41001_, _41000_, _40720_);
  nand (_41002_, _41001_, _40999_);
  or (_41003_, _40721_, _40577_);
  and (_41004_, _41003_, _41002_);
  or (_41005_, _41004_, _40710_);
  not (_41006_, _40708_);
  or (_41007_, _40988_, _40826_);
  and (_41008_, _41007_, _41006_);
  and (_41009_, _41008_, _41005_);
  and (_41010_, _40708_, _40577_);
  or (_41011_, _41010_, _40705_);
  or (_41012_, _41011_, _41009_);
  and (_41013_, _40988_, _40845_);
  or (_41014_, _41013_, _40846_);
  and (_41015_, _41014_, _41012_);
  or (_41016_, _41015_, _40997_);
  and (_41017_, _41016_, _40789_);
  or (_41018_, _41017_, _40978_);
  and (_00145_, _41018_, _42882_);
  and (_41019_, _40977_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_41020_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40575_);
  and (_41021_, _41020_, _40677_);
  or (_41022_, _41021_, _40683_);
  or (_41023_, _40980_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_41024_, _41023_, _40983_);
  nand (_41025_, _40673_, _40586_);
  nand (_41026_, _41025_, _40682_);
  or (_41027_, _41026_, _41024_);
  and (_41028_, _41027_, _41022_);
  and (_41029_, _40676_, _40586_);
  or (_41030_, _41029_, _41028_);
  and (_41031_, _41030_, _40696_);
  and (_41032_, _40705_, _40586_);
  and (_41033_, _41020_, _40706_);
  or (_41034_, _41033_, _40712_);
  and (_41035_, _40720_, _40586_);
  not (_41036_, _40711_);
  or (_41037_, _40998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_41038_, _41037_, _41001_);
  or (_41039_, _41038_, _41036_);
  or (_41040_, _41039_, _41035_);
  and (_41041_, _41040_, _41034_);
  or (_41042_, _41041_, _41032_);
  and (_41043_, _41042_, _40845_);
  or (_41044_, _41043_, _41031_);
  and (_41045_, _41044_, _40789_);
  or (_41046_, _41045_, _41019_);
  and (_00147_, _41046_, _42882_);
  and (_41047_, _40977_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_41048_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_41049_, _41048_, _40677_);
  and (_41050_, _41049_, _40696_);
  not (_41051_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_41052_, _40692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_41053_, _41052_, _41051_);
  nor (_41054_, _40688_, _40575_);
  nor (_41055_, _41054_, _40673_);
  nand (_41056_, _41055_, _41053_);
  or (_41057_, _40674_, _40576_);
  and (_41058_, _41057_, _41056_);
  or (_41059_, _41058_, _40681_);
  or (_41060_, _41048_, _40852_);
  and (_41061_, _41060_, _40888_);
  and (_41062_, _41061_, _41059_);
  and (_41063_, _40679_, _40576_);
  or (_41064_, _41063_, _40676_);
  or (_41065_, _41064_, _41062_);
  and (_41066_, _41065_, _41050_);
  or (_41067_, _41048_, _40706_);
  and (_41068_, _40717_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_41069_, _41068_, _41051_);
  and (_41070_, _40715_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_41071_, _41070_, _40720_);
  nand (_41072_, _41071_, _41069_);
  or (_41073_, _40721_, _40576_);
  and (_41074_, _41073_, _41072_);
  or (_41075_, _41074_, _40710_);
  or (_41076_, _41048_, _40826_);
  and (_41077_, _41076_, _41006_);
  and (_41078_, _41077_, _41075_);
  and (_41079_, _40708_, _40576_);
  or (_41080_, _41079_, _40705_);
  or (_41081_, _41080_, _41078_);
  and (_41082_, _41081_, _40845_);
  and (_41083_, _41082_, _41067_);
  or (_41084_, _41083_, _41066_);
  and (_41085_, _41084_, _40789_);
  or (_41086_, _41085_, _41047_);
  and (_00149_, _41086_, _42882_);
  and (_41087_, _40977_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_41088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_41089_, _41088_, _40677_);
  or (_41090_, _41089_, _40683_);
  or (_41091_, _41052_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_41093_, _41091_, _41055_);
  nand (_41094_, _40673_, _40585_);
  nand (_41096_, _41094_, _40682_);
  or (_41097_, _41096_, _41093_);
  and (_41099_, _41097_, _41090_);
  and (_41100_, _40676_, _40585_);
  or (_41102_, _41100_, _41099_);
  and (_41103_, _41102_, _40696_);
  and (_41105_, _40705_, _40585_);
  and (_41106_, _41088_, _40706_);
  or (_41108_, _41106_, _40712_);
  and (_41109_, _40720_, _40585_);
  or (_41111_, _41068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_41112_, _41111_, _41071_);
  or (_41114_, _41112_, _41036_);
  or (_41115_, _41114_, _41109_);
  and (_41117_, _41115_, _41108_);
  or (_41118_, _41117_, _41105_);
  and (_41120_, _41118_, _40845_);
  or (_41121_, _41120_, _41103_);
  and (_41122_, _41121_, _40789_);
  or (_41123_, _41122_, _41087_);
  and (_00151_, _41123_, _42882_);
  or (_41124_, _40729_, _40724_);
  and (_41125_, _41124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_41126_, _41125_, _40747_);
  and (_00152_, _41126_, _42882_);
  and (_41127_, _40725_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_41128_, _41127_, _40699_);
  and (_00154_, _41128_, _42882_);
  and (_41129_, _40559_, _27045_);
  or (_41130_, _41129_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_41131_, _41130_, _40570_);
  nand (_41132_, _41129_, _31282_);
  and (_41133_, _41132_, _41131_);
  and (_41134_, _40555_, _38465_);
  or (_41135_, _41134_, _41133_);
  and (_00156_, _41135_, _42882_);
  and (_41136_, _40559_, _33296_);
  or (_41137_, _41136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_41138_, _41137_, _40570_);
  nand (_41139_, _41136_, _31282_);
  and (_41140_, _41139_, _41138_);
  nor (_41141_, _40570_, _38449_);
  or (_41142_, _41141_, _41140_);
  and (_00158_, _41142_, _42882_);
  and (_41143_, _40559_, _34765_);
  or (_41144_, _41143_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_41145_, _41144_, _40570_);
  nand (_41146_, _41143_, _31282_);
  and (_41147_, _41146_, _41145_);
  nor (_41148_, _40570_, _38434_);
  or (_41149_, _41148_, _41147_);
  and (_00160_, _41149_, _42882_);
  and (_41150_, _40547_, _27045_);
  or (_41151_, _41150_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_41152_, _41151_, _40544_);
  nand (_41153_, _41150_, _31282_);
  and (_41154_, _41153_, _41152_);
  and (_41155_, _40543_, _38465_);
  or (_41156_, _41155_, _41154_);
  and (_00162_, _41156_, _42882_);
  and (_41157_, _40547_, _32567_);
  or (_41158_, _41157_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_41159_, _41158_, _40544_);
  nand (_41160_, _41157_, _31282_);
  and (_41161_, _41160_, _41159_);
  nor (_41162_, _40544_, _38456_);
  or (_41163_, _41162_, _41161_);
  and (_00163_, _41163_, _42882_);
  nand (_41164_, _40547_, _39293_);
  and (_41165_, _41164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_41166_, _41165_, _40543_);
  and (_41167_, _33329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_41168_, _41167_, _33318_);
  and (_41169_, _41168_, _40547_);
  or (_41170_, _41169_, _41166_);
  nand (_41171_, _40543_, _38449_);
  and (_41172_, _41171_, _42882_);
  and (_00165_, _41172_, _41170_);
  and (_41173_, _40547_, _34004_);
  or (_41174_, _41173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_41175_, _41174_, _40544_);
  nand (_41176_, _41173_, _31282_);
  and (_41177_, _41176_, _41175_);
  nor (_41178_, _40544_, _38442_);
  or (_41179_, _41178_, _41177_);
  and (_00167_, _41179_, _42882_);
  and (_41180_, _40547_, _34765_);
  or (_41181_, _41180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_41182_, _41181_, _40544_);
  nand (_41183_, _41180_, _31282_);
  and (_41184_, _41183_, _41182_);
  nor (_41185_, _40544_, _38434_);
  or (_41186_, _41185_, _41184_);
  and (_00169_, _41186_, _42882_);
  and (_41187_, _40547_, _35549_);
  or (_41188_, _41187_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_41189_, _41188_, _40544_);
  nand (_41190_, _41187_, _31282_);
  and (_41191_, _41190_, _41189_);
  nor (_41192_, _40544_, _38428_);
  or (_41193_, _41192_, _41191_);
  and (_00171_, _41193_, _42882_);
  and (_41194_, _40547_, _36277_);
  or (_41195_, _41194_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_41196_, _41195_, _40544_);
  nand (_41197_, _41194_, _31282_);
  and (_41198_, _41197_, _41196_);
  nor (_41199_, _40544_, _38420_);
  or (_41200_, _41199_, _41198_);
  and (_00173_, _41200_, _42882_);
  and (_41201_, _40531_, _27045_);
  nand (_41202_, _41201_, _31282_);
  or (_41203_, _41201_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_41204_, _41203_, _40536_);
  and (_41205_, _41204_, _41202_);
  and (_41206_, _40535_, _38465_);
  or (_41207_, _41206_, _41205_);
  and (_00174_, _41207_, _42882_);
  and (_41208_, _40531_, _32567_);
  nand (_41209_, _41208_, _31282_);
  or (_41210_, _41208_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_41211_, _41210_, _40536_);
  and (_41212_, _41211_, _41209_);
  nor (_41213_, _40536_, _38456_);
  or (_41214_, _41213_, _41212_);
  and (_00176_, _41214_, _42882_);
  and (_41215_, _33329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_41216_, _41215_, _33318_);
  and (_41217_, _41216_, _40531_);
  nand (_41218_, _40531_, _39293_);
  and (_41219_, _41218_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_41220_, _41219_, _40535_);
  or (_41221_, _41220_, _41217_);
  nand (_41222_, _40535_, _38449_);
  and (_41223_, _41222_, _42882_);
  and (_00178_, _41223_, _41221_);
  and (_41224_, _40531_, _34004_);
  nand (_41225_, _41224_, _31282_);
  or (_41226_, _41224_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_41227_, _41226_, _41225_);
  or (_41228_, _41227_, _40535_);
  nand (_41229_, _40535_, _38442_);
  and (_41230_, _41229_, _42882_);
  and (_00180_, _41230_, _41228_);
  and (_41231_, _40531_, _34765_);
  nand (_41232_, _41231_, _31282_);
  or (_41233_, _41231_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_41234_, _41233_, _40536_);
  and (_41235_, _41234_, _41232_);
  nor (_41236_, _40536_, _38434_);
  or (_41237_, _41236_, _41235_);
  and (_00182_, _41237_, _42882_);
  and (_41238_, _40531_, _35549_);
  nand (_41239_, _41238_, _31282_);
  or (_41240_, _41238_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_41241_, _41240_, _41239_);
  or (_41242_, _41241_, _40535_);
  nand (_41243_, _40535_, _38428_);
  and (_41244_, _41243_, _42882_);
  and (_00184_, _41244_, _41242_);
  and (_41245_, _40531_, _36277_);
  nand (_41246_, _41245_, _31282_);
  or (_41247_, _41245_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_41248_, _41247_, _41246_);
  or (_41249_, _41248_, _40535_);
  nand (_41250_, _40535_, _38420_);
  and (_41251_, _41250_, _42882_);
  and (_00185_, _41251_, _41249_);
  and (_41252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_41253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_41254_, _40571_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_41255_, _41254_, _41253_);
  not (_41256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_41257_, _41256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_41258_, _41257_, _41255_);
  nor (_41259_, _41258_, _41252_);
  or (_41260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_41261_, _41260_, _42882_);
  nor (_00546_, _41261_, _41259_);
  nor (_41262_, _41259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_41263_, _41262_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_41264_, _41262_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_41265_, _41264_, _42882_);
  and (_00548_, _41265_, _41263_);
  not (_41266_, rxd_i);
  and (_41267_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _41266_);
  nor (_41268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_41269_, _41268_);
  and (_41270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_41271_, _41270_, _41269_);
  and (_41272_, _41271_, _41267_);
  not (_41273_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_41274_, _41273_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_41275_, _41274_, _41268_);
  or (_41276_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or (_41277_, _41276_, _41272_);
  and (_41278_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _42882_);
  and (_00551_, _41278_, _41277_);
  and (_41279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_41280_, _41279_, _41269_);
  nor (_41281_, _41268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41282_, _41281_, _41273_);
  nor (_41283_, _41282_, _41280_);
  not (_41284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_41285_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _41284_);
  not (_41286_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_41287_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _41286_);
  and (_41288_, _41287_, _41285_);
  not (_41289_, _41288_);
  or (_41290_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and (_41291_, _41288_, _41280_);
  and (_41292_, _41280_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41293_, _41292_, _41291_);
  and (_41294_, _41293_, _41290_);
  or (_41295_, _41294_, _41283_);
  not (_41296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand (_41297_, _41268_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_41298_, _41297_, _41296_);
  not (_41299_, _41298_);
  or (_41300_, _41299_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_41301_, _41300_, _41295_);
  nand (_00554_, _41301_, _41278_);
  not (_41302_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_41303_, _41280_);
  nor (_41304_, _41273_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_41305_, _41304_);
  not (_41306_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41307_, _41268_, _41306_);
  and (_41308_, _41307_, _41305_);
  and (_41309_, _41308_, _41303_);
  nor (_41310_, _41309_, _41302_);
  and (_41311_, _41309_, rxd_i);
  or (_41312_, _41311_, rst);
  or (_00556_, _41312_, _41310_);
  nor (_41313_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41314_, _41313_, _41285_);
  and (_41315_, _41314_, _41292_);
  nand (_41316_, _41315_, _41266_);
  or (_41317_, _41315_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_41318_, _41317_, _42882_);
  and (_00559_, _41318_, _41316_);
  and (_41319_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41320_, _41319_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41321_, _41320_, _41284_);
  and (_41322_, _41321_, _41292_);
  and (_41323_, _41271_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41324_, _41323_, _41292_);
  nor (_41325_, _41320_, _41303_);
  or (_41326_, _41325_, _41324_);
  and (_41327_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_41328_, _41327_, _41322_);
  and (_00562_, _41328_, _42882_);
  and (_41329_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _42882_);
  nand (_41330_, _41329_, _41306_);
  nand (_41331_, _41278_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand (_00564_, _41331_, _41330_);
  and (_41332_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41306_);
  not (_41333_, _41271_);
  nand (_41334_, _41275_, _41296_);
  and (_41335_, _41334_, _41333_);
  nand (_41336_, _41335_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand (_41337_, _41336_, _41303_);
  or (_41338_, _41288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_41339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_41340_, _41339_, _41291_);
  and (_41341_, _41340_, _41338_);
  and (_41342_, _41341_, _41337_);
  or (_41343_, _41342_, _41298_);
  nand (_41344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_41345_, _41344_, _41280_);
  or (_41346_, _41345_, _41289_);
  and (_41347_, _41346_, _41299_);
  or (_41348_, _41347_, rxd_i);
  and (_41349_, _41348_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41350_, _41349_, _41343_);
  or (_41351_, _41350_, _41332_);
  and (_00567_, _41351_, _42882_);
  and (_41352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_41353_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_41354_, _41254_, _41353_);
  or (_41355_, _41354_, _41257_);
  nor (_41356_, _41355_, _41352_);
  or (_41357_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_41358_, _41357_, _42882_);
  nor (_00570_, _41358_, _41356_);
  nor (_41359_, _41356_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_41360_, _41359_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_41361_, _41359_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_41362_, _41361_, _42882_);
  and (_00572_, _41362_, _41360_);
  not (_41363_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_41364_, _41297_, _41363_);
  nor (_41365_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not (_41366_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_41367_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_41368_, _41367_, _41366_);
  and (_41369_, _41368_, _41365_);
  not (_41370_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_41371_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_41372_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41373_, _41372_, _41371_);
  and (_41374_, _41373_, _41370_);
  and (_41375_, _41374_, _41369_);
  or (_41376_, _41375_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_41377_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41378_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_41379_, _41378_, _41377_);
  and (_41380_, _41269_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_41381_, _41380_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_41382_, _41381_, _41379_);
  not (_41383_, _41382_);
  or (_41384_, _41383_, _41376_);
  and (_41385_, _41379_, _41380_);
  or (_41386_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _41363_);
  or (_41387_, _41386_, _41385_);
  and (_41388_, _41387_, _41384_);
  or (_41389_, _41388_, _41364_);
  not (_41390_, _41364_);
  not (_41391_, _41375_);
  or (_41392_, _41391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_41393_, _41392_, _41376_);
  or (_41394_, _41393_, _41390_);
  nand (_41395_, _41394_, _41389_);
  and (_41396_, _40063_, _32556_);
  and (_41397_, _41396_, _30679_);
  and (_41398_, _41397_, _39227_);
  nor (_41399_, _41398_, rst);
  nand (_41400_, _41399_, _41395_);
  not (_41401_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_41402_, _41398_, _42882_);
  nand (_41403_, _41402_, _41401_);
  and (_00575_, _41403_, _41400_);
  nor (_41404_, _41391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand (_41405_, _41385_, _41404_);
  and (_41406_, _41375_, _41364_);
  or (_41407_, _41363_, rst);
  nor (_41408_, _41407_, _41406_);
  and (_41409_, _41408_, _41405_);
  or (_00578_, _41409_, _41402_);
  or (_41410_, _41383_, _41404_);
  or (_41411_, _41385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_41412_, _41297_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_41413_, _41412_, _41411_);
  and (_41414_, _41413_, _41410_);
  or (_41415_, _41414_, _41406_);
  and (_00580_, _41415_, _41399_);
  and (_41416_, _41381_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_41417_, _41416_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_41418_, _41417_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or (_41419_, _41418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_41420_, _41418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_41421_, _41420_, _41419_);
  and (_00583_, _41421_, _41399_);
  nor (_41422_, _41382_, _41364_);
  and (_41423_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_41424_, _41423_, _41399_);
  and (_41425_, _41402_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_00586_, _41425_, _41424_);
  and (_41426_, _40534_, _38405_);
  or (_41427_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_41428_, _41427_, _42882_);
  nand (_41429_, _41426_, _38485_);
  and (_00588_, _41429_, _41428_);
  and (_41430_, _40530_, _39205_);
  and (_41431_, _41430_, _31304_);
  nand (_41432_, _41431_, _31282_);
  and (_41433_, _40542_, _39227_);
  not (_41434_, _41433_);
  or (_41435_, _41431_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_41436_, _41435_, _41434_);
  and (_41437_, _41436_, _41432_);
  nor (_41438_, _41434_, _38485_);
  or (_41439_, _41438_, _41437_);
  and (_00591_, _41439_, _42882_);
  nor (_41440_, _41298_, _41291_);
  not (_41441_, _41440_);
  nor (_41442_, _41335_, _41280_);
  nor (_41443_, _41442_, _41441_);
  nor (_41444_, _41443_, _41306_);
  or (_41445_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_41446_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _41306_);
  or (_41447_, _41446_, _41440_);
  and (_41448_, _41447_, _42882_);
  and (_01210_, _41448_, _41445_);
  or (_41449_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_41450_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _41306_);
  or (_41451_, _41450_, _41440_);
  and (_41452_, _41451_, _42882_);
  and (_01212_, _41452_, _41449_);
  or (_41453_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_41454_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41306_);
  or (_41455_, _41454_, _41440_);
  and (_41456_, _41455_, _42882_);
  and (_01214_, _41456_, _41453_);
  or (_41457_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_41458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41306_);
  or (_41459_, _41458_, _41440_);
  and (_41460_, _41459_, _42882_);
  and (_01216_, _41460_, _41457_);
  or (_41461_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_41462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41306_);
  or (_41463_, _41462_, _41440_);
  and (_41464_, _41463_, _42882_);
  and (_01218_, _41464_, _41461_);
  or (_41465_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_41466_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41306_);
  or (_41467_, _41466_, _41440_);
  and (_41468_, _41467_, _42882_);
  and (_01220_, _41468_, _41465_);
  or (_41469_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_41470_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41306_);
  or (_41471_, _41470_, _41440_);
  and (_41472_, _41471_, _42882_);
  and (_01222_, _41472_, _41469_);
  or (_41473_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_41474_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _41306_);
  or (_41475_, _41474_, _41440_);
  and (_41476_, _41475_, _42882_);
  and (_01224_, _41476_, _41473_);
  nor (_41477_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_41478_, _41477_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_41479_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or (_41480_, _41288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_41481_, _41480_, _41280_);
  and (_41482_, _41481_, _41479_);
  or (_41483_, _41271_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_41484_, _41483_, _41334_);
  and (_41485_, _41484_, _41303_);
  or (_41486_, _41485_, _41482_);
  or (_41487_, _41486_, _41298_);
  or (_41488_, _41299_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_41489_, _41488_, _41278_);
  and (_41490_, _41489_, _41487_);
  or (_01226_, _41490_, _41478_);
  and (_41491_, _41288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_41492_, _41491_, _41335_);
  or (_41493_, _41492_, _41443_);
  and (_41494_, _41493_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_41495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _41306_);
  nand (_41496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41497_, _41496_, _41440_);
  or (_41498_, _41497_, _41495_);
  or (_41499_, _41498_, _41494_);
  and (_01228_, _41499_, _42882_);
  not (_41500_, _41444_);
  and (_41501_, _41500_, _41329_);
  or (_41502_, _41492_, _41441_);
  and (_41503_, _41278_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_41504_, _41503_, _41502_);
  or (_01229_, _41504_, _41501_);
  or (_41505_, _41322_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_41506_, _41322_, _41266_);
  and (_41507_, _41506_, _42882_);
  and (_01231_, _41507_, _41505_);
  or (_41508_, _41324_, _41286_);
  or (_41509_, _41292_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41510_, _41509_, _42882_);
  and (_01233_, _41510_, _41508_);
  and (_41511_, _41324_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_41512_, _41313_, _41319_);
  and (_41513_, _41512_, _41292_);
  or (_41514_, _41513_, _41511_);
  and (_01235_, _41514_, _42882_);
  and (_41515_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41516_, _41319_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41517_, _41516_, _41325_);
  or (_41518_, _41517_, _41515_);
  and (_01237_, _41518_, _42882_);
  and (_41519_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41306_);
  and (_41520_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41521_, _41520_, _41519_);
  and (_01239_, _41521_, _42882_);
  and (_41522_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41306_);
  and (_41523_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41524_, _41523_, _41522_);
  and (_01241_, _41524_, _42882_);
  and (_41525_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41306_);
  and (_41526_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41527_, _41526_, _41525_);
  and (_01243_, _41527_, _42882_);
  and (_41528_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41306_);
  and (_41529_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41530_, _41529_, _41528_);
  and (_01245_, _41530_, _42882_);
  and (_41531_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41306_);
  and (_41532_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41533_, _41532_, _41531_);
  and (_01247_, _41533_, _42882_);
  and (_41534_, _41278_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_01249_, _41534_, _41478_);
  and (_41535_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41536_, _41535_, _41495_);
  and (_01251_, _41536_, _42882_);
  nor (_41537_, _41381_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41538_, _41537_, _41416_);
  and (_01253_, _41538_, _41399_);
  nor (_41539_, _41416_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_41540_, _41539_, _41417_);
  and (_01255_, _41540_, _41399_);
  nor (_41541_, _41417_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_41542_, _41541_, _41418_);
  and (_01257_, _41542_, _41399_);
  or (_41543_, _41382_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41544_, _41383_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41545_, _41544_, _41543_);
  and (_41546_, _41545_, _41390_);
  and (_41547_, _41375_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41548_, _41547_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41549_, _41548_, _41364_);
  or (_41550_, _41549_, _41546_);
  and (_41551_, _41550_, _41399_);
  nor (_41552_, _41269_, _38464_);
  and (_41553_, _41552_, _41402_);
  or (_01259_, _41553_, _41551_);
  not (_41554_, _41422_);
  and (_41555_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_41556_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_41557_, _41556_, _41555_);
  and (_41558_, _41557_, _41399_);
  nand (_41559_, _41268_, _38456_);
  nand (_41560_, _41269_, _38464_);
  and (_41561_, _41560_, _41402_);
  and (_41562_, _41561_, _41559_);
  or (_01261_, _41562_, _41558_);
  nor (_41563_, _41422_, _41370_);
  and (_41564_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or (_41565_, _41564_, _41563_);
  and (_41566_, _41565_, _41399_);
  nand (_41567_, _41268_, _38449_);
  nand (_41568_, _41269_, _38456_);
  and (_41569_, _41568_, _41402_);
  and (_41570_, _41569_, _41567_);
  or (_01263_, _41570_, _41566_);
  nor (_41571_, _41422_, _41366_);
  and (_41572_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or (_41573_, _41572_, _41571_);
  and (_41574_, _41573_, _41399_);
  nand (_41575_, _41269_, _38449_);
  nand (_41576_, _41268_, _38442_);
  and (_41577_, _41576_, _41402_);
  and (_41578_, _41577_, _41575_);
  or (_01264_, _41578_, _41574_);
  and (_41579_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41580_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or (_41581_, _41580_, _41579_);
  and (_41582_, _41581_, _41399_);
  nand (_41583_, _41268_, _38434_);
  nand (_41584_, _41269_, _38442_);
  and (_41585_, _41584_, _41402_);
  and (_41586_, _41585_, _41583_);
  or (_01266_, _41586_, _41582_);
  and (_41587_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_41588_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or (_41589_, _41588_, _41587_);
  and (_41590_, _41589_, _41399_);
  nand (_41591_, _41269_, _38434_);
  nand (_41592_, _41268_, _38428_);
  and (_41593_, _41592_, _41402_);
  and (_41594_, _41593_, _41591_);
  or (_01268_, _41594_, _41590_);
  and (_41595_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_41596_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or (_41597_, _41596_, _41595_);
  and (_41598_, _41597_, _41399_);
  nand (_41599_, _41268_, _38420_);
  nand (_41600_, _41269_, _38428_);
  and (_41602_, _41600_, _41402_);
  and (_41604_, _41602_, _41599_);
  or (_01270_, _41604_, _41598_);
  and (_41607_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_41609_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_41611_, _41609_, _41607_);
  and (_41613_, _41611_, _41399_);
  nand (_41615_, _41268_, _38485_);
  nand (_41617_, _41269_, _38420_);
  and (_41619_, _41617_, _41402_);
  and (_41621_, _41619_, _41615_);
  or (_01272_, _41621_, _41613_);
  and (_41624_, _41398_, _41269_);
  nand (_41626_, _41624_, _38485_);
  and (_41628_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_41630_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_41632_, _41630_, _41628_);
  or (_41634_, _41632_, _41398_);
  and (_41636_, _41634_, _42882_);
  and (_01274_, _41636_, _41626_);
  and (_41639_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_41641_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_41643_, _41641_, _41639_);
  and (_41645_, _41643_, _41399_);
  or (_41647_, _41256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_41649_, _41647_, _41269_);
  and (_41651_, _41649_, _41402_);
  or (_01276_, _41651_, _41645_);
  nand (_41654_, _41426_, _38464_);
  or (_41656_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_41658_, _41656_, _42882_);
  and (_01278_, _41658_, _41654_);
  or (_41661_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_41663_, _41661_, _42882_);
  nand (_41665_, _41426_, _38456_);
  and (_01280_, _41665_, _41663_);
  or (_41666_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_41667_, _41666_, _42882_);
  nand (_41668_, _41426_, _38449_);
  and (_01282_, _41668_, _41667_);
  or (_41669_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_41670_, _41669_, _42882_);
  nand (_41671_, _41426_, _38442_);
  and (_01284_, _41671_, _41670_);
  or (_41672_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_41673_, _41672_, _42882_);
  nand (_41674_, _41426_, _38434_);
  and (_01286_, _41674_, _41673_);
  or (_41675_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_41676_, _41675_, _42882_);
  nand (_41677_, _41426_, _38428_);
  and (_01288_, _41677_, _41676_);
  or (_41678_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_41679_, _41678_, _42882_);
  nand (_41680_, _41426_, _38420_);
  and (_01290_, _41680_, _41679_);
  not (_41681_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_41682_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41681_);
  or (_41683_, _41682_, _41268_);
  nor (_41684_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41685_, _41684_, _41683_);
  or (_41686_, _41685_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_41687_, _41686_, _41430_);
  nand (_41688_, _39065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_41689_, _41688_, _41430_);
  or (_41690_, _41689_, _39070_);
  and (_41691_, _41690_, _41687_);
  or (_41692_, _41691_, _41433_);
  nand (_41693_, _41433_, _38464_);
  and (_41694_, _41693_, _42882_);
  and (_01292_, _41694_, _41692_);
  or (_41695_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_41696_, _41695_, _41430_);
  not (_41697_, _32567_);
  nor (_41698_, _41697_, _31282_);
  nand (_41699_, _41697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_41700_, _41699_, _41430_);
  or (_41701_, _41700_, _41698_);
  and (_41702_, _41701_, _41696_);
  or (_41703_, _41702_, _41433_);
  nand (_41704_, _41433_, _38456_);
  and (_41705_, _41704_, _42882_);
  and (_01294_, _41705_, _41703_);
  not (_41706_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not (_41707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_41708_, _41281_, _41707_);
  nor (_41709_, _41708_, _41706_);
  and (_41710_, _41708_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_41711_, _41710_, _41709_);
  or (_41712_, _41711_, _41430_);
  or (_41713_, _33296_, _41706_);
  nand (_41714_, _41713_, _41430_);
  or (_41715_, _41714_, _33318_);
  and (_41716_, _41715_, _41712_);
  or (_41717_, _41716_, _41433_);
  nand (_41718_, _41433_, _38449_);
  and (_41719_, _41718_, _42882_);
  and (_01296_, _41719_, _41717_);
  and (_41720_, _41430_, _34004_);
  nand (_41721_, _41720_, _31282_);
  or (_41722_, _41720_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_41723_, _41722_, _41434_);
  and (_41724_, _41723_, _41721_);
  nor (_41725_, _41434_, _38442_);
  or (_41726_, _41725_, _41724_);
  and (_01298_, _41726_, _42882_);
  and (_41727_, _41430_, _34765_);
  nand (_41728_, _41727_, _31282_);
  or (_41729_, _41727_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_41730_, _41729_, _41434_);
  and (_41731_, _41730_, _41728_);
  nor (_41732_, _41434_, _38434_);
  or (_41733_, _41732_, _41731_);
  and (_01299_, _41733_, _42882_);
  and (_41734_, _41430_, _35549_);
  nand (_41735_, _41734_, _31282_);
  or (_41736_, _41734_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_41737_, _41736_, _41434_);
  and (_41738_, _41737_, _41735_);
  nor (_41739_, _41434_, _38428_);
  or (_41740_, _41739_, _41738_);
  and (_01301_, _41740_, _42882_);
  and (_41741_, _41430_, _36277_);
  nand (_41742_, _41741_, _31282_);
  or (_41743_, _41741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_41744_, _41743_, _41434_);
  and (_41745_, _41744_, _41742_);
  nor (_41746_, _41434_, _38420_);
  or (_41747_, _41746_, _41745_);
  and (_01303_, _41747_, _42882_);
  and (_01628_, t2_i, _42882_);
  nor (_41748_, t2_i, rst);
  and (_01631_, _41748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand (_41749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _42882_);
  nor (_01634_, _41749_, t2ex_i);
  and (_01637_, t2ex_i, _42882_);
  and (_41750_, _38403_, _38895_);
  and (_41751_, _41750_, _39993_);
  nand (_41752_, _41751_, _38485_);
  and (_41753_, _41750_, _39840_);
  not (_41754_, _41753_);
  and (_41755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_41756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_41757_, _41756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41758_, _41757_, _41755_);
  not (_41759_, _41758_);
  and (_41760_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_41761_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_41762_, _41761_, _41760_);
  or (_41763_, _41751_, _41762_);
  and (_41764_, _41763_, _41754_);
  and (_41765_, _41764_, _41752_);
  and (_41766_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_41767_, _41766_, _41765_);
  and (_01640_, _41767_, _42882_);
  nand (_41768_, _41753_, _38485_);
  nor (_41769_, _41751_, _41759_);
  or (_41770_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_41771_, _41769_);
  or (_41772_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_41773_, _41772_, _41770_);
  or (_41774_, _41773_, _41753_);
  and (_41775_, _41774_, _42882_);
  and (_01643_, _41775_, _41768_);
  not (_41776_, _41756_);
  or (_41777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_41778_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_41779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _41778_);
  and (_41780_, _41779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_41781_, _41780_, _41777_);
  and (_41782_, _41781_, _41776_);
  and (_41783_, _41750_, _39954_);
  and (_41784_, _39839_, _35549_);
  and (_41785_, _41784_, _41750_);
  nor (_41786_, _41785_, _41783_);
  and (_41787_, _41786_, _41782_);
  and (_41788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_41789_, _41788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_41790_, _41789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_41791_, _41790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_41792_, _41791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_41793_, _41792_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_41794_, _41793_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_41795_, _41794_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_41796_, _41795_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_41797_, _41796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_41798_, _41797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_41799_, _41798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_41800_, _41799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_41801_, _41800_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_41802_, _41801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_41803_, _41802_);
  nand (_41804_, _41803_, _41787_);
  or (_41805_, _41787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_41806_, _41805_, _42882_);
  and (_01646_, _41806_, _41804_);
  nand (_41807_, _41783_, _38485_);
  and (_41808_, _41750_, _35549_);
  and (_41809_, _41808_, _39839_);
  not (_41810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41811_, _41755_, _41810_);
  and (_41812_, _41811_, _41756_);
  and (_41813_, _41812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not (_41814_, _41812_);
  not (_41815_, _41757_);
  and (_41816_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_41817_, _41802_, _41781_);
  and (_41818_, _41817_, _41816_);
  and (_41819_, _41793_, _41781_);
  or (_41820_, _41819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_41821_, _41819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_41822_, _41821_, _41820_);
  or (_41823_, _41822_, _41818_);
  and (_41824_, _41823_, _41814_);
  or (_41825_, _41824_, _41813_);
  nor (_41826_, _41825_, _41783_);
  nor (_41827_, _41826_, _41809_);
  and (_41828_, _41827_, _41807_);
  and (_41829_, _41809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_41830_, _41829_, _41828_);
  and (_01649_, _41830_, _42882_);
  and (_41831_, _41801_, _41781_);
  or (_41832_, _41831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_41833_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand (_41834_, _41833_, _41817_);
  and (_41835_, _41834_, _41832_);
  or (_41836_, _41835_, _41812_);
  or (_41837_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_41838_, _41837_, _41786_);
  and (_41839_, _41838_, _41836_);
  and (_41840_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_41841_, _41785_);
  nor (_41842_, _41841_, _38485_);
  or (_41843_, _41842_, _41840_);
  or (_41844_, _41843_, _41839_);
  and (_01652_, _41844_, _42882_);
  and (_41845_, _41814_, _41781_);
  and (_41846_, _41845_, _41756_);
  nand (_41847_, _41846_, _41802_);
  nand (_41848_, _41847_, _41786_);
  or (_41849_, _41786_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_41850_, _41849_, _42882_);
  and (_01655_, _41850_, _41848_);
  or (_41851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_41852_, _40546_, _38880_);
  or (_41853_, _41852_, _41851_);
  nand (_41854_, _38887_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_41855_, _41854_, _41852_);
  or (_41856_, _41855_, _38888_);
  and (_41857_, _41856_, _41853_);
  and (_41858_, _41750_, _40542_);
  or (_41859_, _41858_, _41857_);
  nand (_41860_, _41858_, _38485_);
  and (_41861_, _41860_, _42882_);
  and (_01658_, _41861_, _41859_);
  or (_41862_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not (_41863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_41864_, _41758_, _41863_);
  and (_41865_, _41864_, _41862_);
  or (_41866_, _41865_, _41751_);
  nand (_41867_, _41751_, _38464_);
  and (_41868_, _41867_, _41866_);
  or (_41869_, _41868_, _41753_);
  or (_41870_, _41754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_41871_, _41870_, _42882_);
  and (_02108_, _41871_, _41869_);
  nand (_41872_, _41751_, _38456_);
  and (_41873_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41874_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_41875_, _41874_, _41873_);
  or (_41876_, _41875_, _41751_);
  and (_41877_, _41876_, _41754_);
  and (_41878_, _41877_, _41872_);
  and (_41879_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_41880_, _41879_, _41878_);
  and (_02109_, _41880_, _42882_);
  nand (_41881_, _41751_, _38449_);
  and (_41882_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_41883_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_41884_, _41883_, _41882_);
  or (_41885_, _41884_, _41751_);
  and (_41886_, _41885_, _41754_);
  and (_41887_, _41886_, _41881_);
  and (_41888_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_41889_, _41888_, _41887_);
  and (_02111_, _41889_, _42882_);
  or (_41890_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_41891_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_41892_, _41891_, _41890_);
  or (_41893_, _41892_, _41751_);
  nand (_41894_, _41751_, _38442_);
  and (_41895_, _41894_, _41893_);
  or (_41896_, _41895_, _41753_);
  or (_41897_, _41754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_41898_, _41897_, _42882_);
  and (_02113_, _41898_, _41896_);
  nand (_41899_, _41751_, _38434_);
  and (_41900_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_41901_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_41902_, _41901_, _41900_);
  or (_41903_, _41902_, _41751_);
  and (_41904_, _41903_, _41754_);
  and (_41905_, _41904_, _41899_);
  and (_41906_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_41907_, _41906_, _41905_);
  and (_02115_, _41907_, _42882_);
  nand (_41908_, _41751_, _38428_);
  and (_41909_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_41910_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_41911_, _41910_, _41909_);
  or (_41912_, _41911_, _41751_);
  and (_41913_, _41912_, _41754_);
  and (_41914_, _41913_, _41908_);
  and (_41915_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_41916_, _41915_, _41914_);
  and (_02116_, _41916_, _42882_);
  nand (_41917_, _41751_, _38420_);
  and (_41918_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_41919_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_41920_, _41919_, _41918_);
  or (_41921_, _41920_, _41751_);
  and (_41922_, _41921_, _41754_);
  and (_41923_, _41922_, _41917_);
  and (_41924_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_41925_, _41924_, _41923_);
  and (_02118_, _41925_, _42882_);
  or (_41926_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_41927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_41928_, _41769_, _41927_);
  and (_41929_, _41928_, _41926_);
  or (_41930_, _41929_, _41753_);
  nand (_41931_, _41753_, _38464_);
  and (_41932_, _41931_, _42882_);
  and (_02120_, _41932_, _41930_);
  nand (_41933_, _41753_, _38456_);
  and (_41934_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_41935_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_41936_, _41935_, _41934_);
  or (_41937_, _41936_, _41753_);
  and (_41938_, _41937_, _42882_);
  and (_02122_, _41938_, _41933_);
  nand (_41939_, _41753_, _38449_);
  and (_41940_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_41941_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_41942_, _41941_, _41940_);
  or (_41943_, _41942_, _41753_);
  and (_41944_, _41943_, _42882_);
  and (_02123_, _41944_, _41939_);
  nand (_41945_, _41753_, _38442_);
  and (_41946_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_41947_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_41948_, _41947_, _41946_);
  or (_41949_, _41948_, _41753_);
  and (_41950_, _41949_, _42882_);
  and (_02125_, _41950_, _41945_);
  nand (_41951_, _41753_, _38434_);
  and (_41952_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_41953_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_41954_, _41953_, _41952_);
  or (_41955_, _41954_, _41753_);
  and (_41956_, _41955_, _42882_);
  and (_02127_, _41956_, _41951_);
  nand (_41957_, _41753_, _38428_);
  and (_41958_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_41959_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_41960_, _41959_, _41958_);
  or (_41961_, _41960_, _41753_);
  and (_41962_, _41961_, _42882_);
  and (_02129_, _41962_, _41957_);
  nand (_41963_, _41753_, _38420_);
  and (_41964_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_41965_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_41966_, _41965_, _41964_);
  or (_41967_, _41966_, _41753_);
  and (_41968_, _41967_, _42882_);
  and (_02130_, _41968_, _41963_);
  or (_41969_, _41781_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_41970_, _41781_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_41971_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_41972_, _41971_, _41802_);
  nand (_41973_, _41972_, _41970_);
  and (_41974_, _41973_, _41969_);
  or (_41975_, _41974_, _41812_);
  nor (_41976_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor (_41977_, _41976_, _41783_);
  and (_41978_, _41977_, _41975_);
  and (_41979_, _41783_, _38465_);
  or (_41980_, _41979_, _41809_);
  or (_41981_, _41980_, _41978_);
  nand (_41982_, _41785_, _41863_);
  and (_41983_, _41982_, _42882_);
  and (_02132_, _41983_, _41981_);
  and (_41984_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41985_, _41984_, _41845_);
  and (_41986_, _41985_, _41802_);
  and (_41987_, _41812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_41988_, _41970_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand (_41989_, _41788_, _41781_);
  and (_41990_, _41989_, _41814_);
  and (_41991_, _41990_, _41988_);
  nor (_41992_, _41991_, _41987_);
  nand (_41993_, _41992_, _41786_);
  or (_41994_, _41993_, _41986_);
  nand (_41995_, _41783_, _38456_);
  or (_41996_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_41997_, _41996_, _42882_);
  and (_41998_, _41997_, _41995_);
  and (_02134_, _41998_, _41994_);
  not (_41999_, _41783_);
  or (_42000_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_42001_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_42002_, _42001_, _41817_);
  and (_42003_, _41989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_42004_, _41989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_42005_, _42004_, _41812_);
  or (_42006_, _42005_, _42003_);
  or (_42007_, _42006_, _42002_);
  nand (_42008_, _42007_, _42000_);
  nand (_42009_, _42008_, _41999_);
  nand (_42010_, _41783_, _38449_);
  and (_42011_, _42010_, _42009_);
  or (_42012_, _42011_, _41785_);
  or (_42013_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_42014_, _42013_, _42882_);
  and (_02136_, _42014_, _42012_);
  or (_42015_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_42016_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_42017_, _42016_, _41817_);
  nand (_42018_, _41789_, _41781_);
  and (_42019_, _42018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_42020_, _42018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_42021_, _42020_, _41812_);
  or (_42022_, _42021_, _42019_);
  or (_42023_, _42022_, _42017_);
  nand (_42024_, _42023_, _42015_);
  nand (_42025_, _42024_, _41999_);
  nand (_42026_, _41783_, _38442_);
  and (_42027_, _42026_, _42025_);
  or (_42028_, _42027_, _41785_);
  or (_42029_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_42030_, _42029_, _42882_);
  and (_02137_, _42030_, _42028_);
  and (_42031_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_42032_, _42031_, _41817_);
  nand (_42033_, _41790_, _41781_);
  and (_42034_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_42035_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_42036_, _42035_, _41812_);
  or (_42037_, _42036_, _42034_);
  or (_42038_, _42037_, _42032_);
  nor (_42039_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor (_42040_, _42039_, _41783_);
  and (_42041_, _42040_, _42038_);
  nor (_42042_, _41999_, _38434_);
  or (_42043_, _42042_, _42041_);
  or (_42044_, _42043_, _41809_);
  or (_42045_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_42046_, _42045_, _42882_);
  and (_02139_, _42046_, _42044_);
  and (_42047_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_42048_, _42047_, _41817_);
  nand (_42049_, _41791_, _41781_);
  and (_42050_, _42049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_42051_, _42049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_42052_, _42051_, _41812_);
  or (_42053_, _42052_, _42050_);
  or (_42054_, _42053_, _42048_);
  nor (_42055_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor (_42056_, _42055_, _41783_);
  and (_42057_, _42056_, _42054_);
  nor (_42058_, _41999_, _38428_);
  or (_42059_, _42058_, _42057_);
  or (_42060_, _42059_, _41809_);
  or (_42061_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_42062_, _42061_, _42882_);
  and (_02141_, _42062_, _42060_);
  nor (_42063_, _41999_, _38420_);
  and (_42064_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_42065_, _42064_, _41817_);
  and (_42066_, _41792_, _41781_);
  nor (_42067_, _42066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_42068_, _42067_, _41819_);
  or (_42069_, _42068_, _41812_);
  or (_42070_, _42069_, _42065_);
  nor (_42071_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_42072_, _42071_, _41783_);
  and (_42073_, _42072_, _42070_);
  or (_42074_, _42073_, _41809_);
  or (_42075_, _42074_, _42063_);
  or (_42076_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_42077_, _42076_, _42882_);
  and (_02143_, _42077_, _42075_);
  and (_42078_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_42079_, _42078_, _41817_);
  nand (_42080_, _41821_, _41927_);
  or (_42081_, _41821_, _41927_);
  and (_42082_, _42081_, _42080_);
  or (_42083_, _42082_, _41812_);
  or (_42084_, _42083_, _42079_);
  nor (_42085_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_42086_, _42085_, _41783_);
  and (_42087_, _42086_, _42084_);
  and (_42088_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_42089_, _42088_, _41809_);
  or (_42090_, _42089_, _42087_);
  nand (_42091_, _41785_, _38464_);
  and (_42092_, _42091_, _42882_);
  and (_02144_, _42092_, _42090_);
  and (_42093_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_42094_, _42093_, _41817_);
  and (_42095_, _41795_, _41781_);
  or (_42096_, _42095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_42097_, _42095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_42098_, _42097_, _42096_);
  or (_42099_, _42098_, _41812_);
  or (_42100_, _42099_, _42094_);
  nor (_42101_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_42102_, _42101_, _41783_);
  and (_42103_, _42102_, _42100_);
  and (_42104_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_42105_, _42104_, _41809_);
  or (_42106_, _42105_, _42103_);
  nand (_42107_, _41809_, _38456_);
  and (_42108_, _42107_, _42882_);
  and (_02145_, _42108_, _42106_);
  and (_42109_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_42110_, _42109_, _41817_);
  nand (_42111_, _41796_, _41781_);
  and (_42112_, _42111_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_42113_, _42111_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_42114_, _42113_, _41812_);
  or (_42115_, _42114_, _42112_);
  or (_42116_, _42115_, _42110_);
  nor (_42117_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_42118_, _42117_, _41783_);
  and (_42119_, _42118_, _42116_);
  and (_42120_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_42121_, _42120_, _41809_);
  or (_42122_, _42121_, _42119_);
  nand (_42123_, _41809_, _38449_);
  and (_42124_, _42123_, _42882_);
  and (_02146_, _42124_, _42122_);
  and (_42125_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_42126_, _42125_, _41817_);
  nand (_42127_, _41797_, _41781_);
  and (_42128_, _42127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor (_42129_, _42127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_42130_, _42129_, _41812_);
  or (_42131_, _42130_, _42128_);
  or (_42132_, _42131_, _42126_);
  nor (_42133_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_42134_, _42133_, _41783_);
  and (_42135_, _42134_, _42132_);
  and (_42136_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_42137_, _42136_, _41809_);
  or (_42138_, _42137_, _42135_);
  nand (_42139_, _41809_, _38442_);
  and (_42140_, _42139_, _42882_);
  and (_02147_, _42140_, _42138_);
  nand (_42141_, _41785_, _38434_);
  and (_42142_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_42143_, _42142_, _41817_);
  nand (_42144_, _41798_, _41781_);
  and (_42145_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_42146_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_42147_, _42146_, _41812_);
  or (_42148_, _42147_, _42145_);
  or (_42149_, _42148_, _42143_);
  nor (_42150_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_42151_, _42150_, _41783_);
  and (_42152_, _42151_, _42149_);
  and (_42153_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_42154_, _42153_, _41809_);
  or (_42155_, _42154_, _42152_);
  and (_42156_, _42155_, _42882_);
  and (_02148_, _42156_, _42141_);
  and (_42157_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_42158_, _42157_, _41817_);
  nand (_42159_, _41799_, _41781_);
  and (_42160_, _42159_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_42161_, _42159_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_42162_, _42161_, _41812_);
  or (_42163_, _42162_, _42160_);
  or (_42164_, _42163_, _42158_);
  nor (_42165_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor (_42166_, _42165_, _41783_);
  and (_42167_, _42166_, _42164_);
  and (_42168_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_42169_, _42168_, _41809_);
  or (_42170_, _42169_, _42167_);
  nand (_42171_, _41809_, _38428_);
  and (_42172_, _42171_, _42882_);
  and (_02149_, _42172_, _42170_);
  and (_42173_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_42174_, _42173_, _41817_);
  and (_42175_, _41800_, _41781_);
  nor (_42176_, _42175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_42177_, _42176_, _41831_);
  or (_42178_, _42177_, _41812_);
  or (_42179_, _42178_, _42174_);
  nor (_42180_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_42181_, _42180_, _41783_);
  and (_42182_, _42181_, _42179_);
  and (_42183_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_42184_, _42183_, _41809_);
  or (_42185_, _42184_, _42182_);
  nand (_42186_, _41809_, _38420_);
  and (_42187_, _42186_, _42882_);
  and (_02150_, _42187_, _42185_);
  and (_42188_, _41852_, _27045_);
  nand (_42189_, _42188_, _31282_);
  or (_42190_, _42188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_42191_, _42190_, _42189_);
  or (_42192_, _42191_, _41858_);
  nand (_42193_, _41858_, _38464_);
  and (_42194_, _42193_, _42882_);
  and (_02151_, _42194_, _42192_);
  not (_42195_, _41858_);
  and (_42196_, _41852_, _32567_);
  or (_42197_, _42196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_42198_, _42197_, _42195_);
  nand (_42199_, _42196_, _31282_);
  and (_42200_, _42199_, _42198_);
  nor (_42201_, _42195_, _38456_);
  or (_42202_, _42201_, _42200_);
  and (_02152_, _42202_, _42882_);
  nand (_42203_, _41852_, _39293_);
  and (_42204_, _42203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_42205_, _42204_, _41858_);
  and (_42206_, _33329_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_42207_, _42206_, _33318_);
  and (_42208_, _42207_, _41852_);
  or (_42209_, _42208_, _42205_);
  nand (_42210_, _41858_, _38449_);
  and (_42211_, _42210_, _42882_);
  and (_02153_, _42211_, _42209_);
  and (_42212_, _41852_, _34004_);
  or (_42213_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_42214_, _42213_, _42195_);
  nand (_42215_, _42212_, _31282_);
  and (_42216_, _42215_, _42214_);
  nor (_42217_, _42195_, _38442_);
  or (_42218_, _42217_, _42216_);
  and (_02154_, _42218_, _42882_);
  and (_42219_, _41852_, _34765_);
  or (_42220_, _42219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_42221_, _42220_, _42195_);
  nand (_42222_, _42219_, _31282_);
  and (_42223_, _42222_, _42221_);
  nor (_42224_, _42195_, _38434_);
  or (_42225_, _42224_, _42223_);
  and (_02155_, _42225_, _42882_);
  and (_42226_, _41852_, _35549_);
  nand (_42227_, _42226_, _31282_);
  or (_42228_, _42226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_42229_, _42228_, _42227_);
  or (_42230_, _42229_, _41858_);
  nand (_42231_, _41858_, _38428_);
  and (_42232_, _42231_, _42882_);
  and (_02156_, _42232_, _42230_);
  not (_42233_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_42234_, _41755_, _42233_);
  or (_42235_, _42234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_42236_, _42235_, _41852_);
  nand (_42237_, _39006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_42238_, _42237_, _41852_);
  or (_42239_, _42238_, _39007_);
  and (_42240_, _42239_, _42236_);
  or (_42241_, _42240_, _41858_);
  nand (_42242_, _41858_, _38420_);
  and (_42243_, _42242_, _42882_);
  and (_02157_, _42243_, _42241_);
  and (_42244_, _30646_, _27527_);
  not (_42245_, _38487_);
  and (_42246_, _42245_, _38399_);
  not (_42247_, _42246_);
  not (_42248_, _38398_);
  nor (_42249_, _42248_, _38357_);
  not (_42250_, _36450_);
  and (_42251_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_42252_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_42253_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_42254_, _42253_, _42252_);
  and (_42255_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_42256_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_42257_, _42256_, _42255_);
  and (_42258_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_42259_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_42260_, _42259_, _42258_);
  and (_42261_, _42260_, _42257_);
  and (_42262_, _42261_, _42254_);
  nor (_42263_, _36636_, _42250_);
  not (_42264_, _42263_);
  nor (_42265_, _42264_, _42262_);
  nor (_42266_, _42265_, _42251_);
  not (_42267_, _42266_);
  and (_42268_, _42267_, _42249_);
  not (_42269_, _42268_);
  not (_42270_, _38257_);
  and (_42271_, _42248_, _38357_);
  nor (_42272_, _38901_, _38948_);
  nor (_42273_, _42272_, _38954_);
  and (_42274_, _42273_, _27714_);
  nor (_42275_, _30657_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_42276_, _42275_, _33329_);
  not (_42277_, _42276_);
  nor (_42278_, _42277_, _42274_);
  nor (_42279_, _42273_, _27714_);
  and (_42280_, _37960_, _27023_);
  nor (_42281_, _37960_, _27023_);
  nor (_42282_, _42281_, _42280_);
  not (_42283_, _42282_);
  nor (_42284_, _42283_, _42279_);
  and (_42285_, _42284_, _42278_);
  not (_42286_, _42285_);
  and (_42287_, _42273_, _38262_);
  and (_42288_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_42289_, _42273_, _37960_);
  and (_42290_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_42291_, _42290_, _42288_);
  nor (_42292_, _42273_, _38262_);
  and (_42293_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_42294_, _42273_, _37960_);
  and (_42295_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_42296_, _42295_, _42293_);
  and (_42297_, _42296_, _42291_);
  and (_42298_, _42297_, _42286_);
  and (_42299_, _42285_, _38485_);
  nor (_42300_, _42299_, _42298_);
  and (_42301_, _42300_, _42271_);
  nor (_42302_, _42301_, _42270_);
  and (_42303_, _42302_, _42269_);
  and (_42304_, _42303_, _42247_);
  and (_42305_, _38246_, _38317_);
  nor (_42306_, _42305_, _38325_);
  not (_42307_, _42306_);
  nor (_42308_, _42307_, _38273_);
  and (_42309_, _42308_, _38319_);
  and (_42310_, _38246_, _37707_);
  nor (_42311_, _42310_, _38320_);
  and (_42312_, _42311_, _38341_);
  and (_42313_, _42312_, _42309_);
  and (_42314_, _42313_, _38268_);
  nor (_42315_, _42314_, _36407_);
  nor (_42316_, _38339_, _38335_);
  not (_42317_, _38243_);
  nor (_42318_, _42317_, _42316_);
  nor (_42319_, _42318_, _42315_);
  not (_42320_, _42319_);
  and (_42321_, _42320_, _42304_);
  and (_42322_, _42249_, _38257_);
  and (_42323_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_42324_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_42325_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_42326_, _42325_, _42324_);
  and (_42327_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_42328_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_42329_, _42328_, _42327_);
  and (_42330_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_42331_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_42332_, _42331_, _42330_);
  and (_42333_, _42332_, _42329_);
  and (_42334_, _42333_, _42326_);
  nor (_42335_, _42334_, _42264_);
  nor (_42336_, _42335_, _42323_);
  not (_42337_, _42336_);
  and (_42338_, _42337_, _42322_);
  and (_42339_, _38398_, _38357_);
  and (_42340_, _42339_, _38257_);
  and (_42341_, _38904_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_42342_, _42341_, _38966_);
  not (_42343_, _42342_);
  and (_42344_, _42343_, _42340_);
  nor (_42345_, _42344_, _42338_);
  and (_42346_, _42271_, _38257_);
  nor (_42347_, _42286_, _38434_);
  and (_42348_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_42349_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_42350_, _42349_, _42348_);
  and (_42351_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_42352_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_42353_, _42352_, _42351_);
  and (_42354_, _42353_, _42350_);
  nor (_42355_, _42354_, _42285_);
  nor (_42356_, _42355_, _42347_);
  not (_42357_, _42356_);
  and (_42358_, _42357_, _42346_);
  not (_42359_, _42358_);
  not (_42360_, _38519_);
  and (_42361_, _42360_, _38400_);
  and (_42362_, _42270_, _38398_);
  nor (_42363_, _42362_, _42361_);
  and (_42364_, _42363_, _42359_);
  and (_42365_, _42364_, _42345_);
  not (_42366_, _42365_);
  and (_42367_, _42366_, _42321_);
  and (_42368_, _42271_, _42270_);
  and (_42369_, _42340_, _38190_);
  or (_42370_, _42369_, _42368_);
  and (_42371_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_42372_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_42373_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_42374_, _42373_, _42372_);
  and (_42375_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_42376_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_42377_, _42376_, _42375_);
  and (_42378_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_42379_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_42380_, _42379_, _42378_);
  and (_42381_, _42380_, _42377_);
  and (_42382_, _42381_, _42374_);
  nor (_42383_, _42382_, _42264_);
  nor (_42384_, _42383_, _42371_);
  not (_42385_, _42384_);
  and (_42386_, _42385_, _42322_);
  not (_42387_, _38501_);
  and (_42388_, _42387_, _38400_);
  and (_42389_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_42390_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_42391_, _42390_, _42389_);
  and (_42392_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_42393_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_42394_, _42393_, _42392_);
  and (_42395_, _42394_, _42391_);
  and (_42396_, _42395_, _42286_);
  and (_42397_, _42285_, _38456_);
  nor (_42398_, _42397_, _42396_);
  and (_42399_, _42398_, _42346_);
  or (_42400_, _42399_, _42388_);
  or (_42401_, _42400_, _42386_);
  nor (_42402_, _42401_, _42370_);
  nor (_42403_, _42402_, _42320_);
  nor (_42404_, _42403_, _42367_);
  not (_42405_, _27845_);
  and (_42406_, _27549_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42407_, _42406_, _42405_);
  nor (_42408_, _26902_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42409_, _42408_, _42407_);
  nand (_42410_, _42409_, _42404_);
  or (_42411_, _42409_, _42404_);
  and (_42412_, _42411_, _42410_);
  not (_42413_, _42412_);
  not (_42414_, _42273_);
  and (_42415_, _42340_, _42414_);
  and (_42416_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_42417_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_42418_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_42419_, _42418_, _42417_);
  and (_42420_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_42421_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_42422_, _42421_, _42420_);
  and (_42423_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_42424_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_42425_, _42424_, _42423_);
  and (_42426_, _42425_, _42422_);
  and (_42427_, _42426_, _42419_);
  nor (_42428_, _42427_, _42264_);
  nor (_42429_, _42428_, _42416_);
  not (_42430_, _42429_);
  and (_42431_, _42430_, _42322_);
  nor (_42432_, _42431_, _42415_);
  not (_42433_, _38513_);
  and (_42434_, _42433_, _38400_);
  and (_42435_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_42436_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_42437_, _42436_, _42435_);
  and (_42438_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_42439_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_42440_, _42439_, _42438_);
  and (_42441_, _42440_, _42437_);
  nor (_42442_, _42441_, _42285_);
  nor (_42443_, _42286_, _38442_);
  nor (_42444_, _42443_, _42442_);
  not (_42445_, _42444_);
  and (_42446_, _42445_, _42346_);
  nor (_42447_, _42446_, _42434_);
  and (_42448_, _42447_, _42432_);
  not (_42449_, _42448_);
  and (_42450_, _42449_, _42321_);
  and (_42451_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_42452_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_42453_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_42454_, _42453_, _42452_);
  and (_42455_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_42456_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_42457_, _42456_, _42455_);
  and (_42458_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_42459_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_42460_, _42459_, _42458_);
  and (_42461_, _42460_, _42457_);
  and (_42462_, _42461_, _42454_);
  nor (_42463_, _42462_, _42264_);
  nor (_42464_, _42463_, _42451_);
  not (_42465_, _42464_);
  and (_42466_, _42465_, _42322_);
  and (_42467_, _42285_, _38465_);
  and (_42468_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_42469_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_42470_, _42469_, _42468_);
  and (_42471_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_42472_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_42473_, _42472_, _42471_);
  and (_42474_, _42473_, _42470_);
  nor (_42475_, _42474_, _42285_);
  nor (_42476_, _42475_, _42467_);
  not (_42477_, _42476_);
  and (_42478_, _42477_, _42346_);
  nor (_42479_, _42478_, _42466_);
  not (_42480_, _38495_);
  and (_42481_, _42480_, _38400_);
  and (_42482_, _42340_, _37960_);
  nor (_42483_, _42482_, _42481_);
  and (_42484_, _42483_, _42479_);
  nor (_42485_, _42484_, _42320_);
  nor (_42486_, _42485_, _42450_);
  and (_42487_, _42406_, _27714_);
  nor (_42488_, _27023_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42489_, _42488_, _42487_);
  not (_42490_, _42489_);
  and (_42491_, _42490_, _42486_);
  nor (_42492_, _42490_, _42486_);
  nor (_42493_, _42492_, _42491_);
  and (_42494_, _42493_, _42413_);
  nor (_42495_, _42271_, _38257_);
  and (_42496_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_42497_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_42498_, _42497_, _42496_);
  and (_42499_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_42500_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_42501_, _42500_, _42499_);
  and (_42502_, _42501_, _42498_);
  and (_42503_, _42502_, _42286_);
  and (_42504_, _42285_, _38420_);
  nor (_42505_, _42504_, _42503_);
  and (_42506_, _42505_, _42346_);
  nor (_42507_, _42506_, _42495_);
  not (_42508_, _38531_);
  and (_42509_, _42508_, _38400_);
  and (_42510_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_42511_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_42512_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_42513_, _42512_, _42511_);
  and (_42514_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_42515_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_42516_, _42515_, _42514_);
  and (_42517_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_42518_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_42519_, _42518_, _42517_);
  and (_42520_, _42519_, _42516_);
  and (_42521_, _42520_, _42513_);
  nor (_42522_, _42521_, _42264_);
  nor (_42523_, _42522_, _42510_);
  not (_42524_, _42523_);
  and (_42525_, _42524_, _42322_);
  nor (_42526_, _42525_, _42509_);
  and (_42527_, _42526_, _42507_);
  and (_42528_, _42527_, _42321_);
  nor (_42529_, _42449_, _42321_);
  nor (_42530_, _42529_, _42528_);
  nor (_42531_, _42406_, _27714_);
  and (_42532_, _42406_, _27242_);
  nor (_42533_, _42532_, _42531_);
  not (_42534_, _42533_);
  and (_42535_, _42534_, _42530_);
  nor (_42536_, _42534_, _42530_);
  nor (_42537_, _42536_, _42535_);
  and (_42538_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_42539_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_42540_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_42541_, _42540_, _42539_);
  and (_42542_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_42543_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_42544_, _42543_, _42542_);
  and (_42545_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_42546_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_42547_, _42546_, _42545_);
  and (_42548_, _42547_, _42544_);
  and (_42549_, _42548_, _42541_);
  nor (_42550_, _42549_, _42264_);
  nor (_42551_, _42550_, _42538_);
  not (_42552_, _42551_);
  and (_42553_, _42552_, _42322_);
  and (_42554_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  not (_42555_, _42554_);
  and (_42556_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_42557_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_42558_, _42557_, _42556_);
  and (_42559_, _42558_, _42555_);
  and (_42560_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_42561_, _42560_, _42285_);
  and (_42562_, _42561_, _42559_);
  and (_42563_, _42285_, _38428_);
  or (_42564_, _42563_, _42562_);
  not (_42565_, _42564_);
  and (_42566_, _42565_, _42346_);
  nor (_42567_, _42566_, _42553_);
  nor (_42568_, _38525_, _38398_);
  nor (_42569_, _42568_, _42270_);
  or (_42570_, _42249_, _42271_);
  nor (_42571_, _42570_, _42569_);
  not (_42572_, _42571_);
  and (_42573_, _42572_, _42567_);
  not (_42574_, _42573_);
  and (_42575_, _42574_, _42321_);
  and (_42576_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_42577_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_42578_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_42579_, _42578_, _42577_);
  and (_42580_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_42581_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_42582_, _42581_, _42580_);
  and (_42583_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_42584_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_42585_, _42584_, _42583_);
  and (_42586_, _42585_, _42582_);
  and (_42587_, _42586_, _42579_);
  nor (_42588_, _42587_, _42264_);
  nor (_42589_, _42588_, _42576_);
  not (_42590_, _42589_);
  and (_42591_, _42590_, _42322_);
  and (_42592_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_42593_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_42594_, _42593_, _42592_);
  and (_42595_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_42596_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_42597_, _42596_, _42595_);
  and (_42598_, _42597_, _42594_);
  nor (_42599_, _42598_, _42285_);
  not (_42600_, _38449_);
  and (_42601_, _42285_, _42600_);
  nor (_42602_, _42601_, _42599_);
  not (_42603_, _42602_);
  and (_42604_, _42603_, _42346_);
  nor (_42605_, _42604_, _42591_);
  not (_42606_, _38507_);
  and (_42607_, _42606_, _38400_);
  and (_42608_, _42340_, _38167_);
  nor (_42609_, _42608_, _42607_);
  and (_42610_, _42609_, _42605_);
  nor (_42611_, _42610_, _42320_);
  nor (_42612_, _42611_, _42575_);
  and (_42613_, _42406_, _38879_);
  nor (_42614_, _26781_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42615_, _42614_, _42613_);
  not (_42616_, _42615_);
  nor (_42617_, _42616_, _42612_);
  and (_42618_, _42616_, _42612_);
  nor (_42619_, _42618_, _42617_);
  and (_42620_, _42619_, _42537_);
  and (_42621_, _42620_, _42494_);
  and (_42622_, _42621_, _42244_);
  nor (_42623_, _42365_, _42321_);
  nor (_42624_, _42406_, _27845_);
  not (_42625_, _42624_);
  and (_42626_, _42625_, _42623_);
  nor (_42627_, _42625_, _42623_);
  nor (_42628_, _42627_, _42626_);
  nor (_42629_, _42574_, _42321_);
  nor (_42630_, _42406_, _38879_);
  not (_42631_, _42630_);
  and (_42632_, _42631_, _42629_);
  nor (_42633_, _42631_, _42629_);
  nor (_42634_, _42633_, _42632_);
  and (_42635_, _42634_, _42628_);
  nor (_42636_, _42304_, _27549_);
  and (_42637_, _42304_, _27549_);
  nor (_42638_, _42637_, _42636_);
  not (_42639_, _42638_);
  nor (_42640_, _42527_, _42321_);
  nor (_42641_, _42406_, _27242_);
  not (_42642_, _42641_);
  nor (_42643_, _42642_, _42640_);
  and (_42644_, _42642_, _42640_);
  nor (_42645_, _42644_, _42643_);
  and (_42646_, _42645_, _42639_);
  and (_42647_, _42646_, _42635_);
  and (_42648_, _42647_, _42622_);
  not (_42649_, _42612_);
  not (_42650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_42651_, _42486_, _42650_);
  and (_42652_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_42653_, _42652_, _42404_);
  or (_42654_, _42653_, _42651_);
  and (_42655_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_42656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_42657_, _42486_, _42656_);
  nand (_42658_, _42657_, _42404_);
  or (_42659_, _42658_, _42655_);
  and (_42660_, _42659_, _42654_);
  or (_42661_, _42660_, _42649_);
  not (_42662_, _42530_);
  not (_42663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_42664_, _42486_, _42663_);
  and (_42665_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_42666_, _42665_, _42404_);
  or (_42667_, _42666_, _42664_);
  and (_42668_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not (_42669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_42670_, _42486_, _42669_);
  nand (_42671_, _42670_, _42404_);
  or (_42672_, _42671_, _42668_);
  and (_42673_, _42672_, _42667_);
  or (_42674_, _42673_, _42612_);
  and (_42675_, _42674_, _42662_);
  and (_42676_, _42675_, _42661_);
  not (_42677_, _42404_);
  not (_42678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_42679_, _42486_, _42678_);
  or (_42680_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_42681_, _42680_, _42679_);
  or (_42682_, _42681_, _42677_);
  or (_42683_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_42684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_42685_, _42486_, _42684_);
  and (_42686_, _42685_, _42683_);
  or (_42687_, _42686_, _42404_);
  and (_42688_, _42687_, _42682_);
  or (_42689_, _42688_, _42649_);
  not (_42690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_42691_, _42486_, _42690_);
  or (_42692_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_42693_, _42692_, _42691_);
  or (_42694_, _42693_, _42677_);
  or (_42695_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_42696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_42697_, _42486_, _42696_);
  and (_42698_, _42697_, _42695_);
  or (_42699_, _42698_, _42404_);
  and (_42700_, _42699_, _42694_);
  or (_42701_, _42700_, _42612_);
  and (_42702_, _42701_, _42530_);
  and (_42703_, _42702_, _42689_);
  nor (_42704_, _42703_, _42676_);
  nor (_42705_, _42704_, _42648_);
  not (_42706_, _42622_);
  nor (_42707_, _42648_, _42706_);
  and (_42708_, _42648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  or (_42709_, _42708_, _42707_);
  or (_42710_, _42709_, _42705_);
  nor (_42711_, _42707_, rst);
  and (_42712_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_42713_, _42712_, _28723_);
  nor (_42714_, _42713_, _31282_);
  nand (_42715_, _28723_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42716_, _20040_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42717_, _42716_, _42715_);
  nor (_42718_, _38485_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_42719_, _42718_, _42717_);
  or (_42720_, _42719_, _42714_);
  and (_40016_, _42720_, _42882_);
  or (_42721_, _40016_, _42711_);
  and (_02563_, _42721_, _42710_);
  not (_42722_, _42244_);
  nor (_42723_, _42489_, _42722_);
  nor (_42724_, _42722_, _42409_);
  and (_42725_, _42724_, _42723_);
  and (_42726_, _42533_, _42244_);
  nor (_42727_, _42722_, _42615_);
  and (_42728_, _42727_, _42726_);
  and (_42729_, _42728_, _42725_);
  and (_42730_, _42720_, _42244_);
  and (_42731_, _42730_, _42729_);
  not (_42732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_42733_, _42729_, _42732_);
  or (_02573_, _42733_, _42731_);
  nor (_42734_, _42727_, _42726_);
  nor (_42735_, _42724_, _42723_);
  and (_42736_, _42735_, _42244_);
  and (_42737_, _42736_, _42734_);
  and (_42738_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _28635_);
  and (_42739_, _42738_, _28690_);
  not (_42740_, _42739_);
  nor (_42741_, _42740_, _31282_);
  not (_42742_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42743_, _38464_, _42742_);
  or (_42744_, _18878_, _42742_);
  and (_42745_, _42744_, _42740_);
  and (_42746_, _42745_, _42743_);
  or (_42747_, _42746_, _42741_);
  and (_42748_, _42747_, _42737_);
  not (_42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_42750_, _42737_, _42749_);
  or (_02796_, _42750_, _42748_);
  nand (_42751_, _42738_, _28657_);
  nor (_42752_, _42751_, _31282_);
  nor (_42753_, _38456_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42754_, _42738_, _28744_);
  and (_42755_, _42738_, _28723_);
  or (_42756_, _42755_, _42712_);
  or (_42757_, _42756_, _42754_);
  and (_42758_, _42757_, _19871_);
  or (_42759_, _42758_, _42753_);
  or (_42760_, _42759_, _42752_);
  and (_42761_, _42760_, _42737_);
  not (_42762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_42763_, _42737_, _42762_);
  or (_02801_, _42763_, _42761_);
  not (_42764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_42765_, _42737_, _42764_);
  nand (_42766_, _42738_, _28755_);
  nor (_42767_, _42766_, _31282_);
  nor (_42768_, _38449_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42769_, _42738_, _28646_);
  or (_42770_, _42769_, _42756_);
  and (_42771_, _42770_, _18516_);
  or (_42772_, _42771_, _42768_);
  or (_42773_, _42772_, _42767_);
  and (_42774_, _42773_, _42737_);
  or (_02806_, _42774_, _42765_);
  and (_42775_, _42755_, _31859_);
  nor (_42776_, _38442_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_42777_, _42754_, _42712_);
  or (_42778_, _42777_, _42769_);
  and (_42779_, _42778_, _19544_);
  or (_42780_, _42779_, _42776_);
  or (_42781_, _42780_, _42775_);
  and (_42782_, _42781_, _42737_);
  not (_42783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_42784_, _42737_, _42783_);
  or (_02811_, _42784_, _42782_);
  not (_42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_42786_, _42737_, _42785_);
  nand (_42787_, _42712_, _28690_);
  nor (_42788_, _42787_, _31282_);
  nor (_42789_, _38434_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42790_, _28690_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42791_, _18714_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42792_, _42791_, _42790_);
  or (_42793_, _42792_, _42789_);
  or (_42794_, _42793_, _42788_);
  and (_42795_, _42794_, _42737_);
  or (_02815_, _42795_, _42786_);
  nand (_42796_, _42712_, _28657_);
  nor (_42797_, _42796_, _31282_);
  nor (_42798_, _38428_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42799_, _28657_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42800_, _19696_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42801_, _42800_, _42799_);
  or (_42802_, _42801_, _42798_);
  or (_42803_, _42802_, _42797_);
  and (_42804_, _42803_, _42737_);
  not (_42805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_42806_, _42737_, _42805_);
  or (_02820_, _42806_, _42804_);
  nand (_42807_, _42712_, _28755_);
  nor (_42808_, _42807_, _31282_);
  nor (_42809_, _38420_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42810_, _28755_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42811_, _19054_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42812_, _42811_, _42810_);
  or (_42813_, _42812_, _42809_);
  or (_42814_, _42813_, _42808_);
  and (_42815_, _42814_, _42737_);
  not (_42816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_42817_, _42737_, _42816_);
  or (_02825_, _42817_, _42815_);
  not (_42818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_42819_, _42737_, _42818_);
  and (_42820_, _42737_, _42720_);
  or (_02827_, _42820_, _42819_);
  and (_42821_, _42747_, _42244_);
  and (_42822_, _42723_, _42409_);
  and (_42823_, _42822_, _42734_);
  and (_42824_, _42823_, _42821_);
  not (_42825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_42826_, _42823_, _42825_);
  or (_02835_, _42826_, _42824_);
  and (_42828_, _42760_, _42244_);
  and (_42829_, _42823_, _42828_);
  not (_42831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_42833_, _42823_, _42831_);
  or (_02838_, _42833_, _42829_);
  and (_42835_, _42773_, _42244_);
  and (_42837_, _42823_, _42835_);
  not (_42839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_42841_, _42823_, _42839_);
  or (_02841_, _42841_, _42837_);
  and (_42842_, _42781_, _42244_);
  and (_42843_, _42823_, _42842_);
  not (_42844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_42845_, _42823_, _42844_);
  or (_02845_, _42845_, _42843_);
  and (_42846_, _42794_, _42244_);
  and (_42847_, _42823_, _42846_);
  not (_42848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_42849_, _42823_, _42848_);
  or (_02849_, _42849_, _42847_);
  and (_42850_, _42803_, _42244_);
  and (_42851_, _42823_, _42850_);
  not (_42852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_42853_, _42823_, _42852_);
  or (_02852_, _42853_, _42851_);
  and (_42854_, _42814_, _42244_);
  and (_42855_, _42823_, _42854_);
  not (_42856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_42857_, _42823_, _42856_);
  or (_02855_, _42857_, _42855_);
  and (_42858_, _42823_, _42730_);
  nor (_42859_, _42823_, _42656_);
  or (_02858_, _42859_, _42858_);
  and (_42860_, _42724_, _42489_);
  and (_42861_, _42860_, _42734_);
  and (_42862_, _42861_, _42821_);
  not (_42863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_42864_, _42861_, _42863_);
  or (_02864_, _42864_, _42862_);
  and (_42865_, _42861_, _42828_);
  not (_42866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_42867_, _42861_, _42866_);
  or (_02868_, _42867_, _42865_);
  and (_42868_, _42861_, _42835_);
  not (_42869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_42871_, _42861_, _42869_);
  or (_02871_, _42871_, _42868_);
  and (_42874_, _42861_, _42842_);
  not (_42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_42878_, _42861_, _42876_);
  or (_02875_, _42878_, _42874_);
  and (_42881_, _42861_, _42846_);
  not (_42883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_42884_, _42861_, _42883_);
  or (_02878_, _42884_, _42881_);
  and (_42887_, _42861_, _42850_);
  not (_42888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_42889_, _42861_, _42888_);
  or (_02882_, _42889_, _42887_);
  and (_42890_, _42861_, _42854_);
  not (_42891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_42892_, _42861_, _42891_);
  or (_02885_, _42892_, _42890_);
  and (_42893_, _42861_, _42730_);
  not (_42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_42895_, _42861_, _42894_);
  or (_02888_, _42895_, _42893_);
  and (_42896_, _42734_, _42725_);
  and (_42897_, _42896_, _42821_);
  not (_42898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_42899_, _42896_, _42898_);
  or (_02894_, _42899_, _42897_);
  and (_42900_, _42896_, _42828_);
  not (_42901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_42902_, _42896_, _42901_);
  or (_02898_, _42902_, _42900_);
  and (_42903_, _42896_, _42835_);
  not (_42904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_42905_, _42896_, _42904_);
  or (_02902_, _42905_, _42903_);
  and (_42906_, _42896_, _42842_);
  not (_42907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_42908_, _42896_, _42907_);
  or (_02905_, _42908_, _42906_);
  and (_42909_, _42896_, _42846_);
  not (_42910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_42911_, _42896_, _42910_);
  or (_02909_, _42911_, _42909_);
  and (_42912_, _42896_, _42850_);
  not (_42913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_42914_, _42896_, _42913_);
  or (_02912_, _42914_, _42912_);
  and (_42915_, _42896_, _42854_);
  not (_42916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_42917_, _42896_, _42916_);
  or (_02916_, _42917_, _42915_);
  and (_42918_, _42896_, _42730_);
  nor (_42919_, _42896_, _42650_);
  or (_02919_, _42919_, _42918_);
  and (_42920_, _42727_, _42534_);
  and (_42921_, _42920_, _42735_);
  and (_42922_, _42921_, _42821_);
  not (_42923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_42924_, _42921_, _42923_);
  or (_02926_, _42924_, _42922_);
  and (_42925_, _42921_, _42828_);
  not (_42926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_42927_, _42921_, _42926_);
  or (_02929_, _42927_, _42925_);
  and (_42928_, _42921_, _42835_);
  not (_42929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_42930_, _42921_, _42929_);
  or (_02933_, _42930_, _42928_);
  and (_42931_, _42921_, _42842_);
  not (_42932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_42933_, _42921_, _42932_);
  or (_02937_, _42933_, _42931_);
  and (_42934_, _42921_, _42846_);
  not (_42935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_42936_, _42921_, _42935_);
  or (_02940_, _42936_, _42934_);
  and (_42937_, _42921_, _42850_);
  not (_42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_42939_, _42921_, _42938_);
  or (_02943_, _42939_, _42937_);
  and (_42940_, _42921_, _42854_);
  not (_42941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_42942_, _42921_, _42941_);
  or (_02947_, _42942_, _42940_);
  and (_42943_, _42921_, _42730_);
  not (_42944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_42945_, _42921_, _42944_);
  or (_02950_, _42945_, _42943_);
  and (_42946_, _42920_, _42822_);
  and (_42947_, _42946_, _42821_);
  not (_42948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_42949_, _42946_, _42948_);
  or (_02954_, _42949_, _42947_);
  and (_42950_, _42946_, _42828_);
  not (_42951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_42952_, _42946_, _42951_);
  or (_02957_, _42952_, _42950_);
  and (_42953_, _42946_, _42835_);
  not (_42954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_42955_, _42946_, _42954_);
  or (_02962_, _42955_, _42953_);
  and (_42956_, _42946_, _42842_);
  not (_42957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_42958_, _42946_, _42957_);
  or (_02965_, _42958_, _42956_);
  and (_42959_, _42946_, _42846_);
  not (_42960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_42961_, _42946_, _42960_);
  or (_02968_, _42961_, _42959_);
  and (_42962_, _42946_, _42850_);
  not (_42963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_42964_, _42946_, _42963_);
  or (_02972_, _42964_, _42962_);
  and (_42965_, _42946_, _42854_);
  not (_42966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_42967_, _42946_, _42966_);
  or (_02976_, _42967_, _42965_);
  and (_42968_, _42946_, _42730_);
  nor (_42969_, _42946_, _42669_);
  or (_02978_, _42969_, _42968_);
  and (_42970_, _42920_, _42860_);
  and (_42971_, _42970_, _42821_);
  not (_42972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_42973_, _42970_, _42972_);
  or (_02983_, _42973_, _42971_);
  and (_42974_, _42970_, _42828_);
  not (_42975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_42976_, _42970_, _42975_);
  or (_02987_, _42976_, _42974_);
  and (_42977_, _42970_, _42835_);
  not (_42978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_42979_, _42970_, _42978_);
  or (_02991_, _42979_, _42977_);
  and (_42980_, _42970_, _42842_);
  not (_42981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_42982_, _42970_, _42981_);
  or (_02994_, _42982_, _42980_);
  and (_42983_, _42970_, _42846_);
  not (_42984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_42985_, _42970_, _42984_);
  or (_02999_, _42985_, _42983_);
  and (_42986_, _42970_, _42850_);
  not (_42987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_42988_, _42970_, _42987_);
  or (_03002_, _42988_, _42986_);
  and (_42989_, _42970_, _42854_);
  not (_42990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_42991_, _42970_, _42990_);
  or (_03006_, _42991_, _42989_);
  and (_42992_, _42970_, _42730_);
  not (_42993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_42994_, _42970_, _42993_);
  or (_03009_, _42994_, _42992_);
  and (_42995_, _42920_, _42725_);
  and (_42996_, _42995_, _42821_);
  not (_42997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_42998_, _42995_, _42997_);
  or (_03014_, _42998_, _42996_);
  and (_42999_, _42995_, _42828_);
  not (_43000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_43001_, _42995_, _43000_);
  or (_03018_, _43001_, _42999_);
  and (_43002_, _42995_, _42835_);
  not (_43003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_43004_, _42995_, _43003_);
  or (_03021_, _43004_, _43002_);
  and (_43005_, _42995_, _42842_);
  not (_43006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_43007_, _42995_, _43006_);
  or (_03025_, _43007_, _43005_);
  and (_43008_, _42995_, _42846_);
  not (_43009_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_43010_, _42995_, _43009_);
  or (_03028_, _43010_, _43008_);
  and (_43011_, _42995_, _42850_);
  not (_43012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_43013_, _42995_, _43012_);
  or (_03032_, _43013_, _43011_);
  and (_43014_, _42995_, _42854_);
  not (_43015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_43016_, _42995_, _43015_);
  or (_03036_, _43016_, _43014_);
  and (_43017_, _42995_, _42730_);
  nor (_43018_, _42995_, _42663_);
  or (_03038_, _43018_, _43017_);
  and (_43019_, _42726_, _42615_);
  and (_43020_, _43019_, _42735_);
  and (_43021_, _43020_, _42821_);
  not (_43022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_43023_, _43020_, _43022_);
  or (_03045_, _43023_, _43021_);
  and (_43024_, _43020_, _42828_);
  not (_43025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_43026_, _43020_, _43025_);
  or (_03048_, _43026_, _43024_);
  and (_43027_, _43020_, _42835_);
  not (_43028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_43029_, _43020_, _43028_);
  or (_03051_, _43029_, _43027_);
  and (_43030_, _43020_, _42842_);
  not (_43031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_43032_, _43020_, _43031_);
  or (_03054_, _43032_, _43030_);
  and (_43033_, _43020_, _42846_);
  not (_43034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_43035_, _43020_, _43034_);
  or (_03058_, _43035_, _43033_);
  and (_43036_, _43020_, _42850_);
  not (_43037_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_43038_, _43020_, _43037_);
  or (_03061_, _43038_, _43036_);
  and (_43039_, _43020_, _42854_);
  not (_43040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_43041_, _43020_, _43040_);
  or (_03064_, _43041_, _43039_);
  and (_43042_, _43020_, _42730_);
  nor (_43043_, _43020_, _42678_);
  or (_03067_, _43043_, _43042_);
  and (_43044_, _43019_, _42822_);
  and (_43045_, _43044_, _42821_);
  not (_43046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_43047_, _43044_, _43046_);
  or (_03071_, _43047_, _43045_);
  and (_43048_, _43044_, _42828_);
  not (_43049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_43050_, _43044_, _43049_);
  or (_03074_, _43050_, _43048_);
  and (_43051_, _43044_, _42835_);
  not (_43052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_43053_, _43044_, _43052_);
  or (_03078_, _43053_, _43051_);
  and (_43054_, _43044_, _42842_);
  not (_43055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_43056_, _43044_, _43055_);
  or (_03081_, _43056_, _43054_);
  and (_43057_, _43044_, _42846_);
  not (_43058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_43059_, _43044_, _43058_);
  or (_03085_, _43059_, _43057_);
  and (_43060_, _43044_, _42850_);
  not (_43061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_43062_, _43044_, _43061_);
  or (_03089_, _43062_, _43060_);
  and (_43063_, _43044_, _42854_);
  not (_43064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_43065_, _43044_, _43064_);
  or (_03093_, _43065_, _43063_);
  and (_43066_, _43044_, _42730_);
  not (_43067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_43068_, _43044_, _43067_);
  or (_03096_, _43068_, _43066_);
  and (_43069_, _43019_, _42860_);
  and (_43070_, _43069_, _42821_);
  not (_43071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_43072_, _43069_, _43071_);
  or (_03101_, _43072_, _43070_);
  and (_43073_, _43069_, _42828_);
  not (_43074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_43075_, _43069_, _43074_);
  or (_03105_, _43075_, _43073_);
  and (_43076_, _43069_, _42835_);
  not (_43077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_43078_, _43069_, _43077_);
  or (_03109_, _43078_, _43076_);
  and (_43079_, _43069_, _42842_);
  not (_43080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_43081_, _43069_, _43080_);
  or (_03113_, _43081_, _43079_);
  and (_43082_, _43069_, _42846_);
  not (_43083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_43084_, _43069_, _43083_);
  or (_03118_, _43084_, _43082_);
  and (_43085_, _43069_, _42850_);
  not (_43086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_43087_, _43069_, _43086_);
  or (_03122_, _43087_, _43085_);
  and (_43088_, _43069_, _42854_);
  not (_43089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_43090_, _43069_, _43089_);
  or (_03126_, _43090_, _43088_);
  and (_43091_, _43069_, _42730_);
  nor (_43092_, _43069_, _42684_);
  or (_03129_, _43092_, _43091_);
  and (_43093_, _43019_, _42725_);
  and (_43094_, _43093_, _42821_);
  not (_43095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_43096_, _43093_, _43095_);
  or (_03134_, _43096_, _43094_);
  and (_43097_, _43093_, _42828_);
  not (_43098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_43099_, _43093_, _43098_);
  or (_03138_, _43099_, _43097_);
  and (_43100_, _43093_, _42835_);
  not (_43101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_43102_, _43093_, _43101_);
  or (_03142_, _43102_, _43100_);
  and (_43103_, _43093_, _42842_);
  not (_43104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_43105_, _43093_, _43104_);
  or (_03146_, _43105_, _43103_);
  and (_43106_, _43093_, _42846_);
  not (_43107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_43108_, _43093_, _43107_);
  or (_03150_, _43108_, _43106_);
  and (_43109_, _43093_, _42850_);
  not (_43110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_43111_, _43093_, _43110_);
  or (_03154_, _43111_, _43109_);
  and (_43112_, _43093_, _42854_);
  not (_43113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_43114_, _43093_, _43113_);
  or (_03158_, _43114_, _43112_);
  and (_43115_, _43093_, _42730_);
  not (_43116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_43117_, _43093_, _43116_);
  or (_03161_, _43117_, _43115_);
  and (_43118_, _42735_, _42728_);
  and (_43119_, _43118_, _42821_);
  not (_43120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_43121_, _43118_, _43120_);
  or (_03167_, _43121_, _43119_);
  and (_43122_, _43118_, _42828_);
  not (_43123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_43124_, _43118_, _43123_);
  or (_03171_, _43124_, _43122_);
  and (_43125_, _43118_, _42835_);
  not (_43126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_43127_, _43118_, _43126_);
  or (_03175_, _43127_, _43125_);
  and (_43128_, _43118_, _42842_);
  not (_43129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_43130_, _43118_, _43129_);
  or (_03179_, _43130_, _43128_);
  and (_43131_, _43118_, _42846_);
  not (_43132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_43133_, _43118_, _43132_);
  or (_03183_, _43133_, _43131_);
  and (_43134_, _43118_, _42850_);
  not (_43135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_43136_, _43118_, _43135_);
  or (_03187_, _43136_, _43134_);
  and (_43137_, _43118_, _42854_);
  not (_43138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_43139_, _43118_, _43138_);
  or (_03191_, _43139_, _43137_);
  and (_43140_, _43118_, _42730_);
  nor (_43141_, _43118_, _42690_);
  or (_03194_, _43141_, _43140_);
  and (_43142_, _42822_, _42728_);
  and (_43143_, _43142_, _42821_);
  not (_43144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_43145_, _43142_, _43144_);
  or (_03199_, _43145_, _43143_);
  and (_43146_, _43142_, _42828_);
  not (_43147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_43148_, _43142_, _43147_);
  or (_03203_, _43148_, _43146_);
  and (_43149_, _43142_, _42835_);
  not (_43150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_43151_, _43142_, _43150_);
  or (_03207_, _43151_, _43149_);
  and (_43152_, _43142_, _42842_);
  not (_43153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_43154_, _43142_, _43153_);
  or (_03211_, _43154_, _43152_);
  and (_43155_, _43142_, _42846_);
  not (_43156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_43157_, _43142_, _43156_);
  or (_03215_, _43157_, _43155_);
  and (_43158_, _43142_, _42850_);
  not (_43159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_43160_, _43142_, _43159_);
  or (_03219_, _43160_, _43158_);
  and (_43161_, _43142_, _42854_);
  not (_43162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_43163_, _43142_, _43162_);
  or (_03223_, _43163_, _43161_);
  and (_43164_, _43142_, _42730_);
  not (_43165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_43166_, _43142_, _43165_);
  or (_03226_, _43166_, _43164_);
  and (_43167_, _42860_, _42728_);
  and (_43168_, _43167_, _42821_);
  not (_43169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_43170_, _43167_, _43169_);
  or (_03231_, _43170_, _43168_);
  and (_43171_, _43167_, _42828_);
  not (_43172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_43173_, _43167_, _43172_);
  or (_03235_, _43173_, _43171_);
  and (_43174_, _43167_, _42835_);
  not (_43175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_43176_, _43167_, _43175_);
  or (_03239_, _43176_, _43174_);
  and (_43177_, _43167_, _42842_);
  not (_43178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_43179_, _43167_, _43178_);
  or (_03243_, _43179_, _43177_);
  and (_43180_, _43167_, _42846_);
  not (_43181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_43182_, _43167_, _43181_);
  or (_03247_, _43182_, _43180_);
  and (_43183_, _43167_, _42850_);
  not (_43184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_43185_, _43167_, _43184_);
  or (_03251_, _43185_, _43183_);
  and (_43186_, _43167_, _42854_);
  not (_43187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_43188_, _43167_, _43187_);
  or (_03255_, _43188_, _43186_);
  and (_43189_, _43167_, _42730_);
  nor (_43190_, _43167_, _42696_);
  or (_03258_, _43190_, _43189_);
  and (_43191_, _42821_, _42729_);
  not (_43192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_43193_, _42729_, _43192_);
  or (_03263_, _43193_, _43191_);
  and (_43194_, _42828_, _42729_);
  not (_43195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_43196_, _42729_, _43195_);
  or (_03267_, _43196_, _43194_);
  and (_43197_, _42835_, _42729_);
  not (_43198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_43199_, _42729_, _43198_);
  or (_03271_, _43199_, _43197_);
  and (_43200_, _42842_, _42729_);
  not (_43201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_43202_, _42729_, _43201_);
  or (_03275_, _43202_, _43200_);
  and (_43203_, _42846_, _42729_);
  not (_43204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_43205_, _42729_, _43204_);
  or (_03279_, _43205_, _43203_);
  and (_43206_, _42850_, _42729_);
  not (_43207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_43208_, _42729_, _43207_);
  or (_03283_, _43208_, _43206_);
  and (_43209_, _42854_, _42729_);
  not (_43210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_43211_, _42729_, _43210_);
  or (_03287_, _43211_, _43209_);
  nor (_43212_, _42486_, _42898_);
  and (_43213_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_43214_, _43213_, _42404_);
  or (_43215_, _43214_, _43212_);
  and (_43216_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_43217_, _42486_, _42825_);
  nand (_43218_, _43217_, _42404_);
  or (_43219_, _43218_, _43216_);
  and (_43220_, _43219_, _43215_);
  or (_43221_, _43220_, _42649_);
  nor (_43222_, _42486_, _42997_);
  and (_43223_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_43224_, _43223_, _42404_);
  or (_43225_, _43224_, _43222_);
  and (_43226_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_43227_, _42486_, _42948_);
  nand (_43228_, _43227_, _42404_);
  or (_43229_, _43228_, _43226_);
  and (_43230_, _43229_, _43225_);
  or (_43231_, _43230_, _42612_);
  and (_43232_, _43231_, _42662_);
  and (_43233_, _43232_, _43221_);
  nand (_43234_, _42486_, _43022_);
  or (_43235_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_43236_, _43235_, _43234_);
  or (_43237_, _43236_, _42677_);
  or (_43238_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand (_43239_, _42486_, _43071_);
  and (_43240_, _43239_, _43238_);
  or (_43241_, _43240_, _42404_);
  and (_43242_, _43241_, _43237_);
  or (_43243_, _43242_, _42649_);
  nand (_43244_, _42486_, _43120_);
  or (_43245_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_43246_, _43245_, _43244_);
  or (_43247_, _43246_, _42677_);
  or (_43248_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand (_43249_, _42486_, _43169_);
  and (_43250_, _43249_, _43248_);
  or (_43251_, _43250_, _42404_);
  and (_43252_, _43251_, _43247_);
  or (_43253_, _43252_, _42612_);
  and (_43254_, _43253_, _42530_);
  and (_43255_, _43254_, _43243_);
  or (_43256_, _43255_, _43233_);
  or (_43257_, _43256_, _42648_);
  not (_43258_, _42648_);
  or (_43259_, _43258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_43260_, _43259_, _42711_);
  and (_43261_, _43260_, _43257_);
  and (_40036_, _42747_, _42882_);
  and (_43262_, _40036_, _42707_);
  or (_05081_, _43262_, _43261_);
  nor (_43263_, _42486_, _42901_);
  and (_43264_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_43265_, _43264_, _42404_);
  or (_43266_, _43265_, _43263_);
  and (_43267_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_43268_, _42486_, _42831_);
  nand (_43269_, _43268_, _42404_);
  or (_43270_, _43269_, _43267_);
  and (_43271_, _43270_, _43266_);
  or (_43272_, _43271_, _42649_);
  nor (_43273_, _42486_, _43000_);
  and (_43274_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_43275_, _43274_, _42404_);
  or (_43276_, _43275_, _43273_);
  and (_43277_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_43278_, _42486_, _42951_);
  nand (_43279_, _43278_, _42404_);
  or (_43280_, _43279_, _43277_);
  and (_43281_, _43280_, _43276_);
  or (_43282_, _43281_, _42612_);
  and (_43283_, _43282_, _42662_);
  and (_43284_, _43283_, _43272_);
  nand (_43285_, _42486_, _43025_);
  or (_43286_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_43287_, _43286_, _43285_);
  or (_43288_, _43287_, _42677_);
  or (_43289_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand (_43290_, _42486_, _43074_);
  and (_43291_, _43290_, _43289_);
  or (_43292_, _43291_, _42404_);
  and (_43293_, _43292_, _43288_);
  or (_43294_, _43293_, _42649_);
  nand (_43295_, _42486_, _43123_);
  or (_43296_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_43297_, _43296_, _43295_);
  or (_43298_, _43297_, _42677_);
  or (_43299_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand (_43300_, _42486_, _43172_);
  and (_43301_, _43300_, _43299_);
  or (_43302_, _43301_, _42404_);
  and (_43303_, _43302_, _43298_);
  or (_43304_, _43303_, _42612_);
  and (_43305_, _43304_, _42530_);
  and (_43306_, _43305_, _43294_);
  nor (_43307_, _43306_, _43284_);
  nor (_43308_, _43307_, _42648_);
  and (_43309_, _42648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or (_43310_, _43309_, _42707_);
  or (_43311_, _43310_, _43308_);
  and (_40037_, _42760_, _42882_);
  or (_43312_, _40037_, _42711_);
  and (_05083_, _43312_, _43311_);
  or (_43313_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_43314_, _42486_, _43175_);
  and (_43315_, _43314_, _43313_);
  or (_43316_, _43315_, _42404_);
  nand (_43317_, _42486_, _43126_);
  or (_43318_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_43319_, _43318_, _43317_);
  or (_43320_, _43319_, _42677_);
  and (_43321_, _43320_, _42530_);
  and (_43322_, _43321_, _43316_);
  and (_43323_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_43331_, _42486_, _42954_);
  or (_43337_, _43331_, _42677_);
  or (_43341_, _43337_, _43323_);
  nor (_43348_, _42486_, _43003_);
  and (_43356_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_43360_, _43356_, _42404_);
  or (_43365_, _43360_, _43348_);
  and (_43373_, _43365_, _42662_);
  and (_43379_, _43373_, _43341_);
  or (_43383_, _43379_, _43322_);
  and (_43390_, _43383_, _42649_);
  or (_43398_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_43402_, _42486_, _43077_);
  and (_43407_, _43402_, _43398_);
  or (_43415_, _43407_, _42404_);
  nand (_43416_, _42486_, _43028_);
  or (_43424_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_43433_, _43424_, _43416_);
  or (_43439_, _43433_, _42677_);
  and (_43443_, _43439_, _42530_);
  and (_43450_, _43443_, _43415_);
  and (_43458_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_43462_, _42486_, _42839_);
  or (_43467_, _43462_, _42677_);
  or (_43475_, _43467_, _43458_);
  nor (_43481_, _42486_, _42904_);
  and (_43485_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_43492_, _43485_, _42404_);
  or (_43500_, _43492_, _43481_);
  and (_43504_, _43500_, _42662_);
  and (_43509_, _43504_, _43475_);
  or (_43517_, _43509_, _43450_);
  and (_43518_, _43517_, _42612_);
  or (_43519_, _43518_, _42622_);
  or (_43520_, _43519_, _43390_);
  or (_43521_, _43258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_40039_, _42773_, _42882_);
  or (_43522_, _40039_, _42711_);
  and (_43523_, _43522_, _43521_);
  and (_05084_, _43523_, _43520_);
  nor (_43524_, _42486_, _42907_);
  and (_43525_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_43526_, _43525_, _42404_);
  or (_43527_, _43526_, _43524_);
  and (_43528_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_43529_, _42486_, _42844_);
  nand (_43530_, _43529_, _42404_);
  or (_43531_, _43530_, _43528_);
  and (_43532_, _43531_, _43527_);
  or (_43533_, _43532_, _42649_);
  nor (_43534_, _42486_, _43006_);
  and (_43535_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_43536_, _43535_, _42404_);
  or (_43537_, _43536_, _43534_);
  and (_43538_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_43539_, _42486_, _42957_);
  nand (_43540_, _43539_, _42404_);
  or (_43541_, _43540_, _43538_);
  and (_43542_, _43541_, _43537_);
  or (_43543_, _43542_, _42612_);
  and (_43544_, _43543_, _42662_);
  and (_43545_, _43544_, _43533_);
  nand (_43546_, _42486_, _43031_);
  or (_43547_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_43548_, _43547_, _43546_);
  or (_43549_, _43548_, _42677_);
  or (_43550_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_43551_, _42486_, _43080_);
  and (_43552_, _43551_, _43550_);
  or (_43553_, _43552_, _42404_);
  and (_43554_, _43553_, _43549_);
  or (_43555_, _43554_, _42649_);
  nand (_43556_, _42486_, _43129_);
  or (_43557_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_43558_, _43557_, _43556_);
  or (_43559_, _43558_, _42677_);
  or (_43560_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_43561_, _42486_, _43178_);
  and (_43562_, _43561_, _43560_);
  or (_43563_, _43562_, _42404_);
  and (_43564_, _43563_, _43559_);
  or (_43565_, _43564_, _42612_);
  and (_43566_, _43565_, _42530_);
  and (_43567_, _43566_, _43555_);
  nor (_43568_, _43567_, _43545_);
  nor (_43569_, _43568_, _42648_);
  and (_43570_, _42648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_43571_, _43570_, _42707_);
  or (_43572_, _43571_, _43569_);
  and (_40040_, _42781_, _42882_);
  or (_43573_, _40040_, _42711_);
  and (_05086_, _43573_, _43572_);
  and (_43574_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_43575_, _42486_, _42848_);
  nand (_43576_, _43575_, _42404_);
  or (_43577_, _43576_, _43574_);
  nor (_43578_, _42486_, _42910_);
  and (_43579_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_43580_, _43579_, _42404_);
  or (_43581_, _43580_, _43578_);
  and (_43582_, _43581_, _43577_);
  or (_43583_, _43582_, _42649_);
  nor (_43584_, _42486_, _43009_);
  and (_43585_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_43586_, _43585_, _42404_);
  or (_43587_, _43586_, _43584_);
  and (_43588_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_43589_, _42486_, _42960_);
  nand (_43590_, _43589_, _42404_);
  or (_43591_, _43590_, _43588_);
  and (_43592_, _43591_, _43587_);
  or (_43593_, _43592_, _42612_);
  and (_43594_, _43593_, _42662_);
  and (_43595_, _43594_, _43583_);
  nor (_43596_, _42486_, _43107_);
  and (_43597_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_43598_, _43597_, _42404_);
  or (_43599_, _43598_, _43596_);
  and (_43600_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_43601_, _42486_, _43058_);
  nand (_43602_, _43601_, _42404_);
  or (_43603_, _43602_, _43600_);
  and (_43604_, _43603_, _43599_);
  or (_43605_, _43604_, _42649_);
  nor (_43606_, _42486_, _43204_);
  and (_43607_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_43608_, _43607_, _42404_);
  or (_43609_, _43608_, _43606_);
  and (_43610_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_43611_, _42486_, _43156_);
  nand (_43612_, _43611_, _42404_);
  or (_43613_, _43612_, _43610_);
  and (_43614_, _43613_, _43609_);
  or (_43615_, _43614_, _42612_);
  and (_43616_, _43615_, _42530_);
  and (_43617_, _43616_, _43605_);
  or (_43618_, _43617_, _43595_);
  and (_43619_, _43618_, _42706_);
  and (_43620_, _42794_, _42707_);
  and (_43621_, _42648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or (_43622_, _43621_, _43620_);
  or (_43623_, _43622_, _43619_);
  and (_05088_, _43623_, _42882_);
  nor (_43624_, _42486_, _42913_);
  and (_43625_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_43626_, _43625_, _42404_);
  or (_43627_, _43626_, _43624_);
  and (_43628_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_43629_, _42486_, _42852_);
  nand (_43630_, _43629_, _42404_);
  or (_43631_, _43630_, _43628_);
  and (_43632_, _43631_, _43627_);
  or (_43633_, _43632_, _42649_);
  nor (_43634_, _42486_, _43012_);
  and (_43635_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_43636_, _43635_, _42404_);
  or (_43637_, _43636_, _43634_);
  and (_43638_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_43639_, _42486_, _42963_);
  nand (_43640_, _43639_, _42404_);
  or (_43641_, _43640_, _43638_);
  and (_43642_, _43641_, _43637_);
  or (_43643_, _43642_, _42612_);
  and (_43644_, _43643_, _42662_);
  and (_43645_, _43644_, _43633_);
  nand (_43646_, _42486_, _43037_);
  or (_43647_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_43648_, _43647_, _43646_);
  or (_43649_, _43648_, _42677_);
  or (_43650_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_43651_, _42486_, _43086_);
  and (_43652_, _43651_, _43650_);
  or (_43653_, _43652_, _42404_);
  and (_43654_, _43653_, _43649_);
  or (_43655_, _43654_, _42649_);
  nand (_43656_, _42486_, _43135_);
  or (_43657_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_43658_, _43657_, _43656_);
  or (_43659_, _43658_, _42677_);
  or (_43660_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_43661_, _42486_, _43184_);
  and (_43662_, _43661_, _43660_);
  or (_43663_, _43662_, _42404_);
  and (_43664_, _43663_, _43659_);
  or (_43665_, _43664_, _42612_);
  and (_43666_, _43665_, _42530_);
  and (_43667_, _43666_, _43655_);
  or (_43668_, _43667_, _43645_);
  or (_43669_, _43668_, _42648_);
  or (_43670_, _43258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_43671_, _43670_, _42711_);
  and (_43672_, _43671_, _43669_);
  and (_40042_, _42803_, _42882_);
  and (_43673_, _40042_, _42707_);
  or (_05090_, _43673_, _43672_);
  nor (_43674_, _42486_, _42916_);
  and (_43675_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_43676_, _43675_, _42404_);
  or (_43677_, _43676_, _43674_);
  and (_43678_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_43679_, _42486_, _42856_);
  nand (_43680_, _43679_, _42404_);
  or (_43681_, _43680_, _43678_);
  and (_43682_, _43681_, _43677_);
  or (_43683_, _43682_, _42649_);
  nor (_43684_, _42486_, _43015_);
  and (_43685_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_43686_, _43685_, _42404_);
  or (_43687_, _43686_, _43684_);
  and (_43688_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_43689_, _42486_, _42966_);
  nand (_43690_, _43689_, _42404_);
  or (_43691_, _43690_, _43688_);
  and (_43692_, _43691_, _43687_);
  or (_43693_, _43692_, _42612_);
  and (_43694_, _43693_, _42662_);
  and (_43695_, _43694_, _43683_);
  nand (_43696_, _42486_, _43040_);
  or (_43697_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_43698_, _43697_, _43696_);
  or (_43699_, _43698_, _42677_);
  or (_43700_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_43701_, _42486_, _43089_);
  and (_43702_, _43701_, _43700_);
  or (_43703_, _43702_, _42404_);
  and (_43704_, _43703_, _43699_);
  or (_43705_, _43704_, _42649_);
  nand (_43706_, _42486_, _43138_);
  or (_43707_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_43708_, _43707_, _43706_);
  or (_43709_, _43708_, _42677_);
  or (_43710_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_43711_, _42486_, _43187_);
  and (_43712_, _43711_, _43710_);
  or (_43713_, _43712_, _42404_);
  and (_43714_, _43713_, _43709_);
  or (_43715_, _43714_, _42612_);
  and (_43716_, _43715_, _42530_);
  and (_43717_, _43716_, _43705_);
  or (_43718_, _43717_, _43695_);
  or (_43719_, _43718_, _42648_);
  or (_43720_, _43258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_43721_, _43720_, _42711_);
  and (_43722_, _43721_, _43719_);
  and (_40043_, _42814_, _42882_);
  and (_43723_, _40043_, _42707_);
  or (_05092_, _43723_, _43722_);
  or (_43724_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_43725_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_43726_, _43725_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_43727_, _43726_, _43724_);
  nand (_43728_, _43727_, _42882_);
  or (_43729_, \oc8051_gm_cxrom_1.cell0.data [7], _42882_);
  and (_05100_, _43729_, _43728_);
  or (_43730_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43731_, \oc8051_gm_cxrom_1.cell0.data [0], _43725_);
  nand (_43732_, _43731_, _43730_);
  nand (_43733_, _43732_, _42882_);
  or (_43734_, \oc8051_gm_cxrom_1.cell0.data [0], _42882_);
  and (_05107_, _43734_, _43733_);
  or (_43735_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43736_, \oc8051_gm_cxrom_1.cell0.data [1], _43725_);
  nand (_43737_, _43736_, _43735_);
  nand (_43738_, _43737_, _42882_);
  or (_43739_, \oc8051_gm_cxrom_1.cell0.data [1], _42882_);
  and (_05111_, _43739_, _43738_);
  or (_43740_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43741_, \oc8051_gm_cxrom_1.cell0.data [2], _43725_);
  nand (_43742_, _43741_, _43740_);
  nand (_43743_, _43742_, _42882_);
  or (_43744_, \oc8051_gm_cxrom_1.cell0.data [2], _42882_);
  and (_05115_, _43744_, _43743_);
  or (_43745_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43746_, \oc8051_gm_cxrom_1.cell0.data [3], _43725_);
  nand (_43747_, _43746_, _43745_);
  nand (_43748_, _43747_, _42882_);
  or (_43749_, \oc8051_gm_cxrom_1.cell0.data [3], _42882_);
  and (_05119_, _43749_, _43748_);
  or (_43750_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43751_, \oc8051_gm_cxrom_1.cell0.data [4], _43725_);
  nand (_43752_, _43751_, _43750_);
  nand (_43753_, _43752_, _42882_);
  or (_43754_, \oc8051_gm_cxrom_1.cell0.data [4], _42882_);
  and (_05123_, _43754_, _43753_);
  nor (_43755_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  nor (_43756_, \oc8051_gm_cxrom_1.cell0.data [5], _43725_);
  or (_43757_, _43756_, _43755_);
  nand (_43758_, _43757_, _42882_);
  or (_43759_, \oc8051_gm_cxrom_1.cell0.data [5], _42882_);
  and (_05126_, _43759_, _43758_);
  or (_43760_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43761_, \oc8051_gm_cxrom_1.cell0.data [6], _43725_);
  nand (_43762_, _43761_, _43760_);
  nand (_43763_, _43762_, _42882_);
  or (_43764_, \oc8051_gm_cxrom_1.cell0.data [6], _42882_);
  and (_05130_, _43764_, _43763_);
  or (_43765_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_43766_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_43767_, _43766_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_43768_, _43767_, _43765_);
  nand (_43769_, _43768_, _42882_);
  or (_43770_, \oc8051_gm_cxrom_1.cell1.data [7], _42882_);
  and (_05152_, _43770_, _43769_);
  or (_43771_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43772_, \oc8051_gm_cxrom_1.cell1.data [0], _43766_);
  nand (_43773_, _43772_, _43771_);
  nand (_43774_, _43773_, _42882_);
  or (_43775_, \oc8051_gm_cxrom_1.cell1.data [0], _42882_);
  and (_05159_, _43775_, _43774_);
  or (_43776_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43777_, \oc8051_gm_cxrom_1.cell1.data [1], _43766_);
  nand (_43778_, _43777_, _43776_);
  nand (_43779_, _43778_, _42882_);
  or (_43780_, \oc8051_gm_cxrom_1.cell1.data [1], _42882_);
  and (_05162_, _43780_, _43779_);
  or (_43781_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43782_, \oc8051_gm_cxrom_1.cell1.data [2], _43766_);
  nand (_43783_, _43782_, _43781_);
  nand (_43784_, _43783_, _42882_);
  or (_43785_, \oc8051_gm_cxrom_1.cell1.data [2], _42882_);
  and (_05166_, _43785_, _43784_);
  or (_43786_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43787_, \oc8051_gm_cxrom_1.cell1.data [3], _43766_);
  nand (_43788_, _43787_, _43786_);
  nand (_43789_, _43788_, _42882_);
  or (_43790_, \oc8051_gm_cxrom_1.cell1.data [3], _42882_);
  and (_05170_, _43790_, _43789_);
  or (_43791_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43792_, \oc8051_gm_cxrom_1.cell1.data [4], _43766_);
  nand (_43793_, _43792_, _43791_);
  nand (_43794_, _43793_, _42882_);
  or (_43795_, \oc8051_gm_cxrom_1.cell1.data [4], _42882_);
  and (_05174_, _43795_, _43794_);
  nor (_43796_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  nor (_43797_, \oc8051_gm_cxrom_1.cell1.data [5], _43766_);
  or (_43798_, _43797_, _43796_);
  nand (_43799_, _43798_, _42882_);
  or (_43800_, \oc8051_gm_cxrom_1.cell1.data [5], _42882_);
  and (_05178_, _43800_, _43799_);
  or (_43801_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43802_, \oc8051_gm_cxrom_1.cell1.data [6], _43766_);
  nand (_43803_, _43802_, _43801_);
  nand (_43804_, _43803_, _42882_);
  or (_43805_, \oc8051_gm_cxrom_1.cell1.data [6], _42882_);
  and (_05182_, _43805_, _43804_);
  or (_43806_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_43807_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_43808_, _43807_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_43809_, _43808_, _43806_);
  nand (_43810_, _43809_, _42882_);
  or (_43811_, \oc8051_gm_cxrom_1.cell2.data [7], _42882_);
  and (_05203_, _43811_, _43810_);
  or (_00002_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00003_, \oc8051_gm_cxrom_1.cell2.data [0], _43807_);
  nand (_00004_, _00003_, _00002_);
  nand (_00005_, _00004_, _42882_);
  or (_00006_, \oc8051_gm_cxrom_1.cell2.data [0], _42882_);
  and (_05210_, _00006_, _00005_);
  or (_00007_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00008_, \oc8051_gm_cxrom_1.cell2.data [1], _43807_);
  nand (_00009_, _00008_, _00007_);
  nand (_00010_, _00009_, _42882_);
  or (_00011_, \oc8051_gm_cxrom_1.cell2.data [1], _42882_);
  and (_05214_, _00011_, _00010_);
  or (_00012_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00013_, \oc8051_gm_cxrom_1.cell2.data [2], _43807_);
  nand (_00014_, _00013_, _00012_);
  nand (_00015_, _00014_, _42882_);
  or (_00016_, \oc8051_gm_cxrom_1.cell2.data [2], _42882_);
  and (_05218_, _00016_, _00015_);
  or (_00017_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00018_, \oc8051_gm_cxrom_1.cell2.data [3], _43807_);
  nand (_00019_, _00018_, _00017_);
  nand (_00020_, _00019_, _42882_);
  or (_00021_, \oc8051_gm_cxrom_1.cell2.data [3], _42882_);
  and (_05222_, _00021_, _00020_);
  or (_00022_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00023_, \oc8051_gm_cxrom_1.cell2.data [4], _43807_);
  nand (_00024_, _00023_, _00022_);
  nand (_00025_, _00024_, _42882_);
  or (_00026_, \oc8051_gm_cxrom_1.cell2.data [4], _42882_);
  and (_05226_, _00026_, _00025_);
  nor (_00027_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  nor (_00028_, \oc8051_gm_cxrom_1.cell2.data [5], _43807_);
  or (_00029_, _00028_, _00027_);
  nand (_00030_, _00029_, _42882_);
  or (_00031_, \oc8051_gm_cxrom_1.cell2.data [5], _42882_);
  and (_05230_, _00031_, _00030_);
  or (_00032_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00033_, \oc8051_gm_cxrom_1.cell2.data [6], _43807_);
  nand (_00034_, _00033_, _00032_);
  nand (_00035_, _00034_, _42882_);
  or (_00036_, \oc8051_gm_cxrom_1.cell2.data [6], _42882_);
  and (_05234_, _00036_, _00035_);
  or (_00037_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_00038_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_00039_, _00038_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_00040_, _00039_, _00037_);
  nand (_00041_, _00040_, _42882_);
  or (_00042_, \oc8051_gm_cxrom_1.cell3.data [7], _42882_);
  and (_05255_, _00042_, _00041_);
  or (_00043_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00044_, \oc8051_gm_cxrom_1.cell3.data [0], _00038_);
  nand (_00045_, _00044_, _00043_);
  nand (_00046_, _00045_, _42882_);
  or (_00047_, \oc8051_gm_cxrom_1.cell3.data [0], _42882_);
  and (_05262_, _00047_, _00046_);
  or (_00048_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00049_, \oc8051_gm_cxrom_1.cell3.data [1], _00038_);
  nand (_00050_, _00049_, _00048_);
  nand (_00051_, _00050_, _42882_);
  or (_00052_, \oc8051_gm_cxrom_1.cell3.data [1], _42882_);
  and (_05266_, _00052_, _00051_);
  or (_00053_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00054_, \oc8051_gm_cxrom_1.cell3.data [2], _00038_);
  nand (_00055_, _00054_, _00053_);
  nand (_00056_, _00055_, _42882_);
  or (_00057_, \oc8051_gm_cxrom_1.cell3.data [2], _42882_);
  and (_05270_, _00057_, _00056_);
  or (_00058_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00059_, \oc8051_gm_cxrom_1.cell3.data [3], _00038_);
  nand (_00060_, _00059_, _00058_);
  nand (_00061_, _00060_, _42882_);
  or (_00062_, \oc8051_gm_cxrom_1.cell3.data [3], _42882_);
  and (_05273_, _00062_, _00061_);
  or (_00063_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00064_, \oc8051_gm_cxrom_1.cell3.data [4], _00038_);
  nand (_00065_, _00064_, _00063_);
  nand (_00066_, _00065_, _42882_);
  or (_00067_, \oc8051_gm_cxrom_1.cell3.data [4], _42882_);
  and (_05277_, _00067_, _00066_);
  nor (_00068_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  nor (_00069_, \oc8051_gm_cxrom_1.cell3.data [5], _00038_);
  or (_00070_, _00069_, _00068_);
  nand (_00071_, _00070_, _42882_);
  or (_00072_, \oc8051_gm_cxrom_1.cell3.data [5], _42882_);
  and (_05281_, _00072_, _00071_);
  or (_00073_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00074_, \oc8051_gm_cxrom_1.cell3.data [6], _00038_);
  nand (_00075_, _00074_, _00073_);
  nand (_00076_, _00075_, _42882_);
  or (_00077_, \oc8051_gm_cxrom_1.cell3.data [6], _42882_);
  and (_05285_, _00077_, _00076_);
  or (_00078_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_00079_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_00080_, _00079_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_00081_, _00080_, _00078_);
  nand (_00082_, _00081_, _42882_);
  or (_00083_, \oc8051_gm_cxrom_1.cell4.data [7], _42882_);
  and (_05306_, _00083_, _00082_);
  or (_00084_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00085_, \oc8051_gm_cxrom_1.cell4.data [0], _00079_);
  nand (_00086_, _00085_, _00084_);
  nand (_00087_, _00086_, _42882_);
  or (_00088_, \oc8051_gm_cxrom_1.cell4.data [0], _42882_);
  and (_05313_, _00088_, _00087_);
  or (_00089_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00090_, \oc8051_gm_cxrom_1.cell4.data [1], _00079_);
  nand (_00091_, _00090_, _00089_);
  nand (_00092_, _00091_, _42882_);
  or (_00093_, \oc8051_gm_cxrom_1.cell4.data [1], _42882_);
  and (_05317_, _00093_, _00092_);
  or (_00094_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00095_, \oc8051_gm_cxrom_1.cell4.data [2], _00079_);
  nand (_00096_, _00095_, _00094_);
  nand (_00097_, _00096_, _42882_);
  or (_00098_, \oc8051_gm_cxrom_1.cell4.data [2], _42882_);
  and (_05321_, _00098_, _00097_);
  or (_00099_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00100_, \oc8051_gm_cxrom_1.cell4.data [3], _00079_);
  nand (_00101_, _00100_, _00099_);
  nand (_00102_, _00101_, _42882_);
  or (_00103_, \oc8051_gm_cxrom_1.cell4.data [3], _42882_);
  and (_05325_, _00103_, _00102_);
  or (_00104_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00105_, \oc8051_gm_cxrom_1.cell4.data [4], _00079_);
  nand (_00106_, _00105_, _00104_);
  nand (_00107_, _00106_, _42882_);
  or (_00108_, \oc8051_gm_cxrom_1.cell4.data [4], _42882_);
  and (_05329_, _00108_, _00107_);
  nor (_00109_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  nor (_00110_, \oc8051_gm_cxrom_1.cell4.data [5], _00079_);
  or (_00111_, _00110_, _00109_);
  nand (_00112_, _00111_, _42882_);
  or (_00113_, \oc8051_gm_cxrom_1.cell4.data [5], _42882_);
  and (_05333_, _00113_, _00112_);
  or (_00114_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00115_, \oc8051_gm_cxrom_1.cell4.data [6], _00079_);
  nand (_00116_, _00115_, _00114_);
  nand (_00117_, _00116_, _42882_);
  or (_00118_, \oc8051_gm_cxrom_1.cell4.data [6], _42882_);
  and (_05337_, _00118_, _00117_);
  or (_00119_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_00120_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_00121_, _00120_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_00122_, _00121_, _00119_);
  nand (_00123_, _00122_, _42882_);
  or (_00124_, \oc8051_gm_cxrom_1.cell5.data [7], _42882_);
  and (_05359_, _00124_, _00123_);
  or (_00125_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00126_, \oc8051_gm_cxrom_1.cell5.data [0], _00120_);
  nand (_00127_, _00126_, _00125_);
  nand (_00128_, _00127_, _42882_);
  or (_00129_, \oc8051_gm_cxrom_1.cell5.data [0], _42882_);
  and (_05366_, _00129_, _00128_);
  or (_00131_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00133_, \oc8051_gm_cxrom_1.cell5.data [1], _00120_);
  nand (_00135_, _00133_, _00131_);
  nand (_00137_, _00135_, _42882_);
  or (_00139_, \oc8051_gm_cxrom_1.cell5.data [1], _42882_);
  and (_05370_, _00139_, _00137_);
  or (_00142_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00144_, \oc8051_gm_cxrom_1.cell5.data [2], _00120_);
  nand (_00146_, _00144_, _00142_);
  nand (_00148_, _00146_, _42882_);
  or (_00150_, \oc8051_gm_cxrom_1.cell5.data [2], _42882_);
  and (_05374_, _00150_, _00148_);
  or (_00153_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00155_, \oc8051_gm_cxrom_1.cell5.data [3], _00120_);
  nand (_00157_, _00155_, _00153_);
  nand (_00159_, _00157_, _42882_);
  or (_00161_, \oc8051_gm_cxrom_1.cell5.data [3], _42882_);
  and (_05378_, _00161_, _00159_);
  or (_00164_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00166_, \oc8051_gm_cxrom_1.cell5.data [4], _00120_);
  nand (_00168_, _00166_, _00164_);
  nand (_00170_, _00168_, _42882_);
  or (_00172_, \oc8051_gm_cxrom_1.cell5.data [4], _42882_);
  and (_05382_, _00172_, _00170_);
  nor (_00175_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  nor (_00177_, \oc8051_gm_cxrom_1.cell5.data [5], _00120_);
  or (_00179_, _00177_, _00175_);
  nand (_00181_, _00179_, _42882_);
  or (_00183_, \oc8051_gm_cxrom_1.cell5.data [5], _42882_);
  and (_05386_, _00183_, _00181_);
  or (_00186_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00187_, \oc8051_gm_cxrom_1.cell5.data [6], _00120_);
  nand (_00188_, _00187_, _00186_);
  nand (_00189_, _00188_, _42882_);
  or (_00190_, \oc8051_gm_cxrom_1.cell5.data [6], _42882_);
  and (_05390_, _00190_, _00189_);
  or (_00191_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_00192_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_00193_, _00192_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_00194_, _00193_, _00191_);
  nand (_00195_, _00194_, _42882_);
  or (_00196_, \oc8051_gm_cxrom_1.cell6.data [7], _42882_);
  and (_05412_, _00196_, _00195_);
  or (_00197_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00198_, \oc8051_gm_cxrom_1.cell6.data [0], _00192_);
  nand (_00199_, _00198_, _00197_);
  nand (_00200_, _00199_, _42882_);
  or (_00201_, \oc8051_gm_cxrom_1.cell6.data [0], _42882_);
  and (_05419_, _00201_, _00200_);
  or (_00202_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00203_, \oc8051_gm_cxrom_1.cell6.data [1], _00192_);
  nand (_00204_, _00203_, _00202_);
  nand (_00205_, _00204_, _42882_);
  or (_00206_, \oc8051_gm_cxrom_1.cell6.data [1], _42882_);
  and (_05423_, _00206_, _00205_);
  or (_00207_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00208_, \oc8051_gm_cxrom_1.cell6.data [2], _00192_);
  nand (_00209_, _00208_, _00207_);
  nand (_00210_, _00209_, _42882_);
  or (_00211_, \oc8051_gm_cxrom_1.cell6.data [2], _42882_);
  and (_05427_, _00211_, _00210_);
  or (_00212_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00213_, \oc8051_gm_cxrom_1.cell6.data [3], _00192_);
  nand (_00214_, _00213_, _00212_);
  nand (_00215_, _00214_, _42882_);
  or (_00216_, \oc8051_gm_cxrom_1.cell6.data [3], _42882_);
  and (_05431_, _00216_, _00215_);
  or (_00217_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00218_, \oc8051_gm_cxrom_1.cell6.data [4], _00192_);
  nand (_00219_, _00218_, _00217_);
  nand (_00220_, _00219_, _42882_);
  or (_00221_, \oc8051_gm_cxrom_1.cell6.data [4], _42882_);
  and (_05435_, _00221_, _00220_);
  nor (_00222_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  nor (_00223_, \oc8051_gm_cxrom_1.cell6.data [5], _00192_);
  or (_00224_, _00223_, _00222_);
  nand (_00225_, _00224_, _42882_);
  or (_00226_, \oc8051_gm_cxrom_1.cell6.data [5], _42882_);
  and (_05439_, _00226_, _00225_);
  or (_00227_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00228_, \oc8051_gm_cxrom_1.cell6.data [6], _00192_);
  nand (_00229_, _00228_, _00227_);
  nand (_00230_, _00229_, _42882_);
  or (_00231_, \oc8051_gm_cxrom_1.cell6.data [6], _42882_);
  and (_05443_, _00231_, _00230_);
  or (_00232_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_00233_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_00234_, _00233_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_00235_, _00234_, _00232_);
  nand (_00236_, _00235_, _42882_);
  or (_00237_, \oc8051_gm_cxrom_1.cell7.data [7], _42882_);
  and (_05465_, _00237_, _00236_);
  or (_00238_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00239_, \oc8051_gm_cxrom_1.cell7.data [0], _00233_);
  nand (_00240_, _00239_, _00238_);
  nand (_00241_, _00240_, _42882_);
  or (_00242_, \oc8051_gm_cxrom_1.cell7.data [0], _42882_);
  and (_05472_, _00242_, _00241_);
  or (_00243_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00244_, \oc8051_gm_cxrom_1.cell7.data [1], _00233_);
  nand (_00245_, _00244_, _00243_);
  nand (_00246_, _00245_, _42882_);
  or (_00247_, \oc8051_gm_cxrom_1.cell7.data [1], _42882_);
  and (_05476_, _00247_, _00246_);
  or (_00248_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00249_, \oc8051_gm_cxrom_1.cell7.data [2], _00233_);
  nand (_00250_, _00249_, _00248_);
  nand (_00251_, _00250_, _42882_);
  or (_00252_, \oc8051_gm_cxrom_1.cell7.data [2], _42882_);
  and (_05480_, _00252_, _00251_);
  or (_00253_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00254_, \oc8051_gm_cxrom_1.cell7.data [3], _00233_);
  nand (_00255_, _00254_, _00253_);
  nand (_00256_, _00255_, _42882_);
  or (_00257_, \oc8051_gm_cxrom_1.cell7.data [3], _42882_);
  and (_05484_, _00257_, _00256_);
  or (_00258_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00259_, \oc8051_gm_cxrom_1.cell7.data [4], _00233_);
  nand (_00260_, _00259_, _00258_);
  nand (_00261_, _00260_, _42882_);
  or (_00262_, \oc8051_gm_cxrom_1.cell7.data [4], _42882_);
  and (_05488_, _00262_, _00261_);
  nor (_00263_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  nor (_00264_, \oc8051_gm_cxrom_1.cell7.data [5], _00233_);
  or (_00265_, _00264_, _00263_);
  nand (_00266_, _00265_, _42882_);
  or (_00267_, \oc8051_gm_cxrom_1.cell7.data [5], _42882_);
  and (_05492_, _00267_, _00266_);
  or (_00268_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00269_, \oc8051_gm_cxrom_1.cell7.data [6], _00233_);
  nand (_00270_, _00269_, _00268_);
  nand (_00271_, _00270_, _42882_);
  or (_00272_, \oc8051_gm_cxrom_1.cell7.data [6], _42882_);
  and (_05496_, _00272_, _00271_);
  or (_00273_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_00274_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_00275_, _00274_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_00276_, _00275_, _00273_);
  nand (_00277_, _00276_, _42882_);
  or (_00278_, \oc8051_gm_cxrom_1.cell8.data [7], _42882_);
  and (_05518_, _00278_, _00277_);
  or (_00279_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00280_, \oc8051_gm_cxrom_1.cell8.data [0], _00274_);
  nand (_00281_, _00280_, _00279_);
  nand (_00282_, _00281_, _42882_);
  or (_00283_, \oc8051_gm_cxrom_1.cell8.data [0], _42882_);
  and (_05525_, _00283_, _00282_);
  or (_00284_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00285_, \oc8051_gm_cxrom_1.cell8.data [1], _00274_);
  nand (_00286_, _00285_, _00284_);
  nand (_00287_, _00286_, _42882_);
  or (_00288_, \oc8051_gm_cxrom_1.cell8.data [1], _42882_);
  and (_05529_, _00288_, _00287_);
  or (_00289_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00290_, \oc8051_gm_cxrom_1.cell8.data [2], _00274_);
  nand (_00291_, _00290_, _00289_);
  nand (_00292_, _00291_, _42882_);
  or (_00293_, \oc8051_gm_cxrom_1.cell8.data [2], _42882_);
  and (_05533_, _00293_, _00292_);
  or (_00294_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00295_, \oc8051_gm_cxrom_1.cell8.data [3], _00274_);
  nand (_00296_, _00295_, _00294_);
  nand (_00297_, _00296_, _42882_);
  or (_00298_, \oc8051_gm_cxrom_1.cell8.data [3], _42882_);
  and (_05537_, _00298_, _00297_);
  or (_00299_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00300_, \oc8051_gm_cxrom_1.cell8.data [4], _00274_);
  nand (_00301_, _00300_, _00299_);
  nand (_00302_, _00301_, _42882_);
  or (_00303_, \oc8051_gm_cxrom_1.cell8.data [4], _42882_);
  and (_05541_, _00303_, _00302_);
  nor (_00304_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  nor (_00305_, \oc8051_gm_cxrom_1.cell8.data [5], _00274_);
  or (_00306_, _00305_, _00304_);
  nand (_00307_, _00306_, _42882_);
  or (_00308_, \oc8051_gm_cxrom_1.cell8.data [5], _42882_);
  and (_05545_, _00308_, _00307_);
  or (_00309_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00310_, \oc8051_gm_cxrom_1.cell8.data [6], _00274_);
  nand (_00311_, _00310_, _00309_);
  nand (_00312_, _00311_, _42882_);
  or (_00313_, \oc8051_gm_cxrom_1.cell8.data [6], _42882_);
  and (_05549_, _00313_, _00312_);
  or (_00314_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_00315_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_00316_, _00315_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_00317_, _00316_, _00314_);
  nand (_00318_, _00317_, _42882_);
  or (_00319_, \oc8051_gm_cxrom_1.cell9.data [7], _42882_);
  and (_05571_, _00319_, _00318_);
  or (_00320_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00321_, \oc8051_gm_cxrom_1.cell9.data [0], _00315_);
  nand (_00322_, _00321_, _00320_);
  nand (_00323_, _00322_, _42882_);
  or (_00324_, \oc8051_gm_cxrom_1.cell9.data [0], _42882_);
  and (_05578_, _00324_, _00323_);
  or (_00325_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00326_, \oc8051_gm_cxrom_1.cell9.data [1], _00315_);
  nand (_00327_, _00326_, _00325_);
  nand (_00328_, _00327_, _42882_);
  or (_00329_, \oc8051_gm_cxrom_1.cell9.data [1], _42882_);
  and (_05582_, _00329_, _00328_);
  or (_00330_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00331_, \oc8051_gm_cxrom_1.cell9.data [2], _00315_);
  nand (_00332_, _00331_, _00330_);
  nand (_00333_, _00332_, _42882_);
  or (_00334_, \oc8051_gm_cxrom_1.cell9.data [2], _42882_);
  and (_05586_, _00334_, _00333_);
  or (_00335_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00336_, \oc8051_gm_cxrom_1.cell9.data [3], _00315_);
  nand (_00337_, _00336_, _00335_);
  nand (_00338_, _00337_, _42882_);
  or (_00339_, \oc8051_gm_cxrom_1.cell9.data [3], _42882_);
  and (_05590_, _00339_, _00338_);
  or (_00340_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00341_, \oc8051_gm_cxrom_1.cell9.data [4], _00315_);
  nand (_00342_, _00341_, _00340_);
  nand (_00343_, _00342_, _42882_);
  or (_00344_, \oc8051_gm_cxrom_1.cell9.data [4], _42882_);
  and (_05594_, _00344_, _00343_);
  nor (_00345_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  nor (_00346_, \oc8051_gm_cxrom_1.cell9.data [5], _00315_);
  or (_00347_, _00346_, _00345_);
  nand (_00348_, _00347_, _42882_);
  or (_00349_, \oc8051_gm_cxrom_1.cell9.data [5], _42882_);
  and (_05598_, _00349_, _00348_);
  or (_00350_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00351_, \oc8051_gm_cxrom_1.cell9.data [6], _00315_);
  nand (_00352_, _00351_, _00350_);
  nand (_00353_, _00352_, _42882_);
  or (_00354_, \oc8051_gm_cxrom_1.cell9.data [6], _42882_);
  and (_05602_, _00354_, _00353_);
  or (_00355_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_00356_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_00357_, _00356_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_00358_, _00357_, _00355_);
  nand (_00359_, _00358_, _42882_);
  or (_00360_, \oc8051_gm_cxrom_1.cell10.data [7], _42882_);
  and (_05624_, _00360_, _00359_);
  or (_00361_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00362_, \oc8051_gm_cxrom_1.cell10.data [0], _00356_);
  nand (_00363_, _00362_, _00361_);
  nand (_00364_, _00363_, _42882_);
  or (_00365_, \oc8051_gm_cxrom_1.cell10.data [0], _42882_);
  and (_05631_, _00365_, _00364_);
  or (_00366_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00367_, \oc8051_gm_cxrom_1.cell10.data [1], _00356_);
  nand (_00368_, _00367_, _00366_);
  nand (_00369_, _00368_, _42882_);
  or (_00370_, \oc8051_gm_cxrom_1.cell10.data [1], _42882_);
  and (_05635_, _00370_, _00369_);
  or (_00371_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00372_, \oc8051_gm_cxrom_1.cell10.data [2], _00356_);
  nand (_00373_, _00372_, _00371_);
  nand (_00374_, _00373_, _42882_);
  or (_00375_, \oc8051_gm_cxrom_1.cell10.data [2], _42882_);
  and (_05639_, _00375_, _00374_);
  or (_00376_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00377_, \oc8051_gm_cxrom_1.cell10.data [3], _00356_);
  nand (_00378_, _00377_, _00376_);
  nand (_00379_, _00378_, _42882_);
  or (_00380_, \oc8051_gm_cxrom_1.cell10.data [3], _42882_);
  and (_05643_, _00380_, _00379_);
  or (_00381_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00382_, \oc8051_gm_cxrom_1.cell10.data [4], _00356_);
  nand (_00383_, _00382_, _00381_);
  nand (_00384_, _00383_, _42882_);
  or (_00385_, \oc8051_gm_cxrom_1.cell10.data [4], _42882_);
  and (_05647_, _00385_, _00384_);
  nor (_00386_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  nor (_00387_, \oc8051_gm_cxrom_1.cell10.data [5], _00356_);
  or (_00388_, _00387_, _00386_);
  nand (_00389_, _00388_, _42882_);
  or (_00390_, \oc8051_gm_cxrom_1.cell10.data [5], _42882_);
  and (_05651_, _00390_, _00389_);
  or (_00391_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00392_, \oc8051_gm_cxrom_1.cell10.data [6], _00356_);
  nand (_00393_, _00392_, _00391_);
  nand (_00394_, _00393_, _42882_);
  or (_00395_, \oc8051_gm_cxrom_1.cell10.data [6], _42882_);
  and (_05655_, _00395_, _00394_);
  or (_00396_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_00397_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_00398_, _00397_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_00399_, _00398_, _00396_);
  nand (_00400_, _00399_, _42882_);
  or (_00401_, \oc8051_gm_cxrom_1.cell11.data [7], _42882_);
  and (_05677_, _00401_, _00400_);
  or (_00402_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00403_, \oc8051_gm_cxrom_1.cell11.data [0], _00397_);
  nand (_00404_, _00403_, _00402_);
  nand (_00405_, _00404_, _42882_);
  or (_00406_, \oc8051_gm_cxrom_1.cell11.data [0], _42882_);
  and (_05684_, _00406_, _00405_);
  or (_00407_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00408_, \oc8051_gm_cxrom_1.cell11.data [1], _00397_);
  nand (_00409_, _00408_, _00407_);
  nand (_00410_, _00409_, _42882_);
  or (_00411_, \oc8051_gm_cxrom_1.cell11.data [1], _42882_);
  and (_05688_, _00411_, _00410_);
  or (_00412_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00413_, \oc8051_gm_cxrom_1.cell11.data [2], _00397_);
  nand (_00414_, _00413_, _00412_);
  nand (_00415_, _00414_, _42882_);
  or (_00416_, \oc8051_gm_cxrom_1.cell11.data [2], _42882_);
  and (_05692_, _00416_, _00415_);
  or (_00417_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00418_, \oc8051_gm_cxrom_1.cell11.data [3], _00397_);
  nand (_00419_, _00418_, _00417_);
  nand (_00420_, _00419_, _42882_);
  or (_00421_, \oc8051_gm_cxrom_1.cell11.data [3], _42882_);
  and (_05696_, _00421_, _00420_);
  or (_00422_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00423_, \oc8051_gm_cxrom_1.cell11.data [4], _00397_);
  nand (_00424_, _00423_, _00422_);
  nand (_00425_, _00424_, _42882_);
  or (_00426_, \oc8051_gm_cxrom_1.cell11.data [4], _42882_);
  and (_05700_, _00426_, _00425_);
  nor (_00427_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  nor (_00428_, \oc8051_gm_cxrom_1.cell11.data [5], _00397_);
  or (_00429_, _00428_, _00427_);
  nand (_00430_, _00429_, _42882_);
  or (_00431_, \oc8051_gm_cxrom_1.cell11.data [5], _42882_);
  and (_05704_, _00431_, _00430_);
  or (_00432_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00433_, \oc8051_gm_cxrom_1.cell11.data [6], _00397_);
  nand (_00434_, _00433_, _00432_);
  nand (_00435_, _00434_, _42882_);
  or (_00436_, \oc8051_gm_cxrom_1.cell11.data [6], _42882_);
  and (_05708_, _00436_, _00435_);
  or (_00437_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_00438_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_00439_, _00438_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_00440_, _00439_, _00437_);
  nand (_00441_, _00440_, _42882_);
  or (_00442_, \oc8051_gm_cxrom_1.cell12.data [7], _42882_);
  and (_05730_, _00442_, _00441_);
  or (_00443_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00444_, \oc8051_gm_cxrom_1.cell12.data [0], _00438_);
  nand (_00445_, _00444_, _00443_);
  nand (_00446_, _00445_, _42882_);
  or (_00447_, \oc8051_gm_cxrom_1.cell12.data [0], _42882_);
  and (_05737_, _00447_, _00446_);
  or (_00448_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00449_, \oc8051_gm_cxrom_1.cell12.data [1], _00438_);
  nand (_00450_, _00449_, _00448_);
  nand (_00451_, _00450_, _42882_);
  or (_00452_, \oc8051_gm_cxrom_1.cell12.data [1], _42882_);
  and (_05741_, _00452_, _00451_);
  or (_00453_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00454_, \oc8051_gm_cxrom_1.cell12.data [2], _00438_);
  nand (_00455_, _00454_, _00453_);
  nand (_00456_, _00455_, _42882_);
  or (_00457_, \oc8051_gm_cxrom_1.cell12.data [2], _42882_);
  and (_05745_, _00457_, _00456_);
  or (_00458_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00459_, \oc8051_gm_cxrom_1.cell12.data [3], _00438_);
  nand (_00460_, _00459_, _00458_);
  nand (_00461_, _00460_, _42882_);
  or (_00462_, \oc8051_gm_cxrom_1.cell12.data [3], _42882_);
  and (_05749_, _00462_, _00461_);
  or (_00463_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00464_, \oc8051_gm_cxrom_1.cell12.data [4], _00438_);
  nand (_00465_, _00464_, _00463_);
  nand (_00466_, _00465_, _42882_);
  or (_00467_, \oc8051_gm_cxrom_1.cell12.data [4], _42882_);
  and (_05753_, _00467_, _00466_);
  nor (_00468_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  nor (_00469_, \oc8051_gm_cxrom_1.cell12.data [5], _00438_);
  or (_00470_, _00469_, _00468_);
  nand (_00471_, _00470_, _42882_);
  or (_00472_, \oc8051_gm_cxrom_1.cell12.data [5], _42882_);
  and (_05757_, _00472_, _00471_);
  or (_00473_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00474_, \oc8051_gm_cxrom_1.cell12.data [6], _00438_);
  nand (_00475_, _00474_, _00473_);
  nand (_00476_, _00475_, _42882_);
  or (_00477_, \oc8051_gm_cxrom_1.cell12.data [6], _42882_);
  and (_05761_, _00477_, _00476_);
  or (_00478_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_00479_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_00480_, _00479_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_00481_, _00480_, _00478_);
  nand (_00482_, _00481_, _42882_);
  or (_00483_, \oc8051_gm_cxrom_1.cell13.data [7], _42882_);
  and (_05783_, _00483_, _00482_);
  or (_00484_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00485_, \oc8051_gm_cxrom_1.cell13.data [0], _00479_);
  nand (_00486_, _00485_, _00484_);
  nand (_00487_, _00486_, _42882_);
  or (_00488_, \oc8051_gm_cxrom_1.cell13.data [0], _42882_);
  and (_05790_, _00488_, _00487_);
  or (_00489_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00490_, \oc8051_gm_cxrom_1.cell13.data [1], _00479_);
  nand (_00491_, _00490_, _00489_);
  nand (_00492_, _00491_, _42882_);
  or (_00493_, \oc8051_gm_cxrom_1.cell13.data [1], _42882_);
  and (_05794_, _00493_, _00492_);
  or (_00494_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00495_, \oc8051_gm_cxrom_1.cell13.data [2], _00479_);
  nand (_00496_, _00495_, _00494_);
  nand (_00497_, _00496_, _42882_);
  or (_00498_, \oc8051_gm_cxrom_1.cell13.data [2], _42882_);
  and (_05798_, _00498_, _00497_);
  or (_00499_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00500_, \oc8051_gm_cxrom_1.cell13.data [3], _00479_);
  nand (_00501_, _00500_, _00499_);
  nand (_00502_, _00501_, _42882_);
  or (_00503_, \oc8051_gm_cxrom_1.cell13.data [3], _42882_);
  and (_05802_, _00503_, _00502_);
  or (_00504_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00505_, \oc8051_gm_cxrom_1.cell13.data [4], _00479_);
  nand (_00506_, _00505_, _00504_);
  nand (_00507_, _00506_, _42882_);
  or (_00508_, \oc8051_gm_cxrom_1.cell13.data [4], _42882_);
  and (_05806_, _00508_, _00507_);
  nor (_00509_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  nor (_00510_, \oc8051_gm_cxrom_1.cell13.data [5], _00479_);
  or (_00511_, _00510_, _00509_);
  nand (_00512_, _00511_, _42882_);
  or (_00513_, \oc8051_gm_cxrom_1.cell13.data [5], _42882_);
  and (_05810_, _00513_, _00512_);
  or (_00514_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00515_, \oc8051_gm_cxrom_1.cell13.data [6], _00479_);
  nand (_00516_, _00515_, _00514_);
  nand (_00517_, _00516_, _42882_);
  or (_00518_, \oc8051_gm_cxrom_1.cell13.data [6], _42882_);
  and (_05814_, _00518_, _00517_);
  or (_00519_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_00520_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_00521_, _00520_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_00522_, _00521_, _00519_);
  nand (_00523_, _00522_, _42882_);
  or (_00524_, \oc8051_gm_cxrom_1.cell14.data [7], _42882_);
  and (_05836_, _00524_, _00523_);
  or (_00525_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00526_, \oc8051_gm_cxrom_1.cell14.data [0], _00520_);
  nand (_00527_, _00526_, _00525_);
  nand (_00528_, _00527_, _42882_);
  or (_00529_, \oc8051_gm_cxrom_1.cell14.data [0], _42882_);
  and (_05843_, _00529_, _00528_);
  or (_00530_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00531_, \oc8051_gm_cxrom_1.cell14.data [1], _00520_);
  nand (_00532_, _00531_, _00530_);
  nand (_00533_, _00532_, _42882_);
  or (_00534_, \oc8051_gm_cxrom_1.cell14.data [1], _42882_);
  and (_05847_, _00534_, _00533_);
  or (_00535_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00536_, \oc8051_gm_cxrom_1.cell14.data [2], _00520_);
  nand (_00537_, _00536_, _00535_);
  nand (_00538_, _00537_, _42882_);
  or (_00539_, \oc8051_gm_cxrom_1.cell14.data [2], _42882_);
  and (_05851_, _00539_, _00538_);
  or (_00540_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00541_, \oc8051_gm_cxrom_1.cell14.data [3], _00520_);
  nand (_00542_, _00541_, _00540_);
  nand (_00544_, _00542_, _42882_);
  or (_00545_, \oc8051_gm_cxrom_1.cell14.data [3], _42882_);
  and (_05855_, _00545_, _00544_);
  or (_00547_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00549_, \oc8051_gm_cxrom_1.cell14.data [4], _00520_);
  nand (_00550_, _00549_, _00547_);
  nand (_00552_, _00550_, _42882_);
  or (_00553_, \oc8051_gm_cxrom_1.cell14.data [4], _42882_);
  and (_05859_, _00553_, _00552_);
  nor (_00555_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  nor (_00557_, \oc8051_gm_cxrom_1.cell14.data [5], _00520_);
  or (_00558_, _00557_, _00555_);
  nand (_00560_, _00558_, _42882_);
  or (_00561_, \oc8051_gm_cxrom_1.cell14.data [5], _42882_);
  and (_05863_, _00561_, _00560_);
  or (_00563_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00565_, \oc8051_gm_cxrom_1.cell14.data [6], _00520_);
  nand (_00566_, _00565_, _00563_);
  nand (_00568_, _00566_, _42882_);
  or (_00569_, \oc8051_gm_cxrom_1.cell14.data [6], _42882_);
  and (_05867_, _00569_, _00568_);
  or (_00571_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_00573_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_00574_, _00573_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_00576_, _00574_, _00571_);
  nand (_00577_, _00576_, _42882_);
  or (_00579_, \oc8051_gm_cxrom_1.cell15.data [7], _42882_);
  and (_05889_, _00579_, _00577_);
  or (_00581_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00582_, \oc8051_gm_cxrom_1.cell15.data [0], _00573_);
  nand (_00584_, _00582_, _00581_);
  nand (_00585_, _00584_, _42882_);
  or (_00587_, \oc8051_gm_cxrom_1.cell15.data [0], _42882_);
  and (_05896_, _00587_, _00585_);
  or (_00589_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00590_, \oc8051_gm_cxrom_1.cell15.data [1], _00573_);
  nand (_00592_, _00590_, _00589_);
  nand (_00593_, _00592_, _42882_);
  or (_00594_, \oc8051_gm_cxrom_1.cell15.data [1], _42882_);
  and (_05900_, _00594_, _00593_);
  or (_00595_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00596_, \oc8051_gm_cxrom_1.cell15.data [2], _00573_);
  nand (_00597_, _00596_, _00595_);
  nand (_00598_, _00597_, _42882_);
  or (_00599_, \oc8051_gm_cxrom_1.cell15.data [2], _42882_);
  and (_05904_, _00599_, _00598_);
  or (_00600_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00601_, \oc8051_gm_cxrom_1.cell15.data [3], _00573_);
  nand (_00602_, _00601_, _00600_);
  nand (_00603_, _00602_, _42882_);
  or (_00604_, \oc8051_gm_cxrom_1.cell15.data [3], _42882_);
  and (_05908_, _00604_, _00603_);
  or (_00605_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00606_, \oc8051_gm_cxrom_1.cell15.data [4], _00573_);
  nand (_00607_, _00606_, _00605_);
  nand (_00608_, _00607_, _42882_);
  or (_00609_, \oc8051_gm_cxrom_1.cell15.data [4], _42882_);
  and (_05912_, _00609_, _00608_);
  nor (_00610_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  nor (_00611_, \oc8051_gm_cxrom_1.cell15.data [5], _00573_);
  or (_00612_, _00611_, _00610_);
  nand (_00613_, _00612_, _42882_);
  or (_00614_, \oc8051_gm_cxrom_1.cell15.data [5], _42882_);
  and (_05916_, _00614_, _00613_);
  or (_00615_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00616_, \oc8051_gm_cxrom_1.cell15.data [6], _00573_);
  nand (_00617_, _00616_, _00615_);
  nand (_00618_, _00617_, _42882_);
  or (_00619_, \oc8051_gm_cxrom_1.cell15.data [6], _42882_);
  and (_05920_, _00619_, _00618_);
  nor (_09695_, _38255_, rst);
  and (_00620_, _38246_, _38280_);
  and (_00621_, _00620_, _36920_);
  not (_00622_, _00621_);
  and (_00623_, _38218_, _38226_);
  and (_00624_, _38281_, _38217_);
  nor (_00625_, _00624_, _00623_);
  and (_00626_, _00625_, _00622_);
  and (_00627_, _38280_, _36909_);
  or (_00628_, _38246_, _38217_);
  nand (_00629_, _00628_, _00627_);
  and (_00630_, _00629_, _00626_);
  and (_00631_, _36450_, _42882_);
  not (_00632_, _00631_);
  or (_00633_, _00632_, _00623_);
  or (_09698_, _00633_, _00630_);
  not (_00634_, _37117_);
  and (_00635_, _37357_, _00634_);
  and (_00636_, _00635_, _37630_);
  not (_00637_, _37905_);
  and (_00638_, _38210_, _38145_);
  and (_00639_, _00638_, _38185_);
  and (_00640_, _00639_, _00637_);
  and (_00641_, _00640_, _00636_);
  not (_00642_, _36844_);
  nor (_00643_, _38210_, _00642_);
  nor (_00644_, _37357_, _37117_);
  and (_00645_, _00644_, _37630_);
  and (_00646_, _00645_, _00643_);
  not (_00647_, _38185_);
  not (_00648_, _38145_);
  and (_00649_, _38210_, _00648_);
  and (_00650_, _00649_, _00647_);
  nor (_00651_, _37630_, _00642_);
  and (_00652_, _00651_, _00635_);
  and (_00653_, _00652_, _00650_);
  or (_00654_, _00653_, _00646_);
  or (_00655_, _00654_, _00641_);
  not (_00656_, _37357_);
  and (_00657_, _00656_, _37117_);
  and (_00658_, _00657_, _00651_);
  and (_00659_, _00658_, _00640_);
  and (_00660_, _00639_, _37905_);
  and (_00661_, _37357_, _37117_);
  and (_00662_, _00661_, _37630_);
  and (_00663_, _00662_, _00660_);
  or (_00664_, _00663_, _00659_);
  or (_00665_, _00664_, _00655_);
  and (_00666_, _37905_, _00647_);
  and (_00667_, _00666_, _00638_);
  and (_00668_, _00667_, _00661_);
  and (_00669_, _37630_, _00642_);
  nor (_00670_, _00669_, _00651_);
  and (_00671_, _00670_, _00668_);
  and (_00672_, _00667_, _36844_);
  and (_00673_, _00672_, _00657_);
  or (_00674_, _00673_, _00671_);
  or (_00675_, _00674_, _00665_);
  and (_00676_, _00638_, _00647_);
  not (_00677_, _00676_);
  nor (_00678_, _37630_, _36844_);
  and (_00679_, _00678_, _00657_);
  nor (_00680_, _00679_, _00637_);
  nor (_00681_, _00680_, _00677_);
  not (_00682_, _00681_);
  and (_00683_, _00669_, _00657_);
  and (_00684_, _00683_, _00667_);
  and (_00685_, _00661_, _00651_);
  and (_00686_, _00685_, _00667_);
  nor (_00687_, _00686_, _00684_);
  and (_00688_, _00687_, _00682_);
  not (_00689_, _37630_);
  and (_00690_, _00644_, _00689_);
  and (_00691_, _00690_, _00639_);
  and (_00692_, _00635_, _00689_);
  and (_00693_, _38185_, _36844_);
  and (_00694_, _00693_, _00649_);
  and (_00695_, _00694_, _00692_);
  nor (_00696_, _37630_, _00656_);
  and (_00697_, _00696_, _00643_);
  and (_00698_, _00697_, _00634_);
  or (_00699_, _00698_, _00695_);
  and (_00700_, _00690_, _00667_);
  or (_00701_, _00700_, _00699_);
  or (_00702_, _00701_, _00691_);
  and (_00703_, _00666_, _00649_);
  and (_00704_, _00703_, _00642_);
  and (_00705_, _00704_, _00635_);
  and (_00706_, _37630_, _36844_);
  and (_00707_, _00706_, _00644_);
  and (_00708_, _00650_, _00637_);
  and (_00709_, _00708_, _00707_);
  or (_00710_, _00709_, _00705_);
  and (_00711_, _00669_, _00635_);
  and (_00712_, _00711_, _00667_);
  and (_00713_, _00661_, _00689_);
  and (_00714_, _00713_, _00660_);
  or (_00715_, _00714_, _00712_);
  or (_00716_, _00715_, _00710_);
  nor (_00717_, _00716_, _00702_);
  nand (_00718_, _00717_, _00688_);
  or (_00719_, _00718_, _00675_);
  and (_00720_, _00719_, _36461_);
  not (_00721_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_00722_, _36439_, _18199_);
  and (_00723_, _00722_, _38241_);
  nor (_00724_, _00723_, _00721_);
  or (_00725_, _00724_, rst);
  or (_09701_, _00725_, _00720_);
  nand (_00726_, _37117_, _36385_);
  or (_00727_, _36385_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_00728_, _00727_, _42882_);
  and (_09704_, _00728_, _00726_);
  and (_00729_, \oc8051_top_1.oc8051_sfr1.wait_data , _42882_);
  and (_00730_, _00729_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00731_, _38246_, _38232_);
  or (_00732_, _00731_, _38247_);
  or (_00733_, _00732_, _38316_);
  and (_00734_, _38218_, _38289_);
  or (_00735_, _00734_, _38266_);
  or (_00736_, _00735_, _00733_);
  and (_00737_, _38235_, _38281_);
  and (_00738_, _00623_, _36920_);
  nor (_00739_, _00738_, _00737_);
  nand (_00740_, _00739_, _38341_);
  or (_00741_, _00740_, _00736_);
  and (_00742_, _00741_, _00631_);
  or (_09707_, _00742_, _00730_);
  and (_00743_, _38233_, _38191_);
  and (_00744_, _00743_, _38289_);
  and (_00745_, _38215_, _36920_);
  and (_00746_, _00745_, _38264_);
  or (_00747_, _00746_, _38360_);
  and (_00748_, _38246_, _38227_);
  or (_00749_, _00748_, _38219_);
  or (_00750_, _00749_, _00747_);
  or (_00751_, _00750_, _00744_);
  and (_00752_, _00751_, _36450_);
  and (_00753_, _38350_, _00721_);
  not (_00754_, _38238_);
  and (_00755_, _00754_, _00753_);
  and (_00756_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00757_, _00756_, _00755_);
  or (_00758_, _00757_, _00752_);
  and (_09710_, _00758_, _42882_);
  and (_00759_, _00729_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_00760_, _38235_, _38299_);
  or (_00761_, _38299_, _38265_);
  and (_00762_, _00761_, _38275_);
  or (_00763_, _00762_, _00760_);
  and (_00764_, _00743_, _38307_);
  or (_00765_, _00764_, _00763_);
  and (_00766_, _00761_, _38215_);
  and (_00767_, _38215_, _36909_);
  and (_00768_, _00767_, _38298_);
  or (_00769_, _00768_, _00766_);
  or (_00770_, _00769_, _38368_);
  and (_00771_, _38235_, _38283_);
  and (_00772_, _38317_, _38215_);
  or (_00773_, _00772_, _00771_);
  or (_00774_, _00773_, _00749_);
  or (_00775_, _00774_, _00770_);
  or (_00776_, _00775_, _00765_);
  and (_00777_, _00776_, _00631_);
  or (_09713_, _00777_, _00759_);
  and (_00778_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00779_, _38276_, _36450_);
  or (_00780_, _00779_, _00778_);
  or (_00781_, _00780_, _00755_);
  and (_09716_, _00781_, _42882_);
  and (_00782_, _38307_, _38260_);
  and (_00783_, _38274_, _38245_);
  and (_00784_, _00783_, _36909_);
  or (_00785_, _00784_, _00782_);
  and (_00786_, _00785_, _38243_);
  or (_00787_, _00786_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00788_, _00785_, _00738_);
  and (_00789_, _00788_, _36396_);
  and (_00790_, _38280_, _38192_);
  and (_00791_, _00790_, _38270_);
  and (_00792_, _38226_, _38375_);
  and (_00793_, _38246_, _38281_);
  or (_00794_, _00793_, _00792_);
  or (_00795_, _00794_, _00791_);
  and (_00796_, _00795_, _00753_);
  or (_00797_, _00796_, _00789_);
  or (_00798_, _00797_, _00787_);
  or (_00799_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18199_);
  and (_00800_, _00799_, _42882_);
  and (_09719_, _00800_, _00798_);
  and (_00801_, _00729_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_00802_, _00746_, _38290_);
  or (_00803_, _38307_, _38289_);
  and (_00804_, _00803_, _38359_);
  or (_00805_, _00804_, _38266_);
  or (_00806_, _00805_, _00802_);
  and (_00807_, _38235_, _38307_);
  or (_00808_, _00807_, _38308_);
  and (_00809_, _00767_, _38264_);
  or (_00810_, _00768_, _00809_);
  or (_00811_, _38376_, _38306_);
  or (_00812_, _00811_, _00810_);
  or (_00813_, _00812_, _00808_);
  or (_00814_, _38318_, _38261_);
  or (_00815_, _00814_, _00813_);
  or (_00816_, _00815_, _00806_);
  and (_00817_, _00816_, _00631_);
  or (_09722_, _00817_, _00801_);
  and (_00818_, _00729_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_00819_, _00743_, _38287_);
  and (_00820_, _38218_, _38294_);
  or (_00821_, _00820_, _00744_);
  or (_00822_, _00821_, _00819_);
  or (_00823_, _00822_, _00769_);
  not (_00824_, _38322_);
  and (_00825_, _38235_, _38312_);
  or (_00826_, _00825_, _00824_);
  and (_00827_, _38271_, _38263_);
  or (_00828_, _00827_, _38386_);
  and (_00829_, _38359_, _38265_);
  or (_00830_, _00829_, _00828_);
  or (_00831_, _00830_, _00826_);
  or (_00832_, _00831_, _00823_);
  and (_00833_, _00745_, _38263_);
  and (_00834_, _00745_, _38222_);
  or (_00835_, _00834_, _00833_);
  nor (_00836_, _38366_, _38343_);
  nand (_00837_, _00836_, _38314_);
  or (_00838_, _00837_, _00835_);
  or (_00839_, _00838_, _00765_);
  or (_00840_, _00839_, _00832_);
  and (_00841_, _00840_, _00631_);
  or (_09725_, _00841_, _00818_);
  and (_00842_, _00743_, _38295_);
  or (_00843_, _00842_, _38363_);
  and (_00844_, _00767_, _38225_);
  and (_00845_, _00844_, _37171_);
  or (_00846_, _00845_, _38370_);
  and (_00847_, _38295_, _38215_);
  or (_00848_, _00847_, _00846_);
  or (_00849_, _00848_, _00843_);
  and (_00850_, _00743_, _38227_);
  or (_00851_, _00850_, _00849_);
  and (_00852_, _00851_, _36450_);
  nand (_00853_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_00854_, _00853_, _38251_);
  or (_00855_, _00854_, _00852_);
  and (_09728_, _00855_, _42882_);
  nand (_00856_, _38344_, _38319_);
  or (_00857_, _00856_, _00762_);
  or (_00858_, _38290_, _38267_);
  and (_00859_, _38221_, _36909_);
  and (_00860_, _00859_, _38275_);
  or (_00861_, _00860_, _38308_);
  or (_00862_, _00861_, _00782_);
  or (_00863_, _38321_, _38278_);
  or (_00864_, _00863_, _00862_);
  or (_00865_, _00864_, _00858_);
  or (_00866_, _00865_, _00857_);
  and (_00867_, _00745_, _38226_);
  or (_00868_, _00867_, _38292_);
  or (_00869_, _00868_, _00784_);
  and (_00870_, _00767_, _38221_);
  or (_00871_, _00870_, _38381_);
  or (_00872_, _00871_, _38327_);
  or (_00873_, _00872_, _00869_);
  and (_00874_, _38359_, _37707_);
  and (_00875_, _38362_, _38221_);
  or (_00876_, _00875_, _38366_);
  or (_00877_, _00876_, _00874_);
  or (_00878_, _00877_, _00747_);
  or (_00879_, _00878_, _00873_);
  or (_00880_, _00879_, _00769_);
  or (_00881_, _00880_, _00866_);
  and (_00882_, _00881_, _36450_);
  and (_00883_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00884_, _00786_, _00755_);
  and (_00885_, _38243_, _38339_);
  or (_00886_, _00885_, _00884_);
  or (_00887_, _00886_, _00883_);
  or (_00888_, _00887_, _00882_);
  and (_09731_, _00888_, _42882_);
  nor (_09790_, _38396_, rst);
  nor (_09792_, _38355_, rst);
  or (_09795_, _00632_, _00626_);
  nor (_00889_, _00623_, _00620_);
  or (_09798_, _00889_, _00632_);
  or (_00890_, _00714_, _00705_);
  or (_00891_, _00641_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_00892_, _00891_, _00890_);
  and (_00893_, _00892_, _00723_);
  nor (_00894_, _00722_, _38241_);
  or (_00895_, _00894_, rst);
  or (_09801_, _00895_, _00893_);
  nand (_00896_, _37905_, _36385_);
  or (_00897_, _36385_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_00898_, _00897_, _42882_);
  and (_09804_, _00898_, _00896_);
  not (_00899_, _36385_);
  or (_00900_, _38185_, _00899_);
  or (_00901_, _36385_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_00902_, _00901_, _42882_);
  and (_09807_, _00902_, _00900_);
  nand (_00903_, _38145_, _36385_);
  or (_00904_, _36385_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_00905_, _00904_, _42882_);
  and (_09810_, _00905_, _00903_);
  nand (_00906_, _38210_, _36385_);
  or (_00907_, _36385_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_00908_, _00907_, _42882_);
  and (_09813_, _00908_, _00906_);
  or (_00909_, _36844_, _00899_);
  or (_00910_, _36385_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_00911_, _00910_, _42882_);
  and (_09816_, _00911_, _00909_);
  nand (_00912_, _37630_, _36385_);
  or (_00913_, _36385_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_00914_, _00913_, _42882_);
  and (_09819_, _00914_, _00912_);
  nand (_00915_, _37357_, _36385_);
  or (_00916_, _36385_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_00917_, _00916_, _42882_);
  and (_09822_, _00917_, _00915_);
  and (_00918_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00919_, _00918_, _00796_);
  and (_00920_, _00919_, _42882_);
  and (_00921_, _38311_, _38215_);
  and (_00922_, _00921_, _36909_);
  or (_00923_, _00922_, _00847_);
  and (_00924_, _00743_, _38312_);
  or (_00926_, _00924_, _00748_);
  or (_00927_, _00926_, _00923_);
  or (_00928_, _38295_, _38281_);
  and (_00929_, _00928_, _00743_);
  or (_00930_, _38298_, _38265_);
  and (_00931_, _00930_, _38235_);
  or (_00932_, _00931_, _00929_);
  or (_00933_, _00932_, _00927_);
  and (_00934_, _00743_, _38326_);
  or (_00935_, _38311_, _38280_);
  and (_00936_, _00935_, _00745_);
  or (_00937_, _00936_, _00934_);
  and (_00938_, _38235_, _38223_);
  and (_00939_, _00627_, _38235_);
  or (_00940_, _00939_, _00938_);
  or (_00941_, _00940_, _00937_);
  or (_00942_, _00834_, _00819_);
  or (_00943_, _00846_, _38369_);
  or (_00944_, _00943_, _00942_);
  and (_00945_, _38227_, _38359_);
  or (_00946_, _00945_, _38219_);
  or (_00947_, _00850_, _00820_);
  or (_00948_, _00947_, _00946_);
  and (_00949_, _00935_, _38271_);
  and (_00950_, _38287_, _38359_);
  or (_00951_, _00950_, _00949_);
  or (_00952_, _00951_, _00948_);
  or (_00953_, _00952_, _00944_);
  or (_00954_, _00953_, _00941_);
  or (_00955_, _00954_, _00933_);
  and (_00957_, _00955_, _00631_);
  or (_09825_, _00957_, _00920_);
  and (_00958_, _00729_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_00959_, _00926_, _00835_);
  or (_00960_, _38312_, _38287_);
  and (_00961_, _00960_, _38260_);
  and (_00962_, _38235_, _38331_);
  or (_00963_, _00962_, _00961_);
  or (_00964_, _00963_, _00959_);
  and (_00965_, _38235_, _38287_);
  and (_00966_, _37685_, _37421_);
  and (_00967_, _00767_, _00966_);
  and (_00968_, _00967_, _37171_);
  nor (_00969_, _00968_, _38365_);
  not (_00970_, _00969_);
  or (_00971_, _00970_, _00771_);
  or (_00972_, _00971_, _00965_);
  nand (_00973_, _00739_, _38291_);
  or (_00974_, _00973_, _00972_);
  or (_00975_, _00974_, _00830_);
  or (_00977_, _00975_, _00964_);
  and (_00978_, _00977_, _00631_);
  or (_34273_, _00978_, _00958_);
  or (_00979_, _00784_, _38327_);
  or (_00980_, _00867_, _38381_);
  or (_00981_, _00980_, _00866_);
  or (_00982_, _00981_, _00979_);
  and (_00983_, _00982_, _36450_);
  and (_00984_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00985_, _00984_, _00886_);
  or (_00986_, _00985_, _00983_);
  and (_34275_, _00986_, _42882_);
  and (_00987_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00988_, _00987_, _00884_);
  and (_00989_, _00988_, _42882_);
  and (_00990_, _38342_, _36920_);
  or (_00991_, _00990_, _00785_);
  or (_00992_, _00991_, _00877_);
  or (_00993_, _00992_, _38360_);
  and (_00994_, _00993_, _00631_);
  or (_34278_, _00994_, _00989_);
  and (_00995_, _00842_, _36909_);
  or (_00996_, _00623_, _38237_);
  or (_00997_, _00996_, _00934_);
  or (_00998_, _00997_, _00995_);
  or (_00999_, _00938_, _00825_);
  and (_01000_, _00627_, _38275_);
  or (_01001_, _01000_, _00965_);
  or (_01002_, _01001_, _00999_);
  or (_01003_, _01002_, _00998_);
  or (_01004_, _00923_, _00820_);
  or (_01005_, _01004_, _00943_);
  or (_01006_, _01005_, _01003_);
  and (_01007_, _00743_, _38317_);
  or (_01008_, _01007_, _00850_);
  or (_01009_, _01008_, _00737_);
  or (_01010_, _01009_, _00939_);
  and (_01011_, _38235_, _38289_);
  or (_01012_, _01011_, _38236_);
  or (_01013_, _01012_, _00931_);
  or (_01014_, _01013_, _01010_);
  and (_01015_, _00859_, _38359_);
  or (_01016_, _00870_, _00945_);
  or (_01017_, _01016_, _01015_);
  or (_01018_, _01017_, _00785_);
  and (_01019_, _38327_, _38262_);
  and (_01020_, _00842_, _36920_);
  or (_01021_, _01020_, _38224_);
  or (_01022_, _01021_, _01019_);
  or (_01023_, _01022_, _01018_);
  or (_01024_, _01023_, _01014_);
  or (_01025_, _01024_, _01006_);
  and (_01026_, _01025_, _36450_);
  and (_01027_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_01028_, _38238_, _36396_);
  or (_01029_, _00796_, _01028_);
  or (_01030_, _01029_, _01027_);
  or (_01031_, _01030_, _01026_);
  and (_34280_, _01031_, _42882_);
  and (_01032_, _00627_, _38359_);
  or (_01033_, _38237_, _00945_);
  or (_01034_, _01033_, _38327_);
  or (_01035_, _01034_, _01032_);
  or (_01036_, _01035_, _01004_);
  or (_01037_, _01036_, _00943_);
  and (_01038_, _00767_, _38280_);
  or (_01039_, _00860_, _00748_);
  or (_01040_, _01039_, _01038_);
  or (_01041_, _01040_, _38230_);
  and (_01042_, _00960_, _38218_);
  or (_01043_, _01042_, _38332_);
  or (_01044_, _01043_, _01041_);
  or (_01045_, _01044_, _01014_);
  or (_01046_, _01045_, _01037_);
  and (_01047_, _01046_, _36450_);
  and (_01048_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01049_, _01048_, _01029_);
  or (_01050_, _01049_, _01047_);
  and (_34282_, _01050_, _42882_);
  and (_01051_, _00729_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_01052_, _00850_, _42307_);
  or (_01053_, _01052_, _00804_);
  or (_01054_, _38307_, _38265_);
  and (_01055_, _01054_, _38218_);
  and (_01056_, _38235_, _38265_);
  or (_01057_, _01056_, _00764_);
  or (_01058_, _01057_, _01055_);
  or (_01059_, _01058_, _01053_);
  or (_01060_, _00945_, _38273_);
  or (_01061_, _01060_, _00995_);
  or (_01062_, _00845_, _00746_);
  and (_01063_, _38317_, _38217_);
  and (_01064_, _01063_, _37960_);
  or (_01065_, _01064_, _01062_);
  or (_01066_, _01065_, _01061_);
  and (_01067_, _38218_, _38334_);
  and (_01068_, _38362_, _38295_);
  and (_01069_, _38334_, _38215_);
  or (_01070_, _01069_, _01068_);
  nor (_01071_, _01070_, _01067_);
  nand (_01072_, _01071_, _42311_);
  or (_01073_, _01072_, _01066_);
  or (_01074_, _00858_, _00812_);
  or (_01075_, _01074_, _01073_);
  or (_01076_, _01075_, _01059_);
  and (_01077_, _01076_, _00631_);
  or (_34284_, _01077_, _01051_);
  or (_01078_, _00923_, _38329_);
  or (_01079_, _01067_, _01056_);
  or (_01080_, _01079_, _01021_);
  or (_01081_, _01080_, _01078_);
  or (_01082_, _00744_, _38313_);
  or (_01083_, _00829_, _00827_);
  or (_01084_, _01083_, _01082_);
  and (_01085_, _38218_, _38307_);
  or (_01086_, _00833_, _38219_);
  or (_01087_, _01086_, _01085_);
  or (_01088_, _01087_, _38371_);
  or (_01089_, _01088_, _01084_);
  or (_01090_, _00998_, _00826_);
  or (_01091_, _01090_, _01089_);
  or (_01092_, _01091_, _01081_);
  and (_01093_, _01092_, _00631_);
  and (_01094_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_01095_, _38237_, _36407_);
  or (_01096_, _01095_, _01094_);
  and (_01097_, _01096_, _42882_);
  or (_34286_, _01097_, _01093_);
  and (_01098_, _38326_, _38359_);
  or (_01099_, _01098_, _00744_);
  or (_01100_, _01062_, _00922_);
  or (_01101_, _01100_, _01099_);
  and (_01102_, _38218_, _38295_);
  or (_01103_, _00772_, _01063_);
  or (_01104_, _01103_, _01102_);
  not (_01105_, _38364_);
  or (_01106_, _01105_, _42310_);
  or (_01107_, _01106_, _01104_);
  or (_01108_, _01107_, _01101_);
  not (_01109_, _00934_);
  and (_01110_, _01109_, _38328_);
  not (_01111_, _01110_);
  or (_01112_, _01111_, _01010_);
  or (_01113_, _01112_, _01108_);
  or (_01114_, _00770_, _00765_);
  or (_01115_, _01114_, _01113_);
  and (_01116_, _01115_, _36450_);
  and (_01117_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01118_, _01117_, _38249_);
  or (_01119_, _01118_, _01116_);
  and (_34288_, _01119_, _42882_);
  and (_01120_, _38218_, _38298_);
  or (_01121_, _01120_, _01063_);
  or (_01122_, _01121_, _38327_);
  or (_01123_, _01098_, _42307_);
  or (_01124_, _01123_, _01122_);
  or (_01125_, _01057_, _00802_);
  or (_01126_, _01125_, _01124_);
  or (_01127_, _00939_, _00934_);
  or (_01128_, _38360_, _38366_);
  or (_01129_, _01128_, _00922_);
  or (_01130_, _01129_, _01127_);
  or (_01131_, _01130_, _00769_);
  or (_01132_, _01131_, _00763_);
  or (_01133_, _01132_, _01126_);
  and (_01134_, _01133_, _36450_);
  and (_01135_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01136_, _01135_, _38250_);
  or (_01137_, _01136_, _01134_);
  and (_34290_, _01137_, _42882_);
  and (_01138_, _00729_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_01139_, _42311_);
  or (_01140_, _01052_, _01139_);
  or (_01141_, _01079_, _01055_);
  or (_01142_, _01141_, _01140_);
  not (_01143_, _38245_);
  or (_01144_, _38218_, _01143_);
  and (_01145_, _01144_, _38317_);
  or (_01146_, _00734_, _38261_);
  or (_01147_, _01146_, _01145_);
  or (_01148_, _01147_, _00849_);
  or (_01149_, _01148_, _01142_);
  and (_01150_, _01149_, _00631_);
  or (_34292_, _01150_, _01138_);
  nor (_38955_, _37117_, rst);
  nor (_38956_, _42266_, rst);
  and (_01151_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_01152_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_01153_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_01154_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_01155_, _01154_, _01153_);
  and (_01156_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01157_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_01158_, _01157_, _01156_);
  and (_01159_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_01160_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_01161_, _01160_, _01159_);
  and (_01162_, _01161_, _01158_);
  and (_01163_, _01162_, _01155_);
  nor (_01164_, _01163_, _36636_);
  nor (_01165_, _01164_, _01152_);
  nor (_01166_, _01165_, _42250_);
  nor (_01167_, _01166_, _01151_);
  nor (_38958_, _01167_, rst);
  nor (_38968_, _37905_, rst);
  and (_38969_, _38185_, _42882_);
  nor (_38970_, _38145_, rst);
  nor (_38971_, _38210_, rst);
  and (_38972_, _36844_, _42882_);
  nor (_38973_, _37630_, rst);
  nor (_38974_, _37357_, rst);
  nor (_38975_, _42464_, rst);
  nor (_38976_, _42384_, rst);
  nor (_38978_, _42589_, rst);
  nor (_38979_, _42429_, rst);
  nor (_38980_, _42336_, rst);
  nor (_38981_, _42551_, rst);
  nor (_38982_, _42523_, rst);
  and (_01168_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_01169_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_01170_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_01171_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_01172_, _01171_, _01170_);
  and (_01173_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_01174_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_01175_, _01174_, _01173_);
  and (_01176_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_01177_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_01178_, _01177_, _01176_);
  and (_01179_, _01178_, _01175_);
  and (_01180_, _01179_, _01172_);
  nor (_01181_, _01180_, _36636_);
  nor (_01182_, _01181_, _01169_);
  nor (_01183_, _01182_, _42250_);
  nor (_01184_, _01183_, _01168_);
  nor (_38984_, _01184_, rst);
  and (_01185_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_01186_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_01187_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_01188_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_01189_, _01188_, _01187_);
  and (_01190_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_01191_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_01192_, _01191_, _01190_);
  and (_01193_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_01194_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_01195_, _01194_, _01193_);
  and (_01196_, _01195_, _01192_);
  and (_01197_, _01196_, _01189_);
  nor (_01198_, _01197_, _36636_);
  nor (_01199_, _01198_, _01186_);
  nor (_01200_, _01199_, _42250_);
  nor (_01201_, _01200_, _01185_);
  nor (_38985_, _01201_, rst);
  and (_01202_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_01203_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_01204_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_01205_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01206_, _01205_, _01204_);
  and (_01207_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_01208_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_01209_, _01208_, _01207_);
  and (_01211_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_01213_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_01215_, _01213_, _01211_);
  and (_01217_, _01215_, _01209_);
  and (_01219_, _01217_, _01206_);
  nor (_01221_, _01219_, _36636_);
  nor (_01223_, _01221_, _01203_);
  nor (_01225_, _01223_, _42250_);
  nor (_01227_, _01225_, _01202_);
  nor (_38986_, _01227_, rst);
  and (_01230_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_01232_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_01234_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_01236_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_01238_, _01236_, _01234_);
  and (_01240_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_01242_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_01244_, _01242_, _01240_);
  and (_01246_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_01248_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_01250_, _01248_, _01246_);
  and (_01252_, _01250_, _01244_);
  and (_01254_, _01252_, _01238_);
  nor (_01256_, _01254_, _36636_);
  nor (_01258_, _01256_, _01232_);
  nor (_01260_, _01258_, _42250_);
  nor (_01262_, _01260_, _01230_);
  nor (_38987_, _01262_, rst);
  and (_01265_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_01267_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_01269_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_01271_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_01273_, _01271_, _01269_);
  and (_01275_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_01277_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_01279_, _01277_, _01275_);
  and (_01281_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_01283_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_01285_, _01283_, _01281_);
  and (_01287_, _01285_, _01279_);
  and (_01289_, _01287_, _01273_);
  nor (_01291_, _01289_, _36636_);
  nor (_01293_, _01291_, _01267_);
  nor (_01295_, _01293_, _42250_);
  nor (_01297_, _01295_, _01265_);
  nor (_38988_, _01297_, rst);
  and (_01300_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_01302_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_01304_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_01305_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_01306_, _01305_, _01304_);
  and (_01307_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_01308_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_01309_, _01308_, _01307_);
  and (_01310_, _01309_, _01306_);
  and (_01311_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_01312_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_01313_, _01312_, _01311_);
  and (_01314_, _01313_, _01310_);
  nor (_01315_, _01314_, _36636_);
  nor (_01316_, _01315_, _01302_);
  nor (_01317_, _01316_, _42250_);
  nor (_01318_, _01317_, _01300_);
  nor (_38990_, _01318_, rst);
  and (_01319_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_01320_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_01321_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_01322_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_01323_, _01322_, _01321_);
  and (_01324_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_01325_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_01326_, _01325_, _01324_);
  and (_01327_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_01328_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_01329_, _01328_, _01327_);
  and (_01330_, _01329_, _01326_);
  and (_01331_, _01330_, _01323_);
  nor (_01332_, _01331_, _36636_);
  nor (_01333_, _01332_, _01320_);
  nor (_01334_, _01333_, _42250_);
  nor (_01335_, _01334_, _01319_);
  nor (_38991_, _01335_, rst);
  and (_01336_, _36461_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_01337_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_01338_, _01336_, _38536_);
  and (_01339_, _01338_, _42882_);
  and (_39015_, _01339_, _01337_);
  not (_01340_, _01336_);
  or (_01341_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_01342_, _36461_, _42882_);
  and (_00000_, _01342_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_01343_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _42882_);
  or (_01344_, _01343_, _00000_);
  and (_39016_, _01344_, _01341_);
  nor (_39054_, _42304_, rst);
  nor (_39056_, _42342_, rst);
  and (_39057_, _42300_, _42882_);
  not (_01345_, _38352_);
  nor (_01346_, _38341_, _38350_);
  nor (_01347_, _42448_, _27703_);
  and (_01348_, _42448_, _27703_);
  nor (_01349_, _01348_, _01347_);
  nor (_01350_, _42365_, _27845_);
  and (_01351_, _42365_, _27845_);
  nor (_01352_, _01351_, _01350_);
  nor (_01353_, _01352_, _01349_);
  nor (_01354_, _42573_, _27374_);
  and (_01355_, _42573_, _27374_);
  nor (_01356_, _01355_, _01354_);
  nor (_01357_, _42527_, _27242_);
  and (_01358_, _42527_, _27242_);
  nor (_01359_, _01358_, _01357_);
  nor (_01360_, _01359_, _01356_);
  and (_01361_, _01360_, _01353_);
  and (_01362_, _01361_, _42639_);
  nor (_01363_, _31304_, _39838_);
  and (_01364_, _01363_, _01362_);
  and (_01365_, _01364_, _01346_);
  not (_01366_, _01365_);
  nor (_01367_, _42402_, _26902_);
  and (_01368_, _42402_, _26902_);
  nor (_01369_, _01368_, _01367_);
  and (_01370_, _42484_, _32545_);
  nor (_01371_, _01370_, _01369_);
  nor (_01372_, _42610_, _26781_);
  and (_01373_, _42610_, _26781_);
  nor (_01374_, _01373_, _01372_);
  nor (_01375_, _42484_, _32545_);
  or (_01376_, _01375_, _39217_);
  nor (_01377_, _01376_, _01374_);
  and (_01378_, _01377_, _01362_);
  and (_01379_, _01378_, _01371_);
  nor (_01380_, _27549_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_01381_, _01380_, _01379_);
  not (_01382_, _01381_);
  and (_01383_, _38298_, _38260_);
  nor (_01384_, _01383_, _00783_);
  nor (_01385_, _01384_, _36407_);
  not (_01386_, _38296_);
  and (_01387_, _38223_, _38375_);
  nor (_01388_, _01387_, _00731_);
  nor (_01389_, _01346_, _38248_);
  not (_01390_, _31455_);
  nand (_01391_, _33513_, _01390_);
  or (_01392_, _01391_, _29030_);
  nor (_01393_, _01392_, _34232_);
  and (_01394_, _01393_, _34960_);
  and (_01395_, _01394_, _28569_);
  and (_01396_, _01395_, _01389_);
  and (_01397_, _01396_, _35744_);
  and (_01398_, _01397_, _29216_);
  not (_01399_, _01398_);
  and (_01400_, _01346_, _28931_);
  not (_01401_, _01400_);
  not (_01402_, _38248_);
  nor (_01403_, _01346_, _38297_);
  nor (_01404_, _01403_, _01402_);
  and (_01405_, _01404_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_01406_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_01407_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01408_, _01407_, _01406_);
  nor (_01409_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_01410_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01411_, _01410_, _01409_);
  and (_01412_, _01411_, _01408_);
  and (_01413_, _01412_, _38394_);
  nor (_01414_, _01413_, _01405_);
  and (_01415_, _01414_, _01401_);
  and (_01416_, _01415_, _01399_);
  or (_01417_, _38334_, _38223_);
  or (_01418_, _01417_, _38326_);
  and (_01419_, _01418_, _38246_);
  not (_01420_, _01419_);
  not (_01421_, _00809_);
  nor (_01422_, _01007_, _38306_);
  and (_01423_, _01422_, _01421_);
  and (_01424_, _01423_, _00969_);
  and (_01425_, _01424_, _01420_);
  not (_01426_, _01425_);
  and (_01427_, _01426_, _01416_);
  and (_01428_, _38247_, _36920_);
  not (_01429_, _01428_);
  and (_01430_, _01429_, _38340_);
  nor (_01431_, _01430_, _01416_);
  nor (_01432_, _01431_, _01427_);
  and (_01433_, _01432_, _01388_);
  and (_01434_, _01433_, _01386_);
  nor (_01435_, _38352_, _38243_);
  nor (_01436_, _01435_, _01434_);
  nor (_01437_, _01436_, _01385_);
  not (_01438_, _38875_);
  nor (_01439_, _38901_, _01438_);
  and (_01440_, _01439_, _38883_);
  not (_01441_, _01440_);
  and (_01442_, _01441_, _01404_);
  not (_01443_, _39133_);
  and (_01444_, _01443_, _38394_);
  nor (_01445_, _01444_, _01442_);
  not (_01446_, _01445_);
  nor (_01447_, _01446_, _01437_);
  and (_01448_, _01447_, _01382_);
  and (_01449_, _01448_, _01366_);
  and (_01450_, _01449_, _01345_);
  and (_39061_, _01450_, _42882_);
  and (_39062_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _42882_);
  and (_39063_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _42882_);
  and (_01451_, _00969_, _38341_);
  and (_01452_, _01451_, _01422_);
  nor (_01453_, _01452_, _42317_);
  and (_01454_, _01383_, _36396_);
  not (_01455_, _01454_);
  and (_01456_, _38246_, _38295_);
  and (_01457_, _01456_, _36396_);
  nor (_01458_, _01457_, _38352_);
  and (_01459_, _01458_, _01455_);
  not (_01460_, _01459_);
  nor (_01461_, _01460_, _01453_);
  and (_01462_, _01461_, _42266_);
  not (_01463_, _01167_);
  nor (_01464_, _01461_, _01463_);
  nor (_01465_, _01464_, _01462_);
  and (_01466_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01467_, _01466_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01468_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_01469_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01470_, _01461_, _42523_);
  not (_01471_, _01335_);
  nor (_01472_, _01461_, _01471_);
  nor (_01473_, _01472_, _01470_);
  and (_01474_, _01473_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_01475_, _01473_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_01476_, _01475_, _01474_);
  and (_01477_, _01461_, _42551_);
  not (_01478_, _01318_);
  nor (_01479_, _01461_, _01478_);
  nor (_01480_, _01479_, _01477_);
  and (_01481_, _01480_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_01482_, _01480_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_01483_, _01461_, _42336_);
  not (_01484_, _01297_);
  nor (_01485_, _01461_, _01484_);
  nor (_01486_, _01485_, _01483_);
  nand (_01487_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01488_, _01461_, _42429_);
  not (_01489_, _01262_);
  nor (_01490_, _01461_, _01489_);
  nor (_01491_, _01490_, _01488_);
  and (_01492_, _01491_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_01493_, _01491_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01494_, _01461_, _42589_);
  not (_01495_, _01227_);
  nor (_01496_, _01461_, _01495_);
  nor (_01497_, _01496_, _01494_);
  and (_01498_, _01497_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01499_, _01461_, _42384_);
  not (_01500_, _01201_);
  nor (_01501_, _01461_, _01500_);
  nor (_01502_, _01501_, _01499_);
  and (_01503_, _01502_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01504_, _01461_, _42464_);
  not (_01505_, _01184_);
  nor (_01506_, _01461_, _01505_);
  nor (_01507_, _01506_, _01504_);
  and (_01508_, _01507_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_01509_, _01502_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_01510_, _01509_, _01503_);
  and (_01511_, _01510_, _01508_);
  nor (_01512_, _01511_, _01503_);
  not (_01513_, _01512_);
  nor (_01514_, _01497_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_01515_, _01514_, _01498_);
  and (_01516_, _01515_, _01513_);
  nor (_01517_, _01516_, _01498_);
  nor (_01518_, _01517_, _01493_);
  or (_01519_, _01518_, _01492_);
  or (_01520_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01521_, _01520_, _01487_);
  nand (_01522_, _01521_, _01519_);
  and (_01523_, _01522_, _01487_);
  nor (_01524_, _01523_, _01482_);
  or (_01525_, _01524_, _01481_);
  and (_01526_, _01525_, _01476_);
  nor (_01527_, _01526_, _01474_);
  nor (_01528_, _01527_, _01469_);
  or (_01529_, _01528_, _01468_);
  and (_01530_, _01529_, _01467_);
  and (_01531_, _01530_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01532_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01533_, _01532_, _01531_);
  nor (_01534_, _01533_, _01465_);
  not (_01535_, _01465_);
  nor (_01536_, _01529_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01537_, _01536_, _38558_);
  and (_01538_, _01537_, _38563_);
  and (_01539_, _01538_, _38548_);
  nor (_01540_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01541_, _01540_, _01539_);
  nor (_01542_, _01541_, _01535_);
  nor (_01543_, _01542_, _01534_);
  or (_01544_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_01545_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01546_, _01545_, _01544_);
  and (_01547_, _01546_, _01543_);
  nand (_01548_, _01547_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_01549_, _01547_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_01550_, _38247_);
  and (_01551_, _01388_, _01550_);
  and (_01552_, _01551_, _01423_);
  and (_01553_, _01552_, _01451_);
  nor (_01554_, _01553_, _42317_);
  nor (_01555_, _01554_, _01457_);
  and (_01556_, _38224_, _38243_);
  nor (_01557_, _01556_, _01385_);
  not (_01558_, _01557_);
  and (_01559_, _01558_, _01461_);
  nor (_01560_, _01559_, _01555_);
  and (_01561_, _01560_, _01549_);
  and (_01562_, _01561_, _01548_);
  nor (_01563_, _01345_, _30603_);
  not (_01564_, _38621_);
  and (_01565_, _01556_, _01564_);
  and (_01566_, _01559_, _01555_);
  and (_01567_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01568_, _01567_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01569_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01570_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01571_, _01570_, _01569_);
  and (_01572_, _01571_, _01568_);
  and (_01573_, _01572_, _01467_);
  and (_01574_, _01573_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01575_, _01574_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01576_, _01575_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_01577_, _01576_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_01578_, _01577_, _38536_);
  or (_01579_, _01577_, _38536_);
  and (_01580_, _01579_, _01578_);
  and (_01581_, _01580_, _01566_);
  and (_01582_, _01454_, _42267_);
  or (_01583_, _01582_, _01581_);
  and (_01584_, _01557_, _01461_);
  and (_01585_, _01584_, _01555_);
  and (_01586_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_01587_, _01586_, _01583_);
  nor (_01588_, _01587_, _01565_);
  nand (_01589_, _01588_, _01449_);
  or (_01590_, _01589_, _01563_);
  or (_01591_, _01590_, _01562_);
  nor (_01592_, _36537_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01593_, _01592_, _42250_);
  nor (_01594_, _01593_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_01595_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_01596_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_01597_, _01596_, _01595_);
  not (_01598_, _01597_);
  nor (_01599_, _01598_, _01594_);
  and (_01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_01601_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01602_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01603_, _01602_, _01599_);
  and (_01604_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01605_, _01604_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01606_, _01605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_01607_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_01608_, _01607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01609_, _01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_01610_, _01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01611_, _01610_, _01609_);
  or (_01612_, _01611_, _01449_);
  and (_01613_, _01612_, _42882_);
  and (_39064_, _01613_, _01591_);
  and (_01614_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _42882_);
  and (_01615_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_01616_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_01617_, _36450_, _01616_);
  not (_01618_, _01617_);
  not (_01619_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_01620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_01621_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_01622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01623_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_01624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01625_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01626_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_01627_, _01626_, _01624_);
  and (_01629_, _01627_, _01625_);
  nor (_01630_, _01629_, _01624_);
  nor (_01632_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01633_, _01632_, _01623_);
  not (_01635_, _01633_);
  nor (_01636_, _01635_, _01630_);
  nor (_01638_, _01636_, _01623_);
  not (_01639_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01641_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_01642_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_01644_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_01645_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_01647_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01648_, _01647_, _01645_);
  and (_01650_, _01648_, _01644_);
  and (_01651_, _01650_, _01642_);
  and (_01653_, _01651_, _01641_);
  and (_01654_, _01653_, _01639_);
  and (_01656_, _01654_, _01638_);
  and (_01657_, _01656_, _01622_);
  and (_01659_, _01657_, _01621_);
  and (_01660_, _01659_, _01620_);
  and (_01661_, _01660_, _01619_);
  nor (_01662_, _01661_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01663_, _01661_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_01664_, _01663_, _01662_);
  not (_01665_, _01664_);
  nor (_01666_, _01660_, _01619_);
  nor (_01667_, _01666_, _01661_);
  not (_01668_, _01667_);
  nor (_01669_, _01659_, _01620_);
  or (_01670_, _01669_, _01660_);
  nor (_01671_, _01657_, _01621_);
  nor (_01672_, _01671_, _01659_);
  not (_01673_, _01672_);
  nor (_01674_, _01656_, _01622_);
  nor (_01675_, _01674_, _01657_);
  not (_01676_, _01675_);
  and (_01677_, _01653_, _01638_);
  nor (_01678_, _01677_, _01639_);
  nor (_01679_, _01678_, _01656_);
  not (_01680_, _01679_);
  not (_01681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_01682_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01683_, _01651_, _01638_);
  and (_01684_, _01683_, _01682_);
  nor (_01685_, _01684_, _01681_);
  nor (_01686_, _01685_, _01677_);
  not (_01687_, _01686_);
  and (_01688_, _01648_, _01638_);
  and (_01689_, _01688_, _01644_);
  nor (_01690_, _01689_, _01642_);
  or (_01691_, _01690_, _01683_);
  nor (_01692_, _01688_, _01644_);
  or (_01693_, _01692_, _01689_);
  and (_01694_, _01647_, _01638_);
  nor (_01695_, _01694_, _01645_);
  nor (_01696_, _01695_, _01688_);
  not (_01697_, _01696_);
  not (_01698_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01699_, _01638_, _01698_);
  nor (_01700_, _01638_, _01698_);
  nor (_01701_, _01700_, _01699_);
  not (_01702_, _01701_);
  and (_01703_, _00706_, _00635_);
  and (_01704_, _01703_, _00708_);
  not (_01705_, _01704_);
  or (_01706_, _00711_, _00658_);
  and (_01707_, _01706_, _00708_);
  not (_01708_, _00708_);
  and (_01709_, _00651_, _00644_);
  nor (_01710_, _01709_, _00683_);
  nor (_01711_, _01710_, _01708_);
  nor (_01712_, _01711_, _01707_);
  and (_01713_, _01712_, _01705_);
  and (_01714_, _00713_, _00704_);
  and (_01715_, _00708_, _00661_);
  nor (_01716_, _01715_, _01714_);
  not (_01717_, _00660_);
  nor (_01718_, _00658_, _00707_);
  nor (_01719_, _01718_, _01717_);
  not (_01720_, _00667_);
  and (_01721_, _00678_, _00635_);
  nor (_01722_, _01721_, _00645_);
  nor (_01723_, _01722_, _01720_);
  nor (_01724_, _01723_, _01719_);
  and (_01725_, _01724_, _01716_);
  and (_01726_, _01725_, _01713_);
  and (_01727_, _01726_, _00688_);
  not (_01728_, _00673_);
  and (_01729_, _00703_, _00658_);
  nor (_01730_, _01729_, _00646_);
  and (_01731_, _00657_, _00689_);
  and (_01732_, _00694_, _01731_);
  and (_01733_, _00635_, _00642_);
  and (_01734_, _00649_, _38185_);
  and (_01735_, _01734_, _01733_);
  nor (_01736_, _01735_, _01732_);
  and (_01737_, _01736_, _01730_);
  and (_01738_, _01737_, _01728_);
  and (_01739_, _00672_, _00635_);
  nor (_01740_, _00650_, _00639_);
  and (_01741_, _00683_, _37905_);
  nor (_01742_, _01741_, _00679_);
  nor (_01743_, _01742_, _01740_);
  nor (_01744_, _01743_, _01739_);
  and (_01745_, _01744_, _01738_);
  and (_01746_, _00683_, _00640_);
  and (_01747_, _00678_, _00644_);
  and (_01748_, _01747_, _00708_);
  nor (_01749_, _01748_, _01746_);
  and (_01750_, _00711_, _00660_);
  not (_01751_, _00703_);
  nor (_01752_, _01703_, _00685_);
  nor (_01753_, _01752_, _01751_);
  nor (_01754_, _01753_, _01750_);
  and (_01755_, _01754_, _01749_);
  nor (_01756_, _00712_, _00663_);
  nor (_01757_, _01733_, _00658_);
  nor (_01758_, _01757_, _38210_);
  nor (_01759_, _01758_, _00699_);
  and (_01760_, _01759_, _01756_);
  and (_01761_, _01760_, _01755_);
  and (_01762_, _01761_, _01745_);
  not (_01763_, _00653_);
  not (_01764_, _00671_);
  and (_01765_, _00657_, _00706_);
  and (_01766_, _01765_, _00640_);
  nor (_01767_, _01766_, _00709_);
  and (_01768_, _01767_, _01764_);
  and (_01769_, _01768_, _01763_);
  and (_01770_, _00670_, _00635_);
  nor (_01771_, _01770_, _00652_);
  nor (_01772_, _01771_, _01717_);
  not (_01773_, _01772_);
  not (_01774_, _01765_);
  nor (_01775_, _00660_, _00650_);
  nor (_01776_, _01775_, _01774_);
  and (_01777_, _00669_, _00644_);
  not (_01778_, _01777_);
  nor (_01779_, _00708_, _00660_);
  nor (_01780_, _01779_, _01778_);
  nor (_01781_, _01780_, _01776_);
  and (_01782_, _01781_, _01773_);
  and (_01783_, _01782_, _01769_);
  and (_01784_, _01783_, _01762_);
  and (_01785_, _01784_, _01727_);
  not (_01786_, _01785_);
  nor (_01787_, _01627_, _01625_);
  nor (_01788_, _01787_, _01629_);
  nand (_01789_, _01788_, _01786_);
  and (_01790_, _00657_, _00642_);
  and (_01791_, _01790_, _00640_);
  and (_01792_, _01703_, _00667_);
  or (_01793_, _01792_, _01707_);
  or (_01794_, _00686_, _00663_);
  or (_01795_, _01794_, _01793_);
  or (_01796_, _01795_, _01791_);
  not (_01797_, _00699_);
  nand (_01798_, _01769_, _01797_);
  or (_01799_, _01798_, _01796_);
  nor (_01800_, _01799_, _01785_);
  not (_01801_, _01800_);
  nor (_01802_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01803_, _01802_, _01625_);
  and (_01804_, _01803_, _01801_);
  or (_01805_, _01788_, _01786_);
  and (_01806_, _01805_, _01789_);
  nand (_01807_, _01806_, _01804_);
  and (_01808_, _01807_, _01789_);
  not (_01809_, _01808_);
  and (_01810_, _01635_, _01630_);
  nor (_01811_, _01810_, _01636_);
  and (_01812_, _01811_, _01809_);
  and (_01813_, _01812_, _01702_);
  not (_01814_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_01815_, _01699_, _01814_);
  or (_01816_, _01815_, _01694_);
  and (_01817_, _01816_, _01813_);
  and (_01818_, _01817_, _01697_);
  and (_01819_, _01818_, _01693_);
  and (_01820_, _01819_, _01691_);
  nor (_01821_, _01683_, _01682_);
  or (_01822_, _01821_, _01684_);
  and (_01823_, _01822_, _01820_);
  and (_01824_, _01823_, _01687_);
  and (_01825_, _01824_, _01680_);
  and (_01826_, _01825_, _01676_);
  and (_01827_, _01826_, _01673_);
  and (_01828_, _01827_, _01670_);
  nand (_01829_, _01828_, _01668_);
  nand (_01830_, _01829_, _01665_);
  or (_01831_, _01829_, _01665_);
  and (_01832_, _01831_, _01830_);
  or (_01833_, _01832_, _01618_);
  or (_01834_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_01835_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_01836_, _01835_, _01834_);
  and (_01837_, _01836_, _01833_);
  or (_39066_, _01837_, _01615_);
  nor (_01838_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_39067_, _01838_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_39068_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _42882_);
  not (_01839_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor (_01840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_01841_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01842_, _01841_, _01840_);
  not (_01843_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_01844_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_01845_, _01844_, _01843_);
  and (_01846_, _01845_, _01842_);
  and (_01847_, _01846_, _01839_);
  and (_01848_, \oc8051_top_1.oc8051_rom1.ea_int , _36418_);
  nand (_01849_, _01848_, _36450_);
  nand (_01850_, _01849_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_01851_, _01850_, _01847_);
  and (_39069_, _01851_, _42882_);
  and (_01852_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_01853_, _01852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_39071_, _01853_, _42882_);
  nor (_01854_, _01594_, _42250_);
  or (_01855_, _01785_, _36646_);
  nor (_01856_, _01800_, _36570_);
  nand (_01857_, _01785_, _36646_);
  and (_01858_, _01857_, _01855_);
  nand (_01859_, _01858_, _01856_);
  and (_01860_, _01859_, _01855_);
  nor (_01861_, _01860_, _42250_);
  and (_01862_, _01861_, _36494_);
  nor (_01863_, _01861_, _36494_);
  nor (_01864_, _01863_, _01862_);
  nor (_01865_, _01864_, _01854_);
  and (_01866_, _36657_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_01867_, _01866_, _01854_);
  and (_01868_, _01867_, _01799_);
  or (_01869_, _01868_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01870_, _01869_, _01865_);
  and (_39072_, _01870_, _42882_);
  nor (_01871_, _38179_, _36767_);
  and (_01872_, _37313_, _37062_);
  and (_01873_, _01872_, _01871_);
  nand (_01874_, _01342_, _38101_);
  nor (_01875_, _01874_, _37861_);
  not (_01876_, _38206_);
  and (_01877_, _01876_, _37586_);
  and (_01878_, _01877_, _01875_);
  and (_39075_, _01878_, _01873_);
  nor (_01879_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_01880_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_01881_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_39078_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _42882_);
  and (_01882_, _39078_, _01881_);
  or (_39076_, _01882_, _01880_);
  not (_01883_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01884_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01885_, _01884_, _01883_);
  and (_01886_, _01884_, _01883_);
  nor (_01887_, _01886_, _01885_);
  not (_01888_, _01887_);
  and (_01889_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01890_, _01889_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01891_, _01889_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01892_, _01891_, _01890_);
  or (_01893_, _01892_, _01884_);
  and (_01894_, _01893_, _01888_);
  nor (_01895_, _01885_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01896_, _01885_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_01897_, _01896_, _01895_);
  or (_01898_, _01890_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_39080_, _01898_, _42882_);
  and (_01899_, _39080_, _01897_);
  and (_39079_, _01899_, _01894_);
  not (_01900_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_01901_, _01594_, _01900_);
  and (_01902_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_01903_, _01901_);
  and (_01904_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_01905_, _01904_, _01902_);
  and (_39081_, _01905_, _42882_);
  and (_01906_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01907_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_01908_, _01907_, _01906_);
  and (_39082_, _01908_, _42882_);
  and (_01909_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_01910_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_01911_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _01910_);
  and (_01912_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_01913_, _01912_, _01909_);
  and (_39083_, _01913_, _42882_);
  and (_01914_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_01915_, _01914_, _01911_);
  and (_39084_, _01915_, _42882_);
  or (_01916_, _01910_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_39086_, _01916_, _42882_);
  not (_01917_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_01918_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01919_, _01918_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_01920_, _01910_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_01921_, _01920_, _42882_);
  and (_39087_, _01921_, _01919_);
  or (_01922_, _01910_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_39088_, _01922_, _42882_);
  nor (_01923_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_01924_, _01923_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_01925_, _01924_, _42882_);
  and (_01926_, _39078_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_39089_, _01926_, _01925_);
  and (_01927_, _01900_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_01928_, _01927_, _01924_);
  and (_39090_, _01928_, _42882_);
  nand (_01929_, _01924_, _38621_);
  or (_01930_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_01931_, _01930_, _42882_);
  and (_39091_, _01931_, _01929_);
  nand (_01932_, _38257_, _42882_);
  nor (_39092_, _01932_, _38398_);
  or (_01933_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_01934_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_01935_, _01934_, _42882_);
  and (_39128_, _01935_, _01933_);
  or (_01936_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_01937_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_01938_, _01336_, _01937_);
  and (_01939_, _01938_, _42882_);
  and (_39129_, _01939_, _01936_);
  or (_01940_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_01941_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_01942_, _01336_, _01941_);
  and (_01943_, _01942_, _42882_);
  and (_39130_, _01943_, _01940_);
  or (_01944_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_01945_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_01946_, _01336_, _01945_);
  and (_01947_, _01946_, _42882_);
  and (_39131_, _01947_, _01944_);
  or (_01948_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_01949_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_01950_, _01336_, _01949_);
  and (_01951_, _01950_, _42882_);
  and (_39132_, _01951_, _01948_);
  or (_01952_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_01953_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_01954_, _01336_, _01953_);
  and (_01955_, _01954_, _42882_);
  and (_39134_, _01955_, _01952_);
  or (_01956_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_01957_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01958_, _01957_, _42882_);
  and (_39135_, _01958_, _01956_);
  or (_01959_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_01960_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_01961_, _01336_, _01960_);
  and (_01962_, _01961_, _42882_);
  and (_39136_, _01962_, _01959_);
  or (_01963_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_01964_, _01336_, _38552_);
  and (_01965_, _01964_, _42882_);
  and (_39137_, _01965_, _01963_);
  or (_01966_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_01967_, _01336_, _38558_);
  and (_01968_, _01967_, _42882_);
  and (_39138_, _01968_, _01966_);
  or (_01969_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_01970_, _01336_, _38563_);
  and (_01971_, _01970_, _42882_);
  and (_39139_, _01971_, _01969_);
  or (_01972_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_01973_, _01336_, _38548_);
  and (_01974_, _01973_, _42882_);
  and (_39140_, _01974_, _01972_);
  or (_01975_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_01976_, _01336_, _38569_);
  and (_01977_, _01976_, _42882_);
  and (_39141_, _01977_, _01975_);
  or (_01978_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_01979_, _01336_, _38544_);
  and (_01980_, _01979_, _42882_);
  and (_39142_, _01980_, _01978_);
  or (_01981_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_01982_, _01336_, _38540_);
  and (_01983_, _01982_, _42882_);
  and (_39143_, _01983_, _01981_);
  and (_01984_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_01985_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_01986_, _01985_, _01984_);
  and (_39148_, _01986_, _42882_);
  and (_01987_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_01988_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_01989_, _01988_, _01987_);
  and (_39149_, _01989_, _42882_);
  and (_01990_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_01991_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_01992_, _01991_, _01990_);
  and (_39150_, _01992_, _42882_);
  and (_01993_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_01994_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_01995_, _01994_, _01993_);
  and (_39151_, _01995_, _42882_);
  and (_01996_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_01997_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or (_01998_, _01997_, _01996_);
  and (_39152_, _01998_, _42882_);
  and (_01999_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_02000_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or (_02001_, _02000_, _01999_);
  and (_39153_, _02001_, _42882_);
  and (_02002_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_02003_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or (_02004_, _02003_, _02002_);
  and (_39154_, _02004_, _42882_);
  and (_02005_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_02006_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or (_02007_, _02006_, _02005_);
  and (_39155_, _02007_, _42882_);
  and (_02008_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_02009_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or (_02010_, _02009_, _02008_);
  and (_39156_, _02010_, _42882_);
  and (_02011_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_02012_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or (_02013_, _02012_, _02011_);
  and (_39157_, _02013_, _42882_);
  and (_02014_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_02015_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or (_02016_, _02015_, _02014_);
  and (_39159_, _02016_, _42882_);
  and (_02017_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_02018_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or (_02019_, _02018_, _02017_);
  and (_39160_, _02019_, _42882_);
  and (_02020_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_02021_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or (_02022_, _02021_, _02020_);
  and (_39161_, _02022_, _42882_);
  and (_02023_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_02024_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or (_02025_, _02024_, _02023_);
  and (_39162_, _02025_, _42882_);
  and (_02026_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_02027_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or (_02028_, _02027_, _02026_);
  and (_39163_, _02028_, _42882_);
  and (_39339_, _37960_, _42882_);
  and (_39340_, _38190_, _42882_);
  and (_39341_, _38167_, _42882_);
  nor (_39342_, _42273_, rst);
  and (_02029_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02030_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_02031_, _02030_, _02029_);
  and (_39343_, _02031_, _42882_);
  and (_02032_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_02033_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_02034_, _02033_, _01901_);
  or (_02035_, _02034_, _02032_);
  and (_39344_, _02035_, _42882_);
  and (_02036_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02037_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_02038_, _02037_, _02036_);
  and (_39345_, _02038_, _42882_);
  and (_02039_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02040_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_02041_, _02040_, _02039_);
  and (_39346_, _02041_, _42882_);
  and (_02042_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02043_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_02044_, _02043_, _02042_);
  and (_39348_, _02044_, _42882_);
  and (_02045_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02046_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_02047_, _02046_, _02045_);
  and (_39349_, _02047_, _42882_);
  and (_02048_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02049_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_02050_, _02049_, _02048_);
  and (_39350_, _02050_, _42882_);
  and (_02051_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02052_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_02053_, _02052_, _02051_);
  and (_39351_, _02053_, _42882_);
  and (_02054_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_02055_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_02056_, _02055_, _02054_);
  and (_39352_, _02056_, _42882_);
  and (_02057_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_02058_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_02059_, _02058_, _02057_);
  and (_39353_, _02059_, _42882_);
  and (_02060_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_02061_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_02062_, _02061_, _02060_);
  and (_39354_, _02062_, _42882_);
  and (_02063_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_02064_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_02065_, _02064_, _02063_);
  and (_39355_, _02065_, _42882_);
  and (_02066_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_02067_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_02068_, _02067_, _02066_);
  and (_39356_, _02068_, _42882_);
  and (_02069_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_02070_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_02071_, _02070_, _02069_);
  and (_39357_, _02071_, _42882_);
  and (_02072_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_02073_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_02074_, _02073_, _02072_);
  and (_39359_, _02074_, _42882_);
  and (_02075_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_02076_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_02077_, _02076_, _02075_);
  and (_39360_, _02077_, _42882_);
  and (_02078_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_02079_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_02080_, _02079_, _02078_);
  and (_39361_, _02080_, _42882_);
  and (_02081_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_02082_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_02083_, _02082_, _02081_);
  and (_39362_, _02083_, _42882_);
  and (_02084_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_02085_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_02086_, _02085_, _02084_);
  and (_39363_, _02086_, _42882_);
  and (_02087_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_02088_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_02089_, _02088_, _02087_);
  and (_39364_, _02089_, _42882_);
  and (_02090_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_02091_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_02092_, _02091_, _02090_);
  and (_39365_, _02092_, _42882_);
  and (_02093_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_02094_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_02095_, _02094_, _02093_);
  and (_39366_, _02095_, _42882_);
  and (_02096_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_02097_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_02098_, _02097_, _02096_);
  and (_39367_, _02098_, _42882_);
  and (_02099_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_02100_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_02101_, _02100_, _02099_);
  and (_39368_, _02101_, _42882_);
  and (_02102_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_02103_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_02104_, _02103_, _02102_);
  and (_39370_, _02104_, _42882_);
  and (_02105_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_02106_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_02107_, _02106_, _02105_);
  and (_39371_, _02107_, _42882_);
  and (_02110_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_02112_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_02114_, _02112_, _02110_);
  and (_39372_, _02114_, _42882_);
  and (_02117_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_02119_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_02121_, _02119_, _02117_);
  and (_39373_, _02121_, _42882_);
  and (_02124_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_02126_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_02128_, _02126_, _02124_);
  and (_39374_, _02128_, _42882_);
  and (_02131_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_02133_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_02135_, _02133_, _02131_);
  and (_39375_, _02135_, _42882_);
  and (_02138_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_02140_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_02142_, _02140_, _02138_);
  and (_39376_, _02142_, _42882_);
  nor (_39377_, _42476_, rst);
  and (_39379_, _42398_, _42882_);
  nor (_39380_, _42602_, rst);
  nor (_39381_, _42444_, rst);
  nor (_39382_, _42356_, rst);
  nor (_39383_, _42564_, rst);
  and (_39385_, _42505_, _42882_);
  and (_39401_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _42882_);
  and (_39402_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _42882_);
  and (_39403_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _42882_);
  and (_39404_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _42882_);
  and (_39405_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _42882_);
  and (_39407_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _42882_);
  and (_39408_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _42882_);
  not (_02158_, _01450_);
  and (_02159_, _02158_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_02160_, _01566_, _42465_);
  and (_02161_, _01454_, _01505_);
  or (_02162_, _02161_, _02160_);
  or (_02163_, _01507_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_02164_, _01508_);
  and (_02165_, _01560_, _02164_);
  and (_02166_, _02165_, _02163_);
  or (_02167_, _02166_, _02162_);
  or (_02168_, _01585_, _01556_);
  and (_02169_, _02168_, _31783_);
  or (_02170_, _02169_, _02167_);
  and (_02171_, _02170_, _01449_);
  or (_02172_, _02171_, _02159_);
  and (_39409_, _02172_, _42882_);
  and (_02173_, _02158_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_02174_, _01566_, _42385_);
  and (_02175_, _01454_, _01500_);
  or (_02176_, _02175_, _02174_);
  or (_02177_, _01510_, _01508_);
  not (_02178_, _01511_);
  and (_02179_, _01560_, _02178_);
  and (_02180_, _02179_, _02177_);
  or (_02181_, _02180_, _02176_);
  and (_02182_, _02168_, _32469_);
  or (_02183_, _02182_, _02181_);
  and (_02184_, _02183_, _01449_);
  or (_02185_, _02184_, _02173_);
  and (_39410_, _02185_, _42882_);
  and (_02186_, _02168_, _33165_);
  or (_02187_, _01515_, _01513_);
  not (_02188_, _01516_);
  and (_02189_, _01560_, _02188_);
  nand (_02190_, _02189_, _02187_);
  and (_02191_, _01566_, _42590_);
  and (_02192_, _01454_, _01495_);
  and (_02193_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_02194_, _02193_, _02192_);
  nor (_02195_, _02194_, _02191_);
  and (_02196_, _02195_, _02190_);
  nand (_02197_, _02196_, _01449_);
  or (_02198_, _02197_, _02186_);
  not (_02199_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02200_, _01594_, _02199_);
  and (_02201_, _01594_, _02199_);
  nor (_02202_, _02201_, _02200_);
  or (_02203_, _02202_, _01449_);
  and (_02204_, _02203_, _42882_);
  and (_39411_, _02204_, _02198_);
  and (_02205_, _02168_, _33916_);
  or (_02206_, _01493_, _01492_);
  or (_02207_, _02206_, _01517_);
  nand (_02208_, _02206_, _01517_);
  and (_02209_, _02208_, _01560_);
  nand (_02210_, _02209_, _02207_);
  and (_02211_, _01566_, _42430_);
  and (_02212_, _01454_, _01489_);
  and (_02213_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_02214_, _02213_, _02212_);
  nor (_02215_, _02214_, _02211_);
  and (_02216_, _02215_, _02210_);
  nand (_02217_, _02216_, _01449_);
  or (_02218_, _02217_, _02205_);
  and (_02219_, _02200_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02220_, _02200_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02221_, _02220_, _02219_);
  or (_02222_, _02221_, _01449_);
  and (_02223_, _02222_, _42882_);
  and (_39412_, _02223_, _02218_);
  and (_02224_, _02168_, _34678_);
  or (_02225_, _01521_, _01519_);
  and (_02226_, _01560_, _01522_);
  and (_02227_, _02226_, _02225_);
  and (_02228_, _01566_, _42337_);
  and (_02229_, _01454_, _01484_);
  and (_02230_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_02231_, _02230_, _02229_);
  or (_02232_, _02231_, _02228_);
  nor (_02233_, _02232_, _02227_);
  nand (_02234_, _02233_, _01449_);
  or (_02235_, _02234_, _02224_);
  and (_02236_, _02219_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02237_, _02219_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02238_, _02237_, _02236_);
  or (_02239_, _02238_, _01449_);
  and (_02240_, _02239_, _42882_);
  and (_39413_, _02240_, _02235_);
  and (_02241_, _02168_, _35472_);
  or (_02242_, _01482_, _01481_);
  nand (_02243_, _02242_, _01523_);
  or (_02244_, _02242_, _01523_);
  and (_02245_, _02244_, _01560_);
  nand (_02246_, _02245_, _02243_);
  and (_02247_, _01566_, _42552_);
  and (_02248_, _01454_, _01478_);
  and (_02249_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_02250_, _02249_, _02248_);
  nor (_02251_, _02250_, _02247_);
  and (_02252_, _02251_, _02246_);
  nand (_02253_, _02252_, _01449_);
  or (_02254_, _02253_, _02241_);
  nor (_02255_, _02236_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02256_, _02255_, _01599_);
  or (_02257_, _02256_, _01449_);
  and (_02258_, _02257_, _42882_);
  and (_39414_, _02258_, _02254_);
  nor (_02259_, _01599_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02260_, _01599_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_02261_, _02260_, _02259_);
  or (_02262_, _02261_, _01449_);
  and (_02263_, _02262_, _42882_);
  and (_02264_, _02168_, _36190_);
  and (_02265_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02266_, _01454_, _01471_);
  and (_02267_, _01566_, _42524_);
  or (_02268_, _02267_, _02266_);
  or (_02269_, _02268_, _02265_);
  or (_02270_, _01525_, _01476_);
  not (_02271_, _01526_);
  and (_02272_, _01560_, _02271_);
  and (_02273_, _02272_, _02270_);
  nor (_02274_, _02273_, _02269_);
  nand (_02275_, _02274_, _01449_);
  or (_02276_, _02275_, _02264_);
  and (_39415_, _02276_, _02263_);
  and (_02277_, _02168_, _30614_);
  or (_02278_, _01468_, _01469_);
  or (_02279_, _02278_, _01527_);
  nand (_02280_, _02278_, _01527_);
  and (_02281_, _02280_, _01560_);
  and (_02282_, _02281_, _02279_);
  and (_02283_, _01454_, _01463_);
  and (_02284_, _01566_, _42267_);
  and (_02285_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_02286_, _02285_, _02284_);
  nor (_02287_, _02286_, _02283_);
  nand (_02288_, _02287_, _01449_);
  or (_02289_, _02288_, _02282_);
  or (_02290_, _02289_, _02277_);
  nor (_02291_, _02260_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_02292_, _02260_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_02293_, _02292_, _02291_);
  or (_02294_, _02293_, _01449_);
  and (_02295_, _02294_, _42882_);
  and (_39416_, _02295_, _02290_);
  nor (_02296_, _01345_, _31782_);
  not (_02297_, _38660_);
  and (_02298_, _01556_, _02297_);
  and (_02299_, _01529_, _38552_);
  nor (_02300_, _01529_, _38552_);
  nor (_02301_, _02300_, _02299_);
  nand (_02302_, _02301_, _01535_);
  or (_02303_, _02301_, _01535_);
  and (_02304_, _02303_, _01560_);
  and (_02305_, _02304_, _02302_);
  and (_02306_, _01566_, _00689_);
  and (_02307_, _01454_, _42465_);
  or (_02308_, _02307_, _02306_);
  and (_02309_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_02310_, _02309_, _02308_);
  nand (_02311_, _02310_, _01449_);
  or (_02312_, _02311_, _02305_);
  or (_02313_, _02312_, _02298_);
  or (_02314_, _02313_, _02296_);
  or (_02315_, _02292_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_02316_, _01601_, _01599_);
  and (_02317_, _02316_, _02315_);
  or (_02318_, _02317_, _01449_);
  and (_02319_, _02318_, _42882_);
  and (_39418_, _02319_, _02314_);
  nor (_02320_, _01345_, _32458_);
  and (_02321_, _01529_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02322_, _02321_, _01535_);
  and (_02323_, _01536_, _01465_);
  nor (_02324_, _02323_, _02322_);
  nand (_02325_, _02324_, _38558_);
  or (_02326_, _02324_, _38558_);
  and (_02327_, _02326_, _01560_);
  and (_02328_, _02327_, _02325_);
  not (_02329_, _38693_);
  nand (_02330_, _01556_, _02329_);
  and (_02331_, _01566_, _00656_);
  and (_02332_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_02333_, _01454_, _42385_);
  or (_02334_, _02333_, _02332_);
  nor (_02335_, _02334_, _02331_);
  and (_02336_, _02335_, _02330_);
  nand (_02337_, _02336_, _01449_);
  or (_02338_, _02337_, _02328_);
  or (_02339_, _02338_, _02320_);
  nand (_02340_, _02316_, _01681_);
  or (_02341_, _02316_, _01681_);
  and (_02342_, _02341_, _02340_);
  or (_02343_, _02342_, _01449_);
  and (_02344_, _02343_, _42882_);
  and (_39419_, _02344_, _02339_);
  nor (_02345_, _01345_, _33154_);
  and (_02346_, _01537_, _01465_);
  and (_02347_, _02322_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_02348_, _02347_, _02346_);
  nand (_02349_, _02348_, _38563_);
  or (_02350_, _02348_, _38563_);
  and (_02351_, _02350_, _01560_);
  and (_02352_, _02351_, _02349_);
  not (_02353_, _38724_);
  and (_02354_, _01556_, _02353_);
  and (_02355_, _01566_, _00634_);
  and (_02357_, _01454_, _42590_);
  or (_02358_, _02357_, _02355_);
  and (_02359_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_02360_, _02359_, _02358_);
  nor (_02361_, _02360_, _02354_);
  nand (_02362_, _02361_, _01449_);
  or (_02363_, _02362_, _02352_);
  or (_02364_, _02363_, _02345_);
  nor (_02365_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_02366_, _02365_, _01604_);
  or (_02367_, _02366_, _01449_);
  and (_02368_, _02367_, _42882_);
  and (_39420_, _02368_, _02364_);
  nor (_02369_, _01345_, _33906_);
  and (_02370_, _01530_, _01535_);
  and (_02371_, _01538_, _01465_);
  nor (_02372_, _02371_, _02370_);
  nand (_02373_, _02372_, _38548_);
  or (_02374_, _02372_, _38548_);
  and (_02375_, _02374_, _01560_);
  and (_02376_, _02375_, _02373_);
  not (_02377_, _38756_);
  and (_02378_, _01556_, _02377_);
  and (_02379_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02380_, _01573_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_02381_, _02380_, _01574_);
  and (_02382_, _02381_, _01566_);
  and (_02383_, _01454_, _42430_);
  or (_02384_, _02383_, _02382_);
  or (_02385_, _02384_, _02379_);
  nor (_02386_, _02385_, _02378_);
  nand (_02387_, _02386_, _01449_);
  or (_02388_, _02387_, _02376_);
  or (_02389_, _02388_, _02369_);
  nor (_02390_, _01604_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02391_, _02390_, _01605_);
  or (_02392_, _02391_, _01449_);
  and (_02393_, _02392_, _42882_);
  and (_39421_, _02393_, _02389_);
  nor (_02394_, _01345_, _34667_);
  and (_02395_, _01531_, _01535_);
  and (_02396_, _01539_, _01465_);
  nor (_02397_, _02396_, _02395_);
  nand (_02398_, _02397_, _38569_);
  or (_02399_, _02397_, _38569_);
  and (_02400_, _02399_, _01560_);
  and (_02401_, _02400_, _02398_);
  not (_02402_, _38787_);
  nand (_02403_, _01556_, _02402_);
  and (_02404_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_02405_, _01574_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_02406_, _02405_, _01575_);
  and (_02407_, _02406_, _01566_);
  and (_02408_, _01454_, _42337_);
  or (_02409_, _02408_, _02407_);
  nor (_02410_, _02409_, _02404_);
  and (_02411_, _02410_, _02403_);
  nand (_02412_, _02411_, _01449_);
  or (_02413_, _02412_, _02401_);
  or (_02414_, _02413_, _02394_);
  nor (_02415_, _01605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_02416_, _02415_, _01606_);
  or (_02417_, _02416_, _01449_);
  and (_02418_, _02417_, _42882_);
  and (_39422_, _02418_, _02414_);
  nor (_02419_, _01345_, _35461_);
  and (_02420_, _02395_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_02421_, _02396_, _38569_);
  nor (_02422_, _02421_, _02420_);
  nand (_02423_, _02422_, _38544_);
  or (_02424_, _02422_, _38544_);
  and (_02425_, _02424_, _01560_);
  and (_02426_, _02425_, _02423_);
  not (_02427_, _38821_);
  nand (_02428_, _01556_, _02427_);
  and (_02429_, _01454_, _42552_);
  nor (_02430_, _01575_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_02431_, _02430_, _01576_);
  and (_02432_, _02431_, _01566_);
  and (_02433_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_02434_, _02433_, _02432_);
  nor (_02435_, _02434_, _02429_);
  and (_02436_, _02435_, _02428_);
  nand (_02437_, _02436_, _01449_);
  or (_02438_, _02437_, _02426_);
  or (_02439_, _02438_, _02419_);
  nor (_02440_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_02441_, _02440_, _01607_);
  or (_02442_, _02441_, _01449_);
  and (_02443_, _02442_, _42882_);
  and (_39423_, _02443_, _02439_);
  nor (_02444_, _01345_, _36179_);
  nor (_02445_, _01543_, _38540_);
  and (_02446_, _01543_, _38540_);
  or (_02447_, _02446_, _02445_);
  and (_02448_, _02447_, _01560_);
  and (_02449_, _01556_, _38847_);
  or (_02450_, _01576_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02451_, _02450_, _01577_);
  and (_02452_, _02451_, _01566_);
  and (_02453_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_02454_, _01454_, _42524_);
  or (_02455_, _02454_, _02453_);
  or (_02456_, _02455_, _02452_);
  nor (_02457_, _02456_, _02449_);
  nand (_02458_, _02457_, _01449_);
  or (_02459_, _02458_, _02448_);
  or (_02460_, _02459_, _02444_);
  nor (_02461_, _01607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_02462_, _02461_, _01608_);
  or (_02463_, _02462_, _01449_);
  and (_02464_, _02463_, _42882_);
  and (_39424_, _02464_, _02460_);
  and (_02465_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_02466_, _01803_, _01801_);
  nor (_02467_, _02466_, _01804_);
  or (_02468_, _02467_, _01618_);
  or (_02469_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_02470_, _02469_, _01835_);
  and (_02471_, _02470_, _02468_);
  or (_39425_, _02471_, _02465_);
  or (_02472_, _01806_, _01804_);
  and (_02473_, _02472_, _01807_);
  or (_02474_, _02473_, _01618_);
  or (_02475_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_02476_, _02475_, _01835_);
  and (_02477_, _02476_, _02474_);
  and (_02478_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39426_, _02478_, _02477_);
  or (_02479_, _01811_, _01809_);
  nor (_02480_, _01812_, _01618_);
  and (_02481_, _02480_, _02479_);
  nor (_02482_, _01617_, _01941_);
  or (_02483_, _02482_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02484_, _02483_, _02481_);
  or (_02485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _36418_);
  and (_02486_, _02485_, _42882_);
  and (_39427_, _02486_, _02484_);
  and (_02487_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02488_, _01812_, _01702_);
  nor (_02489_, _02488_, _01813_);
  or (_02490_, _02489_, _01618_);
  or (_02491_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_02492_, _02491_, _01835_);
  and (_02493_, _02492_, _02490_);
  or (_39429_, _02493_, _02487_);
  and (_02494_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02495_, _01816_, _01813_);
  nor (_02496_, _02495_, _01817_);
  or (_02497_, _02496_, _01618_);
  or (_02498_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_02499_, _02498_, _01835_);
  and (_02500_, _02499_, _02497_);
  or (_39430_, _02500_, _02494_);
  and (_02501_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02502_, _01817_, _01697_);
  nor (_02503_, _02502_, _01818_);
  or (_02504_, _02503_, _01618_);
  or (_02505_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_02506_, _02505_, _01835_);
  and (_02507_, _02506_, _02504_);
  or (_39431_, _02507_, _02501_);
  nor (_02508_, _01818_, _01693_);
  nor (_02509_, _02508_, _01819_);
  or (_02510_, _02509_, _01618_);
  or (_02511_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_02512_, _02511_, _01835_);
  and (_02513_, _02512_, _02510_);
  and (_02514_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39432_, _02514_, _02513_);
  nor (_02515_, _01819_, _01691_);
  nor (_02516_, _02515_, _01820_);
  or (_02517_, _02516_, _01618_);
  or (_02518_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_02519_, _02518_, _01835_);
  and (_02520_, _02519_, _02517_);
  and (_02521_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_39433_, _02521_, _02520_);
  and (_02522_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_02523_, _01822_, _01820_);
  nor (_02524_, _02523_, _01823_);
  or (_02525_, _02524_, _01618_);
  or (_02526_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02527_, _02526_, _01835_);
  and (_02528_, _02527_, _02525_);
  or (_39434_, _02528_, _02522_);
  and (_02529_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_02530_, _01823_, _01687_);
  nor (_02531_, _02530_, _01824_);
  or (_02532_, _02531_, _01618_);
  or (_02533_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_02534_, _02533_, _01835_);
  and (_02535_, _02534_, _02532_);
  or (_39435_, _02535_, _02529_);
  nor (_02536_, _01824_, _01680_);
  nor (_02537_, _02536_, _01825_);
  or (_02538_, _02537_, _01618_);
  or (_02539_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_02540_, _02539_, _01835_);
  and (_02541_, _02540_, _02538_);
  and (_02543_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_39436_, _02543_, _02541_);
  nor (_02544_, _01825_, _01676_);
  nor (_02545_, _02544_, _01826_);
  or (_02546_, _02545_, _01618_);
  or (_02547_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_02548_, _02547_, _01835_);
  and (_02549_, _02548_, _02546_);
  and (_02550_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_39437_, _02550_, _02549_);
  nor (_02551_, _01826_, _01673_);
  nor (_02552_, _02551_, _01827_);
  or (_02553_, _02552_, _01618_);
  or (_02554_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_02555_, _02554_, _01835_);
  and (_02556_, _02555_, _02553_);
  and (_02557_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_39438_, _02557_, _02556_);
  and (_02558_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_02559_, _01827_, _01670_);
  nor (_02560_, _02559_, _01828_);
  or (_02561_, _02560_, _01618_);
  or (_02562_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_02564_, _02562_, _01835_);
  and (_02565_, _02564_, _02561_);
  or (_39440_, _02565_, _02558_);
  or (_02566_, _01828_, _01668_);
  and (_02567_, _02566_, _01829_);
  or (_02568_, _02567_, _01618_);
  or (_02569_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02570_, _02569_, _01835_);
  and (_02571_, _02570_, _02568_);
  and (_02572_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_39441_, _02572_, _02571_);
  and (_02574_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_02575_, _02574_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_39442_, _02575_, _42882_);
  and (_02576_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_02577_, _02576_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_39443_, _02577_, _42882_);
  and (_02578_, _01846_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_02579_, _02578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_39444_, _02579_, _42882_);
  and (_02580_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_02581_, _02580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39445_, _02581_, _42882_);
  and (_02582_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_02583_, _02582_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_39446_, _02583_, _42882_);
  and (_02584_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_02585_, _02584_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_39447_, _02585_, _42882_);
  and (_02586_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_02587_, _02586_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_39448_, _02587_, _42882_);
  nor (_02588_, _01800_, _42250_);
  nand (_02589_, _02588_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_02590_, _02588_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_02591_, _02590_, _01835_);
  and (_39449_, _02591_, _02589_);
  or (_02592_, _01858_, _01856_);
  and (_02593_, _02592_, _01859_);
  or (_02594_, _02593_, _42250_);
  or (_02595_, _36450_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_02596_, _02595_, _01835_);
  and (_39450_, _02596_, _02594_);
  and (_02597_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_02598_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_02599_, _02598_, _39078_);
  or (_39466_, _02599_, _02597_);
  and (_02600_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_02601_, _02033_, _39078_);
  or (_39467_, _02601_, _02600_);
  and (_02602_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_02603_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_02604_, _02603_, _39078_);
  or (_39468_, _02604_, _02602_);
  and (_02605_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_02606_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_02607_, _02606_, _39078_);
  or (_39469_, _02607_, _02605_);
  and (_02608_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_02609_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_02610_, _02609_, _39078_);
  or (_39470_, _02610_, _02608_);
  and (_02611_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_02612_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_02613_, _02612_, _39078_);
  or (_39472_, _02613_, _02611_);
  and (_02614_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_02615_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_02616_, _02615_, _39078_);
  or (_39473_, _02616_, _02614_);
  and (_39474_, _01887_, _42882_);
  nor (_39475_, _01897_, rst);
  and (_39476_, _01893_, _42882_);
  and (_02617_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02618_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_02619_, _02618_, _02617_);
  and (_39477_, _02619_, _42882_);
  and (_02620_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_02621_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_02622_, _02621_, _02620_);
  and (_39478_, _02622_, _42882_);
  and (_02623_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02624_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_02625_, _02624_, _02623_);
  and (_39479_, _02625_, _42882_);
  and (_02626_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02627_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_02628_, _02627_, _02626_);
  and (_39480_, _02628_, _42882_);
  and (_02629_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02630_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_02631_, _02630_, _02629_);
  and (_39481_, _02631_, _42882_);
  and (_02632_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02633_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_02634_, _02633_, _02632_);
  and (_39483_, _02634_, _42882_);
  and (_02635_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02636_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_02637_, _02636_, _02635_);
  and (_39484_, _02637_, _42882_);
  and (_02638_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02639_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_02640_, _02639_, _02638_);
  and (_39485_, _02640_, _42882_);
  and (_02641_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_02642_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_02643_, _02642_, _02641_);
  and (_39486_, _02643_, _42882_);
  and (_02644_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_02645_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_02646_, _02645_, _02644_);
  and (_39487_, _02646_, _42882_);
  and (_02647_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_02648_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_02649_, _02648_, _02647_);
  and (_39488_, _02649_, _42882_);
  and (_02650_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_02651_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_02652_, _02651_, _02650_);
  and (_39489_, _02652_, _42882_);
  and (_02653_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_02654_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_02655_, _02654_, _02653_);
  and (_39490_, _02655_, _42882_);
  and (_02656_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_02657_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_02658_, _02657_, _02656_);
  and (_39491_, _02658_, _42882_);
  and (_02659_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_02660_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_02661_, _02660_, _02659_);
  and (_39492_, _02661_, _42882_);
  and (_02662_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_02663_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_02664_, _02663_, _02662_);
  and (_39494_, _02664_, _42882_);
  and (_02665_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_02666_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_02667_, _02666_, _02665_);
  and (_39495_, _02667_, _42882_);
  and (_02668_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_02669_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_02670_, _02669_, _02668_);
  and (_39496_, _02670_, _42882_);
  and (_02671_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_02672_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_02673_, _02672_, _02671_);
  and (_39497_, _02673_, _42882_);
  and (_02674_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_02675_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_02676_, _02675_, _02674_);
  and (_39498_, _02676_, _42882_);
  and (_02677_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_02678_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_02679_, _02678_, _02677_);
  and (_39499_, _02679_, _42882_);
  and (_02680_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_02681_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_02682_, _02681_, _02680_);
  and (_39500_, _02682_, _42882_);
  and (_02683_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_02684_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_02685_, _02684_, _02683_);
  and (_39501_, _02685_, _42882_);
  and (_02686_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_02687_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_02688_, _02687_, _02686_);
  and (_39502_, _02688_, _42882_);
  and (_02689_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_02690_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_02691_, _02690_, _02689_);
  and (_39503_, _02691_, _42882_);
  and (_02692_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_02693_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_02694_, _02693_, _02692_);
  and (_39505_, _02694_, _42882_);
  and (_02696_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_02697_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_02698_, _02697_, _02696_);
  and (_39506_, _02698_, _42882_);
  and (_02699_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_02700_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_02701_, _02700_, _02699_);
  and (_39507_, _02701_, _42882_);
  and (_02702_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_02703_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_02704_, _02703_, _02702_);
  and (_39508_, _02704_, _42882_);
  and (_02705_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_02706_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_02707_, _02706_, _02705_);
  and (_39509_, _02707_, _42882_);
  and (_02708_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_02709_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_02710_, _02709_, _02708_);
  and (_39510_, _02710_, _42882_);
  and (_02711_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02712_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_02713_, _02712_, _02711_);
  and (_39511_, _02713_, _42882_);
  and (_02714_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02715_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_02716_, _02715_, _02714_);
  and (_39512_, _02716_, _42882_);
  and (_02717_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02718_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_02719_, _02718_, _02717_);
  and (_39513_, _02719_, _42882_);
  and (_02720_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02721_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_02722_, _02721_, _02720_);
  and (_39514_, _02722_, _42882_);
  and (_02723_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02724_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_02725_, _02724_, _02723_);
  and (_39516_, _02725_, _42882_);
  and (_02726_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02727_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_02728_, _02727_, _02726_);
  and (_39517_, _02728_, _42882_);
  and (_02729_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02730_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_02731_, _02730_, _02729_);
  and (_39518_, _02731_, _42882_);
  and (_02732_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02733_, _42476_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02734_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_02735_, _02734_, _01910_);
  and (_02736_, _02735_, _02733_);
  or (_02737_, _02736_, _02732_);
  and (_39519_, _02737_, _42882_);
  and (_02738_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02739_, _42398_, _01917_);
  or (_02740_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_02741_, _02740_, _01910_);
  and (_02742_, _02741_, _02739_);
  or (_02743_, _02742_, _02738_);
  and (_39520_, _02743_, _42882_);
  and (_02744_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02745_, _42602_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02746_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_02747_, _02746_, _01910_);
  and (_02748_, _02747_, _02745_);
  or (_02749_, _02748_, _02744_);
  and (_39521_, _02749_, _42882_);
  and (_02750_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02751_, _42444_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02752_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_02753_, _02752_, _01910_);
  and (_02754_, _02753_, _02751_);
  or (_02755_, _02754_, _02750_);
  and (_39522_, _02755_, _42882_);
  and (_02756_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02757_, _42356_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02758_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_02759_, _02758_, _01910_);
  and (_02760_, _02759_, _02757_);
  or (_02761_, _02760_, _02756_);
  and (_39523_, _02761_, _42882_);
  and (_02762_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02763_, _42564_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02764_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_02765_, _02764_, _01910_);
  and (_02766_, _02765_, _02763_);
  or (_02767_, _02766_, _02762_);
  and (_39524_, _02767_, _42882_);
  and (_02768_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02769_, _42505_, _01917_);
  or (_02770_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_02771_, _02770_, _01910_);
  and (_02772_, _02771_, _02769_);
  or (_02773_, _02772_, _02768_);
  and (_39525_, _02773_, _42882_);
  and (_02774_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02775_, _42300_, _01917_);
  or (_02776_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_02777_, _02776_, _01910_);
  and (_02778_, _02777_, _02775_);
  or (_02779_, _02778_, _02774_);
  and (_39527_, _02779_, _42882_);
  and (_02780_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_02781_, _02780_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02782_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _01910_);
  and (_02783_, _02782_, _42882_);
  and (_39528_, _02783_, _02781_);
  and (_02784_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_02785_, _02784_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02786_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _01910_);
  and (_02787_, _02786_, _42882_);
  and (_39529_, _02787_, _02785_);
  and (_02788_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_02789_, _02788_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02790_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _01910_);
  and (_02791_, _02790_, _42882_);
  and (_39530_, _02791_, _02789_);
  and (_02792_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_02793_, _02792_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02794_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _01910_);
  and (_02795_, _02794_, _42882_);
  and (_39531_, _02795_, _02793_);
  and (_02797_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_02798_, _02797_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02799_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _01910_);
  and (_02800_, _02799_, _42882_);
  and (_39532_, _02800_, _02798_);
  and (_02802_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_02803_, _02802_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02804_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _01910_);
  and (_02805_, _02804_, _42882_);
  and (_39533_, _02805_, _02803_);
  and (_02807_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_02808_, _02807_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02809_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _01910_);
  and (_02810_, _02809_, _42882_);
  and (_39534_, _02810_, _02808_);
  nand (_02812_, _01924_, _31782_);
  or (_02813_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_02814_, _02813_, _42882_);
  and (_39535_, _02814_, _02812_);
  nand (_02816_, _01924_, _32458_);
  or (_02817_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_02818_, _02817_, _42882_);
  and (_39536_, _02818_, _02816_);
  nand (_02819_, _01924_, _33154_);
  or (_02821_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_02822_, _02821_, _42882_);
  and (_39538_, _02822_, _02819_);
  nand (_02823_, _01924_, _33906_);
  or (_02824_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_02826_, _02824_, _42882_);
  and (_39539_, _02826_, _02823_);
  nand (_02828_, _01924_, _34667_);
  or (_02829_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_02830_, _02829_, _42882_);
  and (_39540_, _02830_, _02828_);
  nand (_02831_, _01924_, _35461_);
  or (_02833_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_02834_, _02833_, _42882_);
  and (_39541_, _02834_, _02831_);
  nand (_02836_, _01924_, _36179_);
  or (_02837_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_02839_, _02837_, _42882_);
  and (_39542_, _02839_, _02836_);
  nand (_02840_, _01924_, _30603_);
  or (_02842_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_02843_, _02842_, _42882_);
  and (_39543_, _02843_, _02840_);
  nand (_02846_, _01924_, _38660_);
  or (_02847_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_02848_, _02847_, _42882_);
  and (_39544_, _02848_, _02846_);
  nand (_02850_, _01924_, _38693_);
  or (_02851_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_02853_, _02851_, _42882_);
  and (_39545_, _02853_, _02850_);
  nand (_02854_, _01924_, _38724_);
  or (_02856_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_02857_, _02856_, _42882_);
  and (_39546_, _02857_, _02854_);
  nand (_02859_, _01924_, _38756_);
  or (_02860_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_02861_, _02860_, _42882_);
  and (_39547_, _02861_, _02859_);
  nand (_02862_, _01924_, _38787_);
  or (_02863_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_02865_, _02863_, _42882_);
  and (_39549_, _02865_, _02862_);
  nand (_02867_, _01924_, _38821_);
  or (_02869_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_02870_, _02869_, _42882_);
  and (_39550_, _02870_, _02867_);
  not (_02872_, _01924_);
  or (_02873_, _02872_, _38847_);
  or (_02874_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_02876_, _02874_, _42882_);
  and (_39551_, _02876_, _02873_);
  nor (_39760_, _42319_, rst);
  and (_02879_, _42275_, _39022_);
  nand (_02880_, _02879_, _38485_);
  or (_02881_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_02883_, _02881_, _42882_);
  and (_39762_, _02883_, _02880_);
  and (_02884_, _42275_, _39280_);
  nand (_02886_, _02884_, _38485_);
  or (_02887_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_02889_, _02887_, _42882_);
  and (_39763_, _02889_, _02886_);
  and (_02891_, _42275_, _27045_);
  nor (_02892_, _02884_, _02891_);
  and (_02893_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_02895_, _27045_, _27714_);
  not (_02896_, _02895_);
  nor (_02897_, _02896_, _38485_);
  and (_02899_, _33329_, _27703_);
  and (_02900_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or (_02901_, _02900_, _02897_);
  and (_02903_, _02901_, _42275_);
  or (_02904_, _02903_, _02893_);
  and (_39764_, _02904_, _42882_);
  and (_02906_, _42275_, _41396_);
  nand (_02907_, _02906_, _38485_);
  or (_02908_, _02906_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_02910_, _02908_, _42882_);
  and (_39765_, _02910_, _02907_);
  nand (_02911_, _02879_, _38464_);
  or (_02913_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_02915_, _02913_, _42882_);
  and (_39792_, _02915_, _02911_);
  nand (_02917_, _02879_, _38456_);
  or (_02918_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_02920_, _02918_, _42882_);
  and (_39793_, _02920_, _02917_);
  nand (_02921_, _02879_, _38449_);
  or (_02922_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_02923_, _02922_, _42882_);
  and (_39794_, _02923_, _02921_);
  nand (_02925_, _02879_, _38442_);
  or (_02927_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_02928_, _02927_, _42882_);
  and (_39795_, _02928_, _02925_);
  nand (_02930_, _02879_, _38434_);
  or (_02931_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_02932_, _02931_, _42882_);
  and (_39796_, _02932_, _02930_);
  nand (_02934_, _02879_, _38428_);
  or (_02935_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_02938_, _02935_, _42882_);
  and (_39797_, _02938_, _02934_);
  nand (_02939_, _02879_, _38420_);
  or (_02941_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_02942_, _02941_, _42882_);
  and (_39798_, _02942_, _02939_);
  nand (_02944_, _02884_, _38464_);
  or (_02945_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_02946_, _02945_, _42882_);
  and (_39799_, _02946_, _02944_);
  nand (_02949_, _02884_, _38456_);
  or (_02951_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_02952_, _02951_, _42882_);
  and (_39800_, _02952_, _02949_);
  nand (_02953_, _02884_, _38449_);
  or (_02955_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_02956_, _02955_, _42882_);
  and (_39801_, _02956_, _02953_);
  nand (_02958_, _02884_, _38442_);
  or (_02959_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_02961_, _02959_, _42882_);
  and (_39803_, _02961_, _02958_);
  nand (_02963_, _02884_, _38434_);
  or (_02964_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_02966_, _02964_, _42882_);
  and (_39804_, _02966_, _02963_);
  nand (_02967_, _02884_, _38428_);
  or (_02969_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_02970_, _02969_, _42882_);
  and (_39805_, _02970_, _02967_);
  nand (_02973_, _02884_, _38420_);
  or (_02974_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_02975_, _02974_, _42882_);
  and (_39806_, _02975_, _02973_);
  not (_02977_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_02979_, _42275_, _02895_);
  nor (_02980_, _02979_, _02977_);
  and (_02981_, _02979_, _38465_);
  or (_02982_, _02981_, _02980_);
  and (_39807_, _02982_, _42882_);
  and (_02985_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_02986_, _02896_, _38456_);
  and (_02988_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_02989_, _02988_, _02986_);
  and (_02990_, _02989_, _42275_);
  or (_02992_, _02990_, _02985_);
  and (_39808_, _02992_, _42882_);
  and (_02993_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_02995_, _02896_, _38449_);
  and (_02996_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or (_02998_, _02996_, _02995_);
  and (_03000_, _02998_, _42275_);
  or (_03001_, _03000_, _02993_);
  and (_39809_, _03001_, _42882_);
  and (_03003_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_03004_, _02896_, _38442_);
  and (_03005_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_03007_, _03005_, _03004_);
  and (_03008_, _03007_, _42275_);
  or (_03010_, _03008_, _03003_);
  and (_39810_, _03010_, _42882_);
  and (_03012_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_03013_, _02896_, _38434_);
  and (_03015_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or (_03016_, _03015_, _03013_);
  and (_03017_, _03016_, _42275_);
  or (_03019_, _03017_, _03012_);
  and (_39811_, _03019_, _42882_);
  and (_03020_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_03022_, _02896_, _38428_);
  and (_03023_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_03024_, _03023_, _03022_);
  and (_03026_, _03024_, _42275_);
  or (_03027_, _03026_, _03020_);
  and (_39812_, _03027_, _42882_);
  and (_03029_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_03030_, _02896_, _38420_);
  and (_03031_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_03033_, _03031_, _03030_);
  and (_03034_, _03033_, _42275_);
  or (_03035_, _03034_, _03029_);
  and (_39814_, _03035_, _42882_);
  not (_03037_, _02906_);
  nor (_03039_, _03037_, _38464_);
  and (_03040_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_03041_, _03040_, _03039_);
  and (_39815_, _03041_, _42882_);
  nor (_03042_, _03037_, _38456_);
  and (_03043_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_03044_, _03043_, _03042_);
  and (_39816_, _03044_, _42882_);
  nand (_03046_, _02906_, _38449_);
  or (_03047_, _02906_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_03049_, _03047_, _42882_);
  and (_39817_, _03049_, _03046_);
  nor (_03050_, _03037_, _38442_);
  and (_03052_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_03053_, _03052_, _03050_);
  and (_39818_, _03053_, _42882_);
  nand (_03055_, _02906_, _38434_);
  or (_03056_, _02906_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_03057_, _03056_, _42882_);
  and (_39819_, _03057_, _03055_);
  nand (_03059_, _02906_, _38428_);
  or (_03060_, _02906_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_03062_, _03060_, _42882_);
  and (_39820_, _03062_, _03059_);
  nor (_03063_, _03037_, _38420_);
  and (_03065_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_03066_, _03065_, _03063_);
  and (_39821_, _03066_, _42882_);
  not (_03068_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_03069_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_03070_, _03069_, _03068_);
  and (_03072_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _42882_);
  and (_39849_, _03072_, _03070_);
  nor (_03073_, _03070_, rst);
  nand (_03075_, _03069_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03076_, _03069_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03077_, _03076_, _03075_);
  and (_39850_, _03077_, _03073_);
  nor (_03079_, _42527_, _42573_);
  not (_03080_, _42304_);
  and (_03082_, _42365_, _03080_);
  and (_03083_, _03082_, _03079_);
  and (_03084_, _03083_, _42448_);
  and (_03086_, _03084_, _39021_);
  nor (_03087_, _03086_, _01364_);
  not (_03088_, _42527_);
  and (_03090_, _03088_, _42573_);
  nor (_03091_, _42365_, _42304_);
  and (_03092_, _03091_, _42448_);
  and (_03094_, _03092_, _03090_);
  not (_03095_, _42610_);
  and (_03097_, _39113_, _39100_);
  nor (_03098_, _39113_, _39100_);
  or (_03099_, _03098_, _03097_);
  nor (_03100_, _39169_, _39125_);
  and (_03102_, _39169_, _39125_);
  nor (_03103_, _03102_, _03100_);
  nor (_03104_, _03103_, _03099_);
  and (_03106_, _03103_, _03099_);
  nor (_03107_, _03106_, _03104_);
  and (_03108_, _39193_, _39181_);
  nor (_03110_, _39193_, _39181_);
  nor (_03111_, _03110_, _03108_);
  nor (_03112_, _39204_, _39045_);
  and (_03114_, _39204_, _39045_);
  nor (_03115_, _03114_, _03112_);
  or (_03116_, _03115_, _03111_);
  nand (_03119_, _03115_, _03111_);
  and (_03120_, _03119_, _03116_);
  or (_03121_, _03120_, _03107_);
  nand (_03123_, _03120_, _03107_);
  and (_03124_, _03123_, _03121_);
  or (_03125_, _03124_, _03095_);
  and (_03127_, _42484_, _42402_);
  or (_03128_, _42610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03130_, _03128_, _03127_);
  and (_03131_, _03130_, _03125_);
  nor (_03132_, _42484_, _42402_);
  nor (_03133_, _42610_, _38889_);
  and (_03135_, _42610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_03136_, _03135_, _03133_);
  and (_03137_, _03136_, _03132_);
  or (_03139_, _42610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  not (_03140_, _42484_);
  and (_03141_, _03140_, _42402_);
  nand (_03143_, _42610_, _38905_);
  and (_03144_, _03143_, _03141_);
  and (_03145_, _03144_, _03139_);
  or (_03147_, _03145_, _03137_);
  or (_03148_, _03095_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_03149_, _03140_, _42402_);
  or (_03151_, _42610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_03152_, _03151_, _03149_);
  and (_03153_, _03152_, _03148_);
  or (_03155_, _03153_, _03147_);
  or (_03156_, _03155_, _03131_);
  and (_03157_, _03156_, _03094_);
  and (_03159_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_03160_, _03159_, _42610_);
  and (_03162_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_03163_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_03164_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_03165_, _03164_, _03163_);
  or (_03166_, _03165_, _03162_);
  or (_03168_, _03166_, _03160_);
  and (_03169_, _42527_, _42573_);
  and (_03170_, _03091_, _42449_);
  and (_03172_, _03170_, _03169_);
  and (_03173_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03174_, _03173_, _03095_);
  and (_03176_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_03177_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_03178_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_03180_, _03178_, _03177_);
  or (_03181_, _03180_, _03176_);
  or (_03182_, _03181_, _03174_);
  and (_03184_, _03182_, _03172_);
  and (_03185_, _03184_, _03168_);
  and (_03186_, _38244_, _38271_);
  nor (_03188_, _03186_, _38369_);
  not (_03189_, _38288_);
  and (_03190_, _00836_, _03189_);
  and (_03192_, _03190_, _03188_);
  and (_03193_, _38265_, _38260_);
  or (_03195_, _00921_, _00768_);
  or (_03196_, _03195_, _00834_);
  or (_03197_, _03196_, _38300_);
  or (_03198_, _03197_, _00766_);
  nor (_03200_, _03198_, _03193_);
  and (_03201_, _03200_, _38324_);
  and (_03202_, _03201_, _03192_);
  and (_03204_, _03202_, _01110_);
  nor (_03205_, _03204_, _36407_);
  or (_03206_, _03205_, p3_in[0]);
  not (_03208_, _03205_);
  or (_03209_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_03210_, _03209_, _03206_);
  and (_03212_, _03210_, _03127_);
  or (_03213_, _03212_, _03095_);
  or (_03214_, _03205_, p3_in[3]);
  or (_03216_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03217_, _03216_, _03214_);
  and (_03218_, _03217_, _03132_);
  or (_03220_, _03205_, p3_in[2]);
  or (_03221_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03222_, _03221_, _03220_);
  and (_03224_, _03222_, _03149_);
  or (_03225_, _03205_, p3_in[1]);
  or (_03227_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03228_, _03227_, _03225_);
  and (_03229_, _03228_, _03141_);
  or (_03230_, _03229_, _03224_);
  or (_03232_, _03230_, _03218_);
  or (_03233_, _03232_, _03213_);
  and (_03234_, _03092_, _42574_);
  and (_03236_, _03234_, _42527_);
  or (_03237_, _03205_, p3_in[4]);
  or (_03238_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_03240_, _03238_, _03237_);
  and (_03241_, _03240_, _03127_);
  or (_03242_, _03241_, _42610_);
  or (_03244_, _03205_, p3_in[7]);
  or (_03245_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_03246_, _03245_, _03244_);
  and (_03248_, _03246_, _03132_);
  or (_03249_, _03205_, p3_in[6]);
  or (_03250_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03252_, _03250_, _03249_);
  and (_03253_, _03252_, _03149_);
  or (_03254_, _03205_, p3_in[5]);
  or (_03256_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03257_, _03256_, _03254_);
  and (_03259_, _03257_, _03141_);
  or (_03260_, _03259_, _03253_);
  or (_03261_, _03260_, _03248_);
  or (_03262_, _03261_, _03242_);
  and (_03264_, _03262_, _03236_);
  and (_03265_, _03264_, _03233_);
  or (_03266_, _03265_, _03185_);
  or (_03268_, _03205_, p0_in[1]);
  or (_03269_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03270_, _03269_, _03268_);
  and (_03272_, _03270_, _03141_);
  or (_03273_, _03272_, _03095_);
  or (_03274_, _03205_, p0_in[3]);
  or (_03276_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03277_, _03276_, _03274_);
  and (_03278_, _03277_, _03132_);
  or (_03280_, _03205_, p0_in[0]);
  or (_03281_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_03282_, _03281_, _03280_);
  and (_03284_, _03282_, _03127_);
  or (_03285_, _03205_, p0_in[2]);
  or (_03286_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_03288_, _03286_, _03285_);
  and (_03289_, _03288_, _03149_);
  or (_03290_, _03289_, _03284_);
  or (_03291_, _03290_, _03278_);
  or (_03292_, _03291_, _03273_);
  and (_03293_, _03169_, _03082_);
  and (_03294_, _03293_, _42448_);
  or (_03295_, _03205_, p0_in[5]);
  or (_03296_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03297_, _03296_, _03295_);
  and (_03298_, _03297_, _03141_);
  or (_03299_, _03298_, _42610_);
  or (_03300_, _03205_, p0_in[7]);
  or (_03301_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03302_, _03301_, _03300_);
  and (_03303_, _03302_, _03132_);
  or (_03304_, _03205_, p0_in[4]);
  or (_03305_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_03306_, _03305_, _03304_);
  and (_03307_, _03306_, _03127_);
  or (_03308_, _03205_, p0_in[6]);
  or (_03309_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03310_, _03309_, _03308_);
  and (_03311_, _03310_, _03149_);
  or (_03312_, _03311_, _03307_);
  or (_03313_, _03312_, _03303_);
  or (_03314_, _03313_, _03299_);
  and (_03315_, _03314_, _03294_);
  and (_03316_, _03315_, _03292_);
  and (_03317_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_03318_, _03317_, _03095_);
  and (_03319_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_03320_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_03321_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03322_, _03321_, _03320_);
  or (_03323_, _03322_, _03319_);
  or (_03324_, _03323_, _03318_);
  and (_03325_, _42527_, _42574_);
  and (_03326_, _03325_, _03170_);
  and (_03327_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_03328_, _03327_, _42610_);
  and (_03329_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_03330_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03331_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_03332_, _03331_, _03330_);
  or (_03333_, _03332_, _03329_);
  or (_03334_, _03333_, _03328_);
  and (_03335_, _03334_, _03326_);
  and (_03336_, _03335_, _03324_);
  or (_03337_, _03336_, _03316_);
  or (_03338_, _03337_, _03266_);
  and (_03339_, _01379_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_03340_, _03205_, p2_in[1]);
  or (_03341_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_03342_, _03341_, _03340_);
  and (_03343_, _03342_, _03141_);
  or (_03344_, _03343_, _03095_);
  or (_03345_, _03205_, p2_in[3]);
  or (_03346_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03347_, _03346_, _03345_);
  and (_03348_, _03347_, _03132_);
  or (_03349_, _03205_, p2_in[0]);
  or (_03350_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_03351_, _03350_, _03349_);
  and (_03352_, _03351_, _03127_);
  or (_03353_, _03205_, p2_in[2]);
  or (_03354_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03355_, _03354_, _03353_);
  and (_03356_, _03355_, _03149_);
  or (_03357_, _03356_, _03352_);
  or (_03358_, _03357_, _03348_);
  or (_03359_, _03358_, _03344_);
  and (_03360_, _03325_, _03082_);
  and (_03362_, _03360_, _42448_);
  or (_03363_, _03205_, p2_in[5]);
  or (_03364_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03365_, _03364_, _03363_);
  and (_03366_, _03365_, _03141_);
  or (_03367_, _03366_, _42610_);
  or (_03368_, _03205_, p2_in[7]);
  or (_03369_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_03370_, _03369_, _03368_);
  and (_03371_, _03370_, _03132_);
  or (_03372_, _03205_, p2_in[4]);
  or (_03373_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_03374_, _03373_, _03372_);
  and (_03375_, _03374_, _03127_);
  or (_03376_, _03205_, p2_in[6]);
  or (_03377_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03378_, _03377_, _03376_);
  and (_03379_, _03378_, _03149_);
  or (_03380_, _03379_, _03375_);
  or (_03381_, _03380_, _03371_);
  or (_03382_, _03381_, _03367_);
  and (_03383_, _03382_, _03362_);
  and (_03384_, _03383_, _03359_);
  or (_03385_, _03384_, _03339_);
  and (_03386_, _42527_, _03080_);
  nand (_03387_, _03386_, _42449_);
  nor (_03388_, _03092_, _28613_);
  and (_03389_, _03388_, _03387_);
  nor (_03390_, _03362_, _03084_);
  and (_03391_, _03090_, _03082_);
  and (_03392_, _03391_, _42449_);
  nor (_03393_, _03392_, _03294_);
  and (_03394_, _03393_, _03390_);
  and (_03395_, _03394_, _03389_);
  and (_03396_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_03397_, _03396_, _42610_);
  and (_03398_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03399_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03400_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_03401_, _03400_, _03399_);
  or (_03402_, _03401_, _03398_);
  or (_03403_, _03402_, _03397_);
  and (_03404_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03405_, _03404_, _03095_);
  and (_03406_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_03407_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_03408_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03409_, _03408_, _03407_);
  or (_03410_, _03409_, _03406_);
  or (_03411_, _03410_, _03405_);
  and (_03412_, _03411_, _03084_);
  and (_03413_, _03412_, _03403_);
  or (_03414_, _03413_, _03395_);
  or (_03415_, _03414_, _03385_);
  or (_03416_, _03415_, _03338_);
  and (_03417_, _03082_, _42449_);
  and (_03418_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_03419_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_03420_, _03419_, _03418_);
  and (_03421_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_03422_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_03423_, _03422_, _03421_);
  or (_03424_, _03423_, _03420_);
  and (_03425_, _03424_, _42610_);
  and (_03426_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03427_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_03428_, _03427_, _03426_);
  and (_03429_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_03430_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_03431_, _03430_, _03429_);
  or (_03432_, _03431_, _03428_);
  and (_03433_, _03432_, _03095_);
  or (_03434_, _03433_, _03425_);
  and (_03435_, _03434_, _03325_);
  and (_03436_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03437_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_03438_, _03437_, _03436_);
  and (_03439_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_03440_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03441_, _03440_, _03439_);
  or (_03442_, _03441_, _03438_);
  and (_03443_, _03442_, _03095_);
  and (_03444_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_03445_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_03446_, _03445_, _03444_);
  and (_03447_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_03448_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_03449_, _03448_, _03447_);
  or (_03450_, _03449_, _03446_);
  and (_03451_, _03450_, _42610_);
  or (_03452_, _03451_, _03443_);
  and (_03453_, _03452_, _03169_);
  or (_03454_, _03453_, _03435_);
  and (_03455_, _03454_, _03417_);
  or (_03456_, _03205_, p1_in[4]);
  or (_03457_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03458_, _03457_, _03456_);
  and (_03459_, _03458_, _03127_);
  or (_03460_, _03459_, _42610_);
  or (_03461_, _03205_, p1_in[7]);
  or (_03462_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_03463_, _03462_, _03461_);
  and (_03464_, _03463_, _03132_);
  or (_03465_, _03205_, p1_in[6]);
  or (_03466_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03467_, _03466_, _03465_);
  and (_03468_, _03467_, _03149_);
  or (_03469_, _03205_, p1_in[5]);
  or (_03470_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03471_, _03470_, _03469_);
  and (_03472_, _03471_, _03141_);
  or (_03473_, _03472_, _03468_);
  or (_03474_, _03473_, _03464_);
  or (_03475_, _03474_, _03460_);
  and (_03476_, _03169_, _03092_);
  or (_03477_, _03205_, p1_in[0]);
  or (_03478_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_03479_, _03478_, _03477_);
  and (_03480_, _03479_, _03127_);
  or (_03481_, _03480_, _03095_);
  or (_03482_, _03205_, p1_in[3]);
  or (_03483_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03484_, _03483_, _03482_);
  and (_03485_, _03484_, _03132_);
  or (_03486_, _03205_, p1_in[2]);
  or (_03487_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03488_, _03487_, _03486_);
  and (_03489_, _03488_, _03149_);
  or (_03490_, _03205_, p1_in[1]);
  or (_03491_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03492_, _03491_, _03490_);
  and (_03493_, _03492_, _03141_);
  or (_03494_, _03493_, _03489_);
  or (_03495_, _03494_, _03485_);
  or (_03496_, _03495_, _03481_);
  and (_03497_, _03496_, _03476_);
  and (_03498_, _03497_, _03475_);
  and (_03499_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_03500_, _03499_, _42610_);
  and (_03501_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03502_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_03503_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_03504_, _03503_, _03502_);
  or (_03505_, _03504_, _03501_);
  or (_03506_, _03505_, _03500_);
  and (_03507_, _03234_, _03088_);
  and (_03508_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_03509_, _03508_, _03095_);
  and (_03510_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_03511_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_03512_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_03513_, _03512_, _03511_);
  or (_03514_, _03513_, _03510_);
  or (_03515_, _03514_, _03509_);
  and (_03516_, _03515_, _03507_);
  and (_03517_, _03516_, _03506_);
  and (_03518_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03519_, _03518_, _03095_);
  and (_03520_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_03521_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_03522_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03523_, _03522_, _03521_);
  or (_03524_, _03523_, _03520_);
  or (_03525_, _03524_, _03519_);
  and (_03526_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_03527_, _03526_, _42610_);
  and (_03528_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03529_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03530_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_03531_, _03530_, _03529_);
  or (_03532_, _03531_, _03528_);
  or (_03533_, _03532_, _03527_);
  and (_03534_, _03533_, _03392_);
  and (_03535_, _03534_, _03525_);
  or (_03536_, _03535_, _03517_);
  or (_03537_, _03536_, _03498_);
  or (_03538_, _03537_, _03455_);
  or (_03539_, _03538_, _03416_);
  or (_03540_, _03539_, _03157_);
  nand (_03541_, _03339_, _31282_);
  nand (_03542_, _03541_, _03540_);
  nand (_03543_, _03542_, _03087_);
  nand (_03544_, _42610_, _38456_);
  nand (_03545_, _03095_, _38428_);
  and (_03546_, _03545_, _03141_);
  and (_03547_, _03546_, _03544_);
  and (_03548_, _42610_, _42600_);
  nor (_03549_, _42610_, _38420_);
  or (_03550_, _03549_, _03548_);
  and (_03551_, _03550_, _03149_);
  nor (_03552_, _42610_, _38434_);
  and (_03553_, _42610_, _38465_);
  or (_03554_, _03553_, _03552_);
  and (_03555_, _03554_, _03127_);
  nand (_03556_, _42610_, _38442_);
  nand (_03557_, _03095_, _38485_);
  and (_03558_, _03557_, _03132_);
  and (_03559_, _03558_, _03556_);
  or (_03560_, _03559_, _03555_);
  or (_03561_, _03560_, _03551_);
  or (_03563_, _03561_, _03547_);
  or (_03564_, _03563_, _03087_);
  and (_03565_, _03564_, _42882_);
  and (_39851_, _03565_, _03543_);
  nor (_03566_, _42365_, _42574_);
  nor (_03567_, _42527_, _42304_);
  and (_03568_, _42448_, _42610_);
  and (_03569_, _03568_, _03127_);
  and (_03570_, _03569_, _03567_);
  and (_03571_, _03570_, _03566_);
  and (_03572_, _03571_, _01438_);
  and (_03573_, _03569_, _03083_);
  and (_03574_, _03573_, _39018_);
  nor (_03575_, _03574_, _03572_);
  and (_03576_, _03568_, _03132_);
  and (_03577_, _03576_, _03293_);
  nand (_03578_, _03577_, _38533_);
  and (_03579_, _03578_, _03575_);
  nor (_03580_, _03579_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_03581_, _03580_);
  not (_03582_, _39031_);
  and (_03583_, _03132_, _03095_);
  nor (_03584_, _03583_, _03582_);
  and (_03585_, _03584_, _01362_);
  and (_03586_, _03573_, _39021_);
  nor (_03587_, _03586_, _03585_);
  and (_03588_, _03587_, _01382_);
  and (_03589_, _03588_, _03581_);
  and (_03590_, _03293_, _03149_);
  and (_03591_, _03590_, _03568_);
  and (_03592_, _03591_, _38533_);
  or (_03593_, _03592_, rst);
  nor (_39853_, _03593_, _03589_);
  nand (_03594_, _03592_, _30603_);
  and (_03595_, _42449_, _42610_);
  and (_03596_, _03595_, _03127_);
  and (_03597_, _03596_, _03391_);
  and (_03598_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_03599_, _42448_, _42610_);
  and (_03600_, _03599_, _03127_);
  and (_03601_, _03600_, _03391_);
  and (_03602_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_03603_, _03602_, _03598_);
  and (_03604_, _03595_, _03149_);
  and (_03605_, _03604_, _03391_);
  and (_03606_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_03607_, _03599_, _03141_);
  and (_03608_, _03607_, _03391_);
  and (_03609_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_03610_, _03609_, _03606_);
  or (_03611_, _03610_, _03603_);
  and (_03612_, _03596_, _03293_);
  and (_03613_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03614_, _03595_, _03132_);
  and (_03615_, _03614_, _03391_);
  and (_03616_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_03617_, _03616_, _03613_);
  and (_03618_, _03596_, _03360_);
  and (_03619_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03620_, _03583_, _42448_);
  nor (_03621_, _42365_, _42573_);
  and (_03622_, _03621_, _03386_);
  and (_03623_, _03622_, _03620_);
  and (_03624_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_03625_, _03624_, _03619_);
  or (_03626_, _03625_, _03617_);
  or (_03627_, _03626_, _03611_);
  and (_03628_, _03614_, _03293_);
  and (_03629_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_03630_, _03595_, _03141_);
  and (_03631_, _03630_, _03293_);
  and (_03632_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_03633_, _03632_, _03629_);
  and (_03634_, _03607_, _03293_);
  and (_03635_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_03636_, _03604_, _03293_);
  and (_03637_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_03638_, _03637_, _03635_);
  or (_03639_, _03638_, _03633_);
  and (_03640_, _03169_, _03091_);
  and (_03641_, _03640_, _03630_);
  and (_03642_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_03643_, _03596_, _03640_);
  and (_03644_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_03645_, _03644_, _03642_);
  and (_03646_, _03600_, _03293_);
  and (_03647_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_03648_, _03583_, _03294_);
  and (_03649_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_03650_, _03649_, _03647_);
  or (_03651_, _03650_, _03645_);
  or (_03652_, _03651_, _03639_);
  or (_03653_, _03652_, _03627_);
  and (_03654_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_03655_, _03293_, _03132_);
  and (_03656_, _03655_, _03568_);
  and (_03657_, _03656_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_03658_, _03657_, _03654_);
  and (_03659_, _03621_, _03570_);
  and (_03660_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03661_, _03293_, _03141_);
  and (_03662_, _03661_, _03568_);
  and (_03663_, _03662_, _42245_);
  or (_03664_, _03663_, _03660_);
  or (_03665_, _03664_, _03658_);
  and (_03666_, _03569_, _03360_);
  and (_03667_, _03666_, _03370_);
  and (_03668_, _03622_, _03569_);
  and (_03669_, _03668_, _03246_);
  or (_03670_, _03669_, _03667_);
  and (_03671_, _03569_, _03293_);
  and (_03672_, _03671_, _03302_);
  and (_03673_, _03640_, _03569_);
  and (_03674_, _03673_, _03463_);
  or (_03675_, _03674_, _03672_);
  or (_03676_, _03675_, _03670_);
  or (_03677_, _03676_, _03665_);
  and (_03678_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_03679_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03680_, _03679_, _03678_);
  or (_03681_, _03680_, _03677_);
  or (_03682_, _03681_, _03653_);
  and (_03683_, _03682_, _03589_);
  and (_03684_, _03569_, _03386_);
  or (_03685_, _03659_, _03684_);
  or (_03686_, _03685_, _03662_);
  and (_03687_, _03595_, _03655_);
  or (_03688_, _03646_, _03641_);
  or (_03689_, _03634_, _03643_);
  or (_03690_, _03689_, _03688_);
  or (_03691_, _03690_, _03687_);
  or (_03692_, _03691_, _03686_);
  or (_03693_, _03623_, _03573_);
  or (_03694_, _03648_, _03571_);
  or (_03695_, _03694_, _03693_);
  or (_03696_, _03615_, _03605_);
  or (_03697_, _03608_, _03612_);
  or (_03698_, _03697_, _03696_);
  or (_03699_, _03698_, _03656_);
  or (_03700_, _03699_, _03695_);
  and (_03701_, _03595_, _03590_);
  or (_03702_, _03631_, _03618_);
  or (_03703_, _03702_, _03701_);
  and (_03704_, _03392_, _03127_);
  or (_03705_, _03704_, _03591_);
  or (_03706_, _03705_, _03703_);
  or (_03707_, _03706_, _03700_);
  or (_03708_, _03707_, _03692_);
  nand (_03709_, _03708_, _03589_);
  and (_03710_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_03711_, _03710_, _03683_);
  or (_03712_, _03711_, _03592_);
  and (_03713_, _03712_, _42882_);
  and (_39854_, _03713_, _03594_);
  nor (_39935_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_03714_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_03715_, _03069_, rst);
  and (_39936_, _03715_, _03714_);
  nor (_03716_, _03069_, _03068_);
  or (_03717_, _03716_, _03070_);
  and (_03718_, _03075_, _42882_);
  and (_39937_, _03718_, _03717_);
  and (_03719_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_03720_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_03721_, _03720_, _03719_);
  and (_03722_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_03723_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_03724_, _03723_, _03722_);
  or (_03725_, _03724_, _03721_);
  and (_03726_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_03727_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_03728_, _03727_, _03726_);
  and (_03729_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_03730_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_03731_, _03730_, _03729_);
  or (_03732_, _03731_, _03728_);
  or (_03733_, _03732_, _03725_);
  and (_03734_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_03735_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_03736_, _03735_, _03734_);
  and (_03737_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_03738_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or (_03739_, _03738_, _03737_);
  or (_03740_, _03739_, _03736_);
  and (_03741_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_03742_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_03743_, _03742_, _03741_);
  and (_03744_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_03745_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  or (_03746_, _03745_, _03744_);
  or (_03747_, _03746_, _03743_);
  or (_03748_, _03747_, _03740_);
  or (_03749_, _03748_, _03733_);
  and (_03750_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_03751_, _03662_, _42480_);
  or (_03752_, _03751_, _03750_);
  and (_03753_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_03754_, _03577_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_03755_, _03754_, _03753_);
  or (_03756_, _03755_, _03752_);
  and (_03758_, _03666_, _03351_);
  and (_03759_, _03668_, _03210_);
  or (_03760_, _03759_, _03758_);
  and (_03761_, _03671_, _03282_);
  and (_03762_, _03673_, _03479_);
  or (_03763_, _03762_, _03761_);
  or (_03764_, _03763_, _03760_);
  or (_03765_, _03764_, _03756_);
  and (_03766_, _03571_, _03124_);
  and (_03767_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03768_, _03767_, _03766_);
  or (_03769_, _03768_, _03765_);
  or (_03770_, _03769_, _03749_);
  and (_03771_, _03770_, _03589_);
  and (_03772_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or (_03773_, _03772_, _03592_);
  or (_03774_, _03773_, _03771_);
  nand (_03775_, _03592_, _31782_);
  and (_03776_, _03775_, _42882_);
  and (_39938_, _03776_, _03774_);
  and (_03777_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_03778_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_03779_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_03780_, _03779_, _03778_);
  and (_03781_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_03782_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_03783_, _03782_, _03781_);
  or (_03784_, _03783_, _03780_);
  and (_03785_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_03786_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_03787_, _03786_, _03785_);
  and (_03788_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_03789_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_03790_, _03789_, _03788_);
  or (_03791_, _03790_, _03787_);
  or (_03792_, _03791_, _03784_);
  and (_03793_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_03794_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_03795_, _03794_, _03793_);
  and (_03796_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_03797_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_03798_, _03797_, _03796_);
  or (_03799_, _03798_, _03795_);
  and (_03800_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_03801_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03802_, _03801_, _03800_);
  and (_03803_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_03804_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_03805_, _03804_, _03803_);
  or (_03806_, _03805_, _03802_);
  or (_03807_, _03806_, _03799_);
  or (_03808_, _03807_, _03792_);
  and (_03809_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_03810_, _03662_, _42387_);
  or (_03811_, _03810_, _03809_);
  and (_03812_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_03813_, _03577_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_03814_, _03813_, _03812_);
  or (_03815_, _03814_, _03811_);
  and (_03816_, _03666_, _03342_);
  and (_03817_, _03668_, _03228_);
  or (_03818_, _03817_, _03816_);
  and (_03819_, _03671_, _03270_);
  and (_03820_, _03673_, _03492_);
  or (_03821_, _03820_, _03819_);
  or (_03822_, _03821_, _03818_);
  or (_03823_, _03822_, _03815_);
  and (_03824_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03825_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03826_, _03825_, _03824_);
  or (_03827_, _03826_, _03823_);
  or (_03828_, _03827_, _03808_);
  and (_03829_, _03828_, _03589_);
  or (_03830_, _03829_, _03592_);
  or (_03831_, _03830_, _03777_);
  nand (_03832_, _03592_, _32458_);
  and (_03833_, _03832_, _42882_);
  and (_39939_, _03833_, _03831_);
  and (_03834_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_03835_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_03836_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_03837_, _03836_, _03835_);
  and (_03838_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_03839_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_03840_, _03839_, _03838_);
  or (_03841_, _03840_, _03837_);
  and (_03842_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_03843_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_03844_, _03843_, _03842_);
  and (_03845_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_03846_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03847_, _03846_, _03845_);
  or (_03848_, _03847_, _03844_);
  or (_03849_, _03848_, _03841_);
  and (_03850_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_03851_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_03852_, _03851_, _03850_);
  and (_03853_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_03854_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_03855_, _03854_, _03853_);
  or (_03856_, _03855_, _03852_);
  and (_03857_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_03858_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_03859_, _03858_, _03857_);
  and (_03860_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_03861_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_03862_, _03861_, _03860_);
  or (_03863_, _03862_, _03859_);
  or (_03864_, _03863_, _03856_);
  or (_03865_, _03864_, _03849_);
  and (_03866_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_03867_, _03656_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_03868_, _03867_, _03866_);
  and (_03869_, _03662_, _42606_);
  and (_03870_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_03871_, _03870_, _03869_);
  or (_03872_, _03871_, _03868_);
  and (_03873_, _03666_, _03355_);
  and (_03874_, _03668_, _03222_);
  or (_03875_, _03874_, _03873_);
  and (_03876_, _03671_, _03288_);
  and (_03877_, _03673_, _03488_);
  or (_03878_, _03877_, _03876_);
  or (_03879_, _03878_, _03875_);
  or (_03880_, _03879_, _03872_);
  and (_03881_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_03882_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03883_, _03882_, _03881_);
  or (_03884_, _03883_, _03880_);
  or (_03885_, _03884_, _03865_);
  and (_03886_, _03885_, _03589_);
  or (_03887_, _03886_, _03592_);
  or (_03888_, _03887_, _03834_);
  nand (_03889_, _03592_, _33154_);
  and (_03890_, _03889_, _42882_);
  and (_39940_, _03890_, _03888_);
  nand (_03891_, _03592_, _33906_);
  and (_03892_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_03893_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_03894_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_03895_, _03894_, _03893_);
  and (_03896_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_03897_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_03898_, _03897_, _03896_);
  or (_03899_, _03898_, _03895_);
  and (_03900_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_03901_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_03902_, _03901_, _03900_);
  and (_03903_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03904_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03905_, _03904_, _03903_);
  or (_03906_, _03905_, _03902_);
  or (_03907_, _03906_, _03899_);
  and (_03908_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_03909_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or (_03910_, _03909_, _03908_);
  and (_03911_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_03912_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_03913_, _03912_, _03911_);
  or (_03914_, _03913_, _03910_);
  and (_03915_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_03916_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_03917_, _03916_, _03915_);
  and (_03918_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_03919_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or (_03920_, _03919_, _03918_);
  or (_03921_, _03920_, _03917_);
  or (_03922_, _03921_, _03914_);
  or (_03923_, _03922_, _03907_);
  and (_03924_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_03925_, _03656_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_03926_, _03925_, _03924_);
  and (_03927_, _03662_, _42433_);
  and (_03928_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_03929_, _03928_, _03927_);
  or (_03930_, _03929_, _03926_);
  and (_03931_, _03666_, _03347_);
  and (_03932_, _03668_, _03217_);
  or (_03933_, _03932_, _03931_);
  and (_03934_, _03671_, _03277_);
  and (_03935_, _03673_, _03484_);
  or (_03936_, _03935_, _03934_);
  or (_03937_, _03936_, _03933_);
  or (_03938_, _03937_, _03930_);
  and (_03939_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_03940_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_03941_, _03940_, _03939_);
  or (_03942_, _03941_, _03938_);
  or (_03943_, _03942_, _03923_);
  and (_03944_, _03943_, _03589_);
  or (_03945_, _03944_, _03892_);
  or (_03946_, _03945_, _03592_);
  and (_03947_, _03946_, _42882_);
  and (_39941_, _03947_, _03891_);
  nand (_03948_, _03592_, _34667_);
  and (_03949_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_03950_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03951_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_03952_, _03951_, _03950_);
  and (_03953_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_03955_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_03956_, _03955_, _03953_);
  or (_03957_, _03956_, _03952_);
  and (_03958_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_03959_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_03960_, _03959_, _03958_);
  and (_03961_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_03962_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_03963_, _03962_, _03961_);
  or (_03964_, _03963_, _03960_);
  or (_03965_, _03964_, _03957_);
  and (_03966_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_03967_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or (_03968_, _03967_, _03966_);
  and (_03969_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_03970_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_03971_, _03970_, _03969_);
  or (_03972_, _03971_, _03968_);
  and (_03973_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_03974_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_03975_, _03974_, _03973_);
  and (_03976_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_03977_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_03978_, _03977_, _03976_);
  or (_03979_, _03978_, _03975_);
  or (_03980_, _03979_, _03972_);
  or (_03981_, _03980_, _03965_);
  and (_03982_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_03983_, _03662_, _42360_);
  or (_03984_, _03983_, _03982_);
  and (_03985_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_03986_, _03577_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_03987_, _03986_, _03985_);
  or (_03988_, _03987_, _03984_);
  and (_03989_, _03666_, _03374_);
  and (_03990_, _03668_, _03240_);
  or (_03991_, _03990_, _03989_);
  and (_03992_, _03671_, _03306_);
  and (_03993_, _03673_, _03458_);
  or (_03994_, _03993_, _03992_);
  or (_03995_, _03994_, _03991_);
  or (_03996_, _03995_, _03988_);
  and (_03997_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_03998_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_03999_, _03998_, _03997_);
  or (_04000_, _03999_, _03996_);
  or (_04001_, _04000_, _03981_);
  and (_04002_, _04001_, _03589_);
  or (_04003_, _04002_, _03949_);
  or (_04004_, _04003_, _03592_);
  and (_04005_, _04004_, _42882_);
  and (_39943_, _04005_, _03948_);
  nand (_04006_, _03592_, _35461_);
  and (_04007_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_04008_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04009_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_04010_, _04009_, _04008_);
  and (_04011_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_04012_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_04013_, _04012_, _04011_);
  or (_04014_, _04013_, _04010_);
  and (_04015_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04016_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_04017_, _04016_, _04015_);
  and (_04018_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_04019_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_04020_, _04019_, _04018_);
  or (_04021_, _04020_, _04017_);
  or (_04022_, _04021_, _04014_);
  and (_04023_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_04024_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_04025_, _04024_, _04023_);
  and (_04026_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_04027_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_04028_, _04027_, _04026_);
  or (_04029_, _04028_, _04025_);
  and (_04030_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_04031_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_04032_, _04031_, _04030_);
  and (_04033_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_04034_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_04035_, _04034_, _04033_);
  or (_04036_, _04035_, _04032_);
  or (_04037_, _04036_, _04029_);
  or (_04038_, _04037_, _04022_);
  not (_04039_, _38525_);
  and (_04040_, _03662_, _04039_);
  and (_04041_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_04042_, _04041_, _04040_);
  and (_04043_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_04044_, _03577_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_04045_, _04044_, _04043_);
  or (_04046_, _04045_, _04042_);
  and (_04047_, _03666_, _03365_);
  and (_04048_, _03668_, _03257_);
  or (_04049_, _04048_, _04047_);
  and (_04050_, _03671_, _03297_);
  and (_04051_, _03673_, _03471_);
  or (_04052_, _04051_, _04050_);
  or (_04053_, _04052_, _04049_);
  or (_04055_, _04053_, _04046_);
  and (_04056_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_04057_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_04058_, _04057_, _04056_);
  or (_04059_, _04058_, _04055_);
  or (_04060_, _04059_, _04038_);
  and (_04061_, _04060_, _03589_);
  or (_04062_, _04061_, _04007_);
  or (_04063_, _04062_, _03592_);
  and (_04064_, _04063_, _42882_);
  and (_39944_, _04064_, _04006_);
  and (_04065_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_04066_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_04067_, _04066_, _04065_);
  and (_04068_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_04069_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_04070_, _04069_, _04068_);
  or (_04071_, _04070_, _04067_);
  and (_04072_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_04073_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_04074_, _04073_, _04072_);
  and (_04075_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_04076_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_04077_, _04076_, _04075_);
  or (_04078_, _04077_, _04074_);
  or (_04079_, _04078_, _04071_);
  and (_04080_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_04081_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_04082_, _04081_, _04080_);
  and (_04083_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_04084_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_04085_, _04084_, _04083_);
  or (_04086_, _04085_, _04082_);
  and (_04087_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_04088_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_04089_, _04088_, _04087_);
  and (_04090_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_04091_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_04092_, _04091_, _04090_);
  or (_04093_, _04092_, _04089_);
  or (_04094_, _04093_, _04086_);
  or (_04095_, _04094_, _04079_);
  and (_04096_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_04097_, _03656_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_04098_, _04097_, _04096_);
  and (_04099_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_04100_, _03662_, _42508_);
  or (_04101_, _04100_, _04099_);
  or (_04102_, _04101_, _04098_);
  and (_04103_, _03666_, _03378_);
  and (_04104_, _03668_, _03252_);
  or (_04105_, _04104_, _04103_);
  and (_04106_, _03671_, _03310_);
  and (_04107_, _03673_, _03467_);
  or (_04108_, _04107_, _04106_);
  or (_04109_, _04108_, _04105_);
  or (_04110_, _04109_, _04102_);
  and (_04111_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_04112_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_04113_, _04112_, _04111_);
  or (_04114_, _04113_, _04110_);
  or (_04115_, _04114_, _04095_);
  and (_04116_, _04115_, _03589_);
  and (_04117_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or (_04118_, _04117_, _04116_);
  or (_04119_, _04118_, _03592_);
  nand (_04120_, _03592_, _36179_);
  and (_04121_, _04120_, _42882_);
  and (_39945_, _04121_, _04119_);
  and (_40015_, _42648_, _42882_);
  nor (_40019_, _42610_, rst);
  and (_40041_, _42794_, _42882_);
  nor (_40044_, _42484_, rst);
  nor (_40045_, _42402_, rst);
  not (_04122_, _00317_);
  nor (_04123_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_04124_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04125_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _04124_);
  nor (_04126_, _04125_, _04123_);
  nor (_04127_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04128_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _04124_);
  nor (_04129_, _04128_, _04127_);
  nor (_04130_, _04129_, _04126_);
  and (_04131_, _04129_, _04126_);
  nor (_04132_, _02202_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04133_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _04124_);
  nor (_04134_, _04133_, _04132_);
  and (_04135_, _04134_, _04131_);
  nor (_04136_, _04134_, _04131_);
  nor (_04137_, _04136_, _04135_);
  not (_04138_, _04137_);
  nor (_04139_, _02221_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04140_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _04124_);
  nor (_04141_, _04140_, _04139_);
  and (_04142_, _04141_, _04135_);
  nor (_04143_, _04141_, _04135_);
  nor (_04144_, _04143_, _04142_);
  and (_04145_, _04144_, _04138_);
  and (_04146_, _04145_, _04130_);
  and (_04148_, _04146_, _04122_);
  not (_04149_, _00358_);
  not (_04150_, _04129_);
  and (_04151_, _04150_, _04126_);
  and (_04152_, _04145_, _04151_);
  and (_04153_, _04152_, _04149_);
  or (_04154_, _04153_, _04148_);
  not (_04155_, _00399_);
  nor (_04156_, _04150_, _04126_);
  and (_04157_, _04145_, _04156_);
  and (_04158_, _04157_, _04155_);
  not (_04159_, _00040_);
  nor (_04160_, _04144_, _04137_);
  and (_04161_, _04160_, _04156_);
  and (_04162_, _04161_, _04159_);
  or (_04163_, _04162_, _04158_);
  or (_04164_, _04163_, _04154_);
  not (_04165_, _43768_);
  and (_04166_, _04160_, _04130_);
  and (_04167_, _04166_, _04165_);
  not (_04168_, _43809_);
  and (_04169_, _04160_, _04151_);
  and (_04170_, _04169_, _04168_);
  or (_04171_, _04170_, _04167_);
  not (_04172_, _00481_);
  and (_04173_, _04141_, _04137_);
  and (_04174_, _04173_, _04130_);
  and (_04175_, _04174_, _04172_);
  not (_04176_, _00522_);
  and (_04177_, _04173_, _04151_);
  and (_04178_, _04177_, _04176_);
  or (_04179_, _04178_, _04175_);
  not (_04180_, _00122_);
  not (_04181_, _04141_);
  and (_04182_, _04181_, _04137_);
  and (_04183_, _04182_, _04130_);
  and (_04184_, _04183_, _04180_);
  not (_04185_, _00194_);
  and (_04186_, _04182_, _04151_);
  and (_04187_, _04186_, _04185_);
  or (_04188_, _04187_, _04184_);
  or (_04189_, _04188_, _04179_);
  not (_04190_, _00081_);
  and (_04191_, _04143_, _04131_);
  and (_04192_, _04191_, _04190_);
  not (_04193_, _00576_);
  and (_04194_, _04134_, _04156_);
  and (_04195_, _04194_, _04141_);
  and (_04196_, _04195_, _04193_);
  not (_04197_, _00276_);
  and (_04198_, _04181_, _04135_);
  and (_04199_, _04198_, _04197_);
  not (_04200_, _43727_);
  and (_04201_, _04142_, _04200_);
  or (_04202_, _04201_, _04199_);
  or (_04203_, _04202_, _04196_);
  or (_04204_, _04203_, _04192_);
  not (_04205_, _00440_);
  and (_04206_, _04173_, _04131_);
  and (_04207_, _04206_, _04205_);
  not (_04208_, _00235_);
  and (_04209_, _04182_, _04156_);
  and (_04210_, _04209_, _04208_);
  or (_04211_, _04210_, _04207_);
  or (_04212_, _04211_, _04204_);
  or (_04213_, _04212_, _04189_);
  or (_04214_, _04213_, _04171_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _04214_, _04164_);
  and (_04215_, _04157_, _04205_);
  and (_04216_, _04152_, _04155_);
  or (_04217_, _04216_, _04215_);
  and (_04218_, _04146_, _04149_);
  and (_04219_, _04161_, _04190_);
  or (_04220_, _04219_, _04218_);
  or (_04221_, _04220_, _04217_);
  and (_04222_, _04186_, _04208_);
  and (_04223_, _04183_, _04185_);
  or (_04224_, _04223_, _04222_);
  and (_04225_, _04174_, _04176_);
  and (_04226_, _04209_, _04197_);
  or (_04227_, _04226_, _04225_);
  or (_04228_, _04227_, _04224_);
  and (_04229_, _04191_, _04180_);
  and (_04230_, _04142_, _04165_);
  and (_04231_, _04198_, _04122_);
  and (_04232_, _04195_, _04200_);
  or (_04233_, _04232_, _04231_);
  or (_04234_, _04233_, _04230_);
  or (_04235_, _04234_, _04229_);
  and (_04236_, _04177_, _04193_);
  and (_04237_, _04206_, _04172_);
  or (_04238_, _04237_, _04236_);
  or (_04239_, _04238_, _04235_);
  or (_04240_, _04239_, _04228_);
  and (_04241_, _04169_, _04159_);
  and (_04242_, _04166_, _04168_);
  or (_04243_, _04242_, _04241_);
  or (_04244_, _04243_, _04240_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _04244_, _04221_);
  and (_04245_, _04146_, _04155_);
  and (_04247_, _04152_, _04205_);
  or (_04248_, _04247_, _04245_);
  and (_04249_, _04157_, _04172_);
  and (_04250_, _04161_, _04180_);
  or (_04251_, _04250_, _04249_);
  or (_04252_, _04251_, _04248_);
  and (_04253_, _04169_, _04190_);
  and (_04254_, _04166_, _04159_);
  or (_04255_, _04254_, _04253_);
  and (_04256_, _04209_, _04122_);
  and (_04257_, _04186_, _04197_);
  or (_04258_, _04257_, _04256_);
  and (_04259_, _04183_, _04208_);
  and (_04260_, _04177_, _04200_);
  or (_04261_, _04260_, _04259_);
  or (_04262_, _04261_, _04258_);
  and (_04263_, _04191_, _04185_);
  and (_04264_, _04142_, _04168_);
  and (_04265_, _04198_, _04149_);
  and (_04266_, _04195_, _04165_);
  or (_04267_, _04266_, _04265_);
  or (_04268_, _04267_, _04264_);
  or (_04269_, _04268_, _04263_);
  and (_04270_, _04174_, _04193_);
  and (_04271_, _04206_, _04176_);
  or (_04272_, _04271_, _04270_);
  or (_04273_, _04272_, _04269_);
  or (_04274_, _04273_, _04262_);
  or (_04275_, _04274_, _04255_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _04275_, _04252_);
  and (_04276_, _04142_, _04193_);
  and (_04277_, _04161_, _04168_);
  and (_04278_, _04166_, _04200_);
  or (_04279_, _04278_, _04277_);
  and (_04280_, _04169_, _04165_);
  and (_04281_, _04209_, _04185_);
  and (_04282_, _04186_, _04180_);
  or (_04283_, _04282_, _04281_);
  and (_04284_, _04183_, _04190_);
  and (_04285_, _04191_, _04159_);
  or (_04286_, _04285_, _04284_);
  or (_04287_, _04286_, _04283_);
  or (_04288_, _04287_, _04280_);
  or (_04289_, _04288_, _04279_);
  and (_04290_, _04177_, _04172_);
  and (_04291_, _04195_, _04176_);
  or (_04292_, _04291_, _04290_);
  and (_04293_, _04206_, _04155_);
  and (_04294_, _04174_, _04205_);
  or (_04295_, _04294_, _04293_);
  or (_04296_, _04295_, _04292_);
  and (_04297_, _04157_, _04149_);
  and (_04298_, _04152_, _04122_);
  or (_04299_, _04298_, _04297_);
  and (_04300_, _04146_, _04197_);
  and (_04301_, _04198_, _04208_);
  or (_04302_, _04301_, _04300_);
  or (_04303_, _04302_, _04299_);
  or (_04304_, _04303_, _04296_);
  or (_04305_, _04304_, _04289_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _04305_, _04276_);
  not (_04306_, _00404_);
  and (_04307_, _04146_, _04306_);
  not (_04308_, _00127_);
  and (_04309_, _04161_, _04308_);
  or (_04310_, _04309_, _04307_);
  not (_04311_, _00445_);
  and (_04312_, _04152_, _04311_);
  not (_04313_, _00486_);
  and (_04314_, _04157_, _04313_);
  or (_04315_, _04314_, _04312_);
  or (_04316_, _04315_, _04310_);
  not (_04317_, _00045_);
  and (_04318_, _04166_, _04317_);
  not (_04319_, _00086_);
  and (_04320_, _04169_, _04319_);
  or (_04321_, _04320_, _04318_);
  not (_04322_, _00584_);
  and (_04323_, _04174_, _04322_);
  not (_04324_, _00322_);
  and (_04325_, _04209_, _04324_);
  or (_04326_, _04325_, _04323_);
  not (_04327_, _00527_);
  and (_04328_, _04206_, _04327_);
  not (_04329_, _00240_);
  and (_04330_, _04183_, _04329_);
  or (_04331_, _04330_, _04328_);
  or (_04332_, _04331_, _04326_);
  not (_04333_, _00199_);
  and (_04334_, _04191_, _04333_);
  not (_04335_, _43773_);
  and (_04336_, _04195_, _04335_);
  not (_04337_, _00363_);
  and (_04338_, _04198_, _04337_);
  not (_04339_, _00004_);
  and (_04340_, _04142_, _04339_);
  or (_04341_, _04340_, _04338_);
  or (_04342_, _04341_, _04336_);
  or (_04343_, _04342_, _04334_);
  not (_04344_, _00281_);
  and (_04346_, _04186_, _04344_);
  not (_04347_, _43732_);
  and (_04348_, _04177_, _04347_);
  or (_04349_, _04348_, _04346_);
  or (_04350_, _04349_, _04343_);
  or (_04351_, _04350_, _04332_);
  or (_04352_, _04351_, _04321_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _04352_, _04316_);
  not (_04353_, _00409_);
  and (_04354_, _04146_, _04353_);
  not (_04355_, _00135_);
  and (_04356_, _04161_, _04355_);
  or (_04357_, _04356_, _04354_);
  not (_04358_, _00450_);
  and (_04359_, _04152_, _04358_);
  not (_04360_, _00491_);
  and (_04361_, _04157_, _04360_);
  or (_04362_, _04361_, _04359_);
  or (_04363_, _04362_, _04357_);
  not (_04364_, _00050_);
  and (_04365_, _04166_, _04364_);
  not (_04366_, _00091_);
  and (_04367_, _04169_, _04366_);
  or (_04368_, _04367_, _04365_);
  not (_04369_, _00592_);
  and (_04370_, _04174_, _04369_);
  not (_04371_, _00327_);
  and (_04372_, _04209_, _04371_);
  or (_04373_, _04372_, _04370_);
  not (_04374_, _00532_);
  and (_04375_, _04206_, _04374_);
  not (_04376_, _00245_);
  and (_04377_, _04183_, _04376_);
  or (_04378_, _04377_, _04375_);
  or (_04379_, _04378_, _04373_);
  not (_04380_, _00204_);
  and (_04381_, _04191_, _04380_);
  not (_04382_, _43778_);
  and (_04383_, _04195_, _04382_);
  not (_04384_, _00368_);
  and (_04385_, _04198_, _04384_);
  not (_04386_, _00009_);
  and (_04387_, _04142_, _04386_);
  or (_04388_, _04387_, _04385_);
  or (_04389_, _04388_, _04383_);
  or (_04390_, _04389_, _04381_);
  not (_04391_, _00286_);
  and (_04392_, _04186_, _04391_);
  not (_04393_, _43737_);
  and (_04394_, _04177_, _04393_);
  or (_04395_, _04394_, _04392_);
  or (_04396_, _04395_, _04390_);
  or (_04397_, _04396_, _04379_);
  or (_04398_, _04397_, _04368_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _04398_, _04363_);
  not (_04399_, _00455_);
  and (_04400_, _04152_, _04399_);
  not (_04401_, _00146_);
  and (_04402_, _04161_, _04401_);
  or (_04403_, _04402_, _04400_);
  not (_04404_, _00496_);
  and (_04405_, _04157_, _04404_);
  not (_04406_, _00414_);
  and (_04407_, _04146_, _04406_);
  or (_04408_, _04407_, _04405_);
  or (_04409_, _04408_, _04403_);
  not (_04410_, _00096_);
  and (_04411_, _04169_, _04410_);
  not (_04412_, _00055_);
  and (_04413_, _04166_, _04412_);
  or (_04414_, _04413_, _04411_);
  not (_04415_, _00537_);
  and (_04416_, _04206_, _04415_);
  not (_04417_, _43742_);
  and (_04418_, _04177_, _04417_);
  or (_04419_, _04418_, _04416_);
  not (_04420_, _00332_);
  and (_04421_, _04209_, _04420_);
  not (_04422_, _00250_);
  and (_04423_, _04183_, _04422_);
  or (_04424_, _04423_, _04421_);
  or (_04425_, _04424_, _04419_);
  not (_04426_, _00209_);
  and (_04427_, _04191_, _04426_);
  not (_04428_, _00373_);
  and (_04429_, _04198_, _04428_);
  not (_04430_, _43783_);
  and (_04431_, _04195_, _04430_);
  not (_04432_, _00014_);
  and (_04433_, _04142_, _04432_);
  or (_04434_, _04433_, _04431_);
  or (_04435_, _04434_, _04429_);
  or (_04436_, _04435_, _04427_);
  not (_04437_, _00597_);
  and (_04438_, _04174_, _04437_);
  not (_04439_, _00291_);
  and (_04440_, _04186_, _04439_);
  or (_04441_, _04440_, _04438_);
  or (_04442_, _04441_, _04436_);
  or (_04443_, _04442_, _04425_);
  or (_04445_, _04443_, _04414_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _04445_, _04409_);
  not (_04446_, _00419_);
  and (_04447_, _04146_, _04446_);
  not (_04448_, _00157_);
  and (_04449_, _04161_, _04448_);
  or (_04450_, _04449_, _04447_);
  not (_04451_, _00460_);
  and (_04452_, _04152_, _04451_);
  not (_04453_, _00501_);
  and (_04454_, _04157_, _04453_);
  or (_04455_, _04454_, _04452_);
  or (_04456_, _04455_, _04450_);
  not (_04457_, _00060_);
  and (_04458_, _04166_, _04457_);
  not (_04459_, _00101_);
  and (_04460_, _04169_, _04459_);
  or (_04461_, _04460_, _04458_);
  not (_04462_, _00602_);
  and (_04463_, _04174_, _04462_);
  not (_04464_, _00337_);
  and (_04465_, _04209_, _04464_);
  or (_04466_, _04465_, _04463_);
  not (_04467_, _00542_);
  and (_04468_, _04206_, _04467_);
  not (_04469_, _00255_);
  and (_04470_, _04183_, _04469_);
  or (_04471_, _04470_, _04468_);
  or (_04472_, _04471_, _04466_);
  not (_04473_, _00214_);
  and (_04474_, _04191_, _04473_);
  not (_04475_, _43788_);
  and (_04476_, _04195_, _04475_);
  not (_04477_, _00378_);
  and (_04478_, _04198_, _04477_);
  not (_04479_, _00019_);
  and (_04480_, _04142_, _04479_);
  or (_04481_, _04480_, _04478_);
  or (_04482_, _04481_, _04476_);
  or (_04483_, _04482_, _04474_);
  not (_04484_, _00296_);
  and (_04485_, _04186_, _04484_);
  not (_04486_, _43747_);
  and (_04487_, _04177_, _04486_);
  or (_04488_, _04487_, _04485_);
  or (_04489_, _04488_, _04483_);
  or (_04490_, _04489_, _04472_);
  or (_04491_, _04490_, _04461_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _04491_, _04456_);
  not (_04492_, _00424_);
  and (_04493_, _04146_, _04492_);
  not (_04494_, _00168_);
  and (_04495_, _04161_, _04494_);
  or (_04496_, _04495_, _04493_);
  not (_04497_, _00465_);
  and (_04498_, _04152_, _04497_);
  not (_04499_, _00506_);
  and (_04500_, _04157_, _04499_);
  or (_04501_, _04500_, _04498_);
  or (_04502_, _04501_, _04496_);
  not (_04503_, _00065_);
  and (_04504_, _04166_, _04503_);
  not (_04505_, _00106_);
  and (_04506_, _04169_, _04505_);
  or (_04507_, _04506_, _04504_);
  not (_04508_, _00607_);
  and (_04509_, _04174_, _04508_);
  not (_04510_, _00342_);
  and (_04511_, _04209_, _04510_);
  or (_04512_, _04511_, _04509_);
  not (_04513_, _00550_);
  and (_04514_, _04206_, _04513_);
  not (_04515_, _00260_);
  and (_04516_, _04183_, _04515_);
  or (_04517_, _04516_, _04514_);
  or (_04518_, _04517_, _04512_);
  not (_04519_, _00219_);
  and (_04520_, _04191_, _04519_);
  not (_04521_, _43793_);
  and (_04522_, _04195_, _04521_);
  not (_04523_, _00383_);
  and (_04524_, _04198_, _04523_);
  not (_04525_, _00024_);
  and (_04526_, _04142_, _04525_);
  or (_04527_, _04526_, _04524_);
  or (_04528_, _04527_, _04522_);
  or (_04529_, _04528_, _04520_);
  not (_04530_, _00301_);
  and (_04531_, _04186_, _04530_);
  not (_04532_, _43752_);
  and (_04533_, _04177_, _04532_);
  or (_04534_, _04533_, _04531_);
  or (_04535_, _04534_, _04529_);
  or (_04536_, _04535_, _04518_);
  or (_04537_, _04536_, _04507_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _04537_, _04502_);
  not (_04538_, _00511_);
  and (_04539_, _04157_, _04538_);
  not (_04540_, _00429_);
  and (_04541_, _04146_, _04540_);
  or (_04543_, _04541_, _04539_);
  not (_04544_, _00470_);
  and (_04545_, _04152_, _04544_);
  not (_04546_, _00179_);
  and (_04547_, _04161_, _04546_);
  or (_04548_, _04547_, _04545_);
  or (_04549_, _04548_, _04543_);
  not (_04550_, _00111_);
  and (_04551_, _04169_, _04550_);
  not (_04552_, _00070_);
  and (_04553_, _04166_, _04552_);
  or (_04554_, _04553_, _04551_);
  not (_04555_, _00347_);
  and (_04556_, _04209_, _04555_);
  not (_04557_, _00306_);
  and (_04558_, _04186_, _04557_);
  or (_04559_, _04558_, _04556_);
  not (_04560_, _00265_);
  and (_04561_, _04183_, _04560_);
  not (_04562_, _43757_);
  and (_04563_, _04177_, _04562_);
  or (_04564_, _04563_, _04561_);
  or (_04565_, _04564_, _04559_);
  not (_04566_, _00224_);
  and (_04567_, _04191_, _04566_);
  not (_04568_, _00029_);
  and (_04569_, _04142_, _04568_);
  not (_04570_, _00388_);
  and (_04571_, _04198_, _04570_);
  not (_04572_, _43798_);
  and (_04573_, _04195_, _04572_);
  or (_04574_, _04573_, _04571_);
  or (_04575_, _04574_, _04569_);
  or (_04576_, _04575_, _04567_);
  not (_04577_, _00612_);
  and (_04578_, _04174_, _04577_);
  not (_04579_, _00558_);
  and (_04580_, _04206_, _04579_);
  or (_04581_, _04580_, _04578_);
  or (_04582_, _04581_, _04576_);
  or (_04583_, _04582_, _04565_);
  or (_04584_, _04583_, _04554_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _04584_, _04549_);
  not (_04585_, _00434_);
  and (_04586_, _04146_, _04585_);
  not (_04587_, _00475_);
  and (_04588_, _04152_, _04587_);
  or (_04589_, _04588_, _04586_);
  not (_04590_, _00516_);
  and (_04591_, _04157_, _04590_);
  not (_04592_, _00188_);
  and (_04593_, _04161_, _04592_);
  or (_04594_, _04593_, _04591_);
  or (_04595_, _04594_, _04589_);
  not (_04596_, _00116_);
  and (_04597_, _04169_, _04596_);
  not (_04598_, _00075_);
  and (_04599_, _04166_, _04598_);
  or (_04600_, _04599_, _04597_);
  not (_04601_, _00352_);
  and (_04602_, _04209_, _04601_);
  not (_04603_, _00311_);
  and (_04604_, _04186_, _04603_);
  or (_04605_, _04604_, _04602_);
  not (_04606_, _00270_);
  and (_04607_, _04183_, _04606_);
  not (_04608_, _43762_);
  and (_04609_, _04177_, _04608_);
  or (_04610_, _04609_, _04607_);
  or (_04611_, _04610_, _04605_);
  not (_04612_, _00229_);
  and (_04613_, _04191_, _04612_);
  not (_04614_, _00034_);
  and (_04615_, _04142_, _04614_);
  not (_04616_, _00393_);
  and (_04617_, _04198_, _04616_);
  not (_04618_, _43803_);
  and (_04619_, _04195_, _04618_);
  or (_04620_, _04619_, _04617_);
  or (_04621_, _04620_, _04615_);
  or (_04622_, _04621_, _04613_);
  not (_04623_, _00617_);
  and (_04624_, _04174_, _04623_);
  not (_04625_, _00566_);
  and (_04626_, _04206_, _04625_);
  or (_04627_, _04626_, _04624_);
  or (_04628_, _04627_, _04622_);
  or (_04629_, _04628_, _04611_);
  or (_04630_, _04629_, _04600_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _04630_, _04595_);
  and (_04631_, _04157_, _04311_);
  and (_04632_, _04161_, _04319_);
  or (_04633_, _04632_, _04631_);
  and (_04634_, _04152_, _04306_);
  and (_04635_, _04146_, _04337_);
  or (_04636_, _04635_, _04634_);
  or (_04637_, _04636_, _04633_);
  and (_04638_, _04209_, _04344_);
  and (_04639_, _04183_, _04333_);
  or (_04640_, _04639_, _04638_);
  and (_04642_, _04206_, _04313_);
  and (_04643_, _04186_, _04329_);
  or (_04644_, _04643_, _04642_);
  or (_04645_, _04644_, _04640_);
  and (_04646_, _04191_, _04308_);
  and (_04647_, _04198_, _04324_);
  and (_04648_, _04195_, _04347_);
  and (_04649_, _04142_, _04335_);
  or (_04650_, _04649_, _04648_);
  or (_04651_, _04650_, _04647_);
  or (_04652_, _04651_, _04646_);
  and (_04653_, _04177_, _04322_);
  and (_04654_, _04174_, _04327_);
  or (_04655_, _04654_, _04653_);
  or (_04656_, _04655_, _04652_);
  or (_04657_, _04656_, _04645_);
  and (_04658_, _04169_, _04317_);
  and (_04659_, _04166_, _04339_);
  or (_04660_, _04659_, _04658_);
  or (_04661_, _04660_, _04657_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _04661_, _04637_);
  and (_04662_, _04157_, _04358_);
  and (_04663_, _04152_, _04353_);
  or (_04664_, _04663_, _04662_);
  and (_04665_, _04146_, _04384_);
  and (_04666_, _04161_, _04366_);
  or (_04667_, _04666_, _04665_);
  or (_04668_, _04667_, _04664_);
  and (_04669_, _04186_, _04376_);
  and (_04670_, _04183_, _04380_);
  or (_04671_, _04670_, _04669_);
  and (_04672_, _04174_, _04374_);
  and (_04673_, _04209_, _04391_);
  or (_04674_, _04673_, _04672_);
  or (_04675_, _04674_, _04671_);
  and (_04676_, _04191_, _04355_);
  and (_04677_, _04142_, _04382_);
  and (_04678_, _04198_, _04371_);
  and (_04679_, _04195_, _04393_);
  or (_04680_, _04679_, _04678_);
  or (_04681_, _04680_, _04677_);
  or (_04682_, _04681_, _04676_);
  and (_04683_, _04177_, _04369_);
  and (_04684_, _04206_, _04360_);
  or (_04685_, _04684_, _04683_);
  or (_04686_, _04685_, _04682_);
  or (_04687_, _04686_, _04675_);
  and (_04688_, _04169_, _04364_);
  and (_04689_, _04166_, _04386_);
  or (_04690_, _04689_, _04688_);
  or (_04691_, _04690_, _04687_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _04691_, _04668_);
  and (_04692_, _04157_, _04399_);
  and (_04693_, _04161_, _04410_);
  or (_04694_, _04693_, _04692_);
  and (_04695_, _04152_, _04406_);
  and (_04696_, _04146_, _04428_);
  or (_04697_, _04696_, _04695_);
  or (_04698_, _04697_, _04694_);
  and (_04699_, _04177_, _04437_);
  and (_04700_, _04174_, _04415_);
  or (_04701_, _04700_, _04699_);
  and (_04702_, _04209_, _04439_);
  and (_04703_, _04183_, _04426_);
  or (_04704_, _04703_, _04702_);
  or (_04705_, _04704_, _04701_);
  and (_04706_, _04191_, _04401_);
  and (_04707_, _04198_, _04420_);
  and (_04708_, _04195_, _04417_);
  and (_04709_, _04142_, _04430_);
  or (_04710_, _04709_, _04708_);
  or (_04711_, _04710_, _04707_);
  or (_04712_, _04711_, _04706_);
  and (_04713_, _04206_, _04404_);
  and (_04714_, _04186_, _04422_);
  or (_04715_, _04714_, _04713_);
  or (_04716_, _04715_, _04712_);
  or (_04717_, _04716_, _04705_);
  and (_04718_, _04169_, _04412_);
  and (_04719_, _04166_, _04432_);
  or (_04720_, _04719_, _04718_);
  or (_04721_, _04720_, _04717_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _04721_, _04698_);
  and (_04722_, _04152_, _04446_);
  and (_04723_, _04157_, _04451_);
  or (_04724_, _04723_, _04722_);
  and (_04725_, _04146_, _04477_);
  and (_04726_, _04161_, _04459_);
  or (_04727_, _04726_, _04725_);
  or (_04728_, _04727_, _04724_);
  and (_04729_, _04186_, _04469_);
  and (_04730_, _04183_, _04473_);
  or (_04731_, _04730_, _04729_);
  and (_04732_, _04177_, _04462_);
  and (_04733_, _04206_, _04453_);
  or (_04734_, _04733_, _04732_);
  or (_04735_, _04734_, _04731_);
  and (_04736_, _04191_, _04448_);
  and (_04737_, _04195_, _04486_);
  and (_04738_, _04198_, _04464_);
  and (_04739_, _04142_, _04475_);
  or (_04740_, _04739_, _04738_);
  or (_04741_, _04740_, _04737_);
  or (_04742_, _04741_, _04736_);
  and (_04743_, _04174_, _04467_);
  and (_04744_, _04209_, _04484_);
  or (_04745_, _04744_, _04743_);
  or (_04746_, _04745_, _04742_);
  or (_04747_, _04746_, _04735_);
  and (_04748_, _04169_, _04457_);
  and (_04749_, _04166_, _04479_);
  or (_04750_, _04749_, _04748_);
  or (_04751_, _04750_, _04747_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _04751_, _04728_);
  and (_04752_, _04157_, _04497_);
  and (_04753_, _04146_, _04523_);
  or (_04754_, _04753_, _04752_);
  and (_04755_, _04152_, _04492_);
  and (_04756_, _04161_, _04505_);
  or (_04757_, _04756_, _04755_);
  or (_04758_, _04757_, _04754_);
  and (_04759_, _04186_, _04515_);
  and (_04760_, _04183_, _04519_);
  or (_04761_, _04760_, _04759_);
  and (_04762_, _04174_, _04513_);
  and (_04763_, _04209_, _04530_);
  or (_04764_, _04763_, _04762_);
  or (_04765_, _04764_, _04761_);
  and (_04766_, _04191_, _04494_);
  and (_04767_, _04142_, _04521_);
  and (_04768_, _04198_, _04510_);
  and (_04769_, _04195_, _04532_);
  or (_04770_, _04769_, _04768_);
  or (_04771_, _04770_, _04767_);
  or (_04772_, _04771_, _04766_);
  and (_04773_, _04177_, _04508_);
  and (_04774_, _04206_, _04499_);
  or (_04775_, _04774_, _04773_);
  or (_04776_, _04775_, _04772_);
  or (_04777_, _04776_, _04765_);
  and (_04778_, _04169_, _04503_);
  and (_04779_, _04166_, _04525_);
  or (_04780_, _04779_, _04778_);
  or (_04781_, _04780_, _04777_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _04781_, _04758_);
  and (_04782_, _04152_, _04540_);
  and (_04783_, _04157_, _04544_);
  or (_04784_, _04783_, _04782_);
  and (_04785_, _04146_, _04570_);
  and (_04786_, _04161_, _04550_);
  or (_04787_, _04786_, _04785_);
  or (_04788_, _04787_, _04784_);
  and (_04789_, _04186_, _04560_);
  and (_04790_, _04183_, _04566_);
  or (_04791_, _04790_, _04789_);
  and (_04792_, _04177_, _04577_);
  and (_04793_, _04206_, _04538_);
  or (_04794_, _04793_, _04792_);
  or (_04795_, _04794_, _04791_);
  and (_04796_, _04191_, _04546_);
  and (_04797_, _04195_, _04562_);
  and (_04798_, _04198_, _04555_);
  and (_04799_, _04142_, _04572_);
  or (_04800_, _04799_, _04798_);
  or (_04801_, _04800_, _04797_);
  or (_04802_, _04801_, _04796_);
  and (_04803_, _04174_, _04579_);
  and (_04804_, _04209_, _04557_);
  or (_04805_, _04804_, _04803_);
  or (_04806_, _04805_, _04802_);
  or (_04807_, _04806_, _04795_);
  and (_04808_, _04169_, _04552_);
  and (_04809_, _04166_, _04568_);
  or (_04810_, _04809_, _04808_);
  or (_04811_, _04810_, _04807_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _04811_, _04788_);
  and (_04812_, _04157_, _04587_);
  and (_04813_, _04146_, _04616_);
  or (_04814_, _04813_, _04812_);
  and (_04815_, _04152_, _04585_);
  and (_04816_, _04161_, _04596_);
  or (_04817_, _04816_, _04815_);
  or (_04818_, _04817_, _04814_);
  and (_04819_, _04186_, _04606_);
  and (_04820_, _04183_, _04612_);
  or (_04821_, _04820_, _04819_);
  and (_04822_, _04174_, _04625_);
  and (_04823_, _04209_, _04603_);
  or (_04824_, _04823_, _04822_);
  or (_04825_, _04824_, _04821_);
  and (_04826_, _04191_, _04592_);
  and (_04827_, _04142_, _04618_);
  and (_04828_, _04198_, _04601_);
  and (_04829_, _04195_, _04608_);
  or (_04830_, _04829_, _04828_);
  or (_04831_, _04830_, _04827_);
  or (_04832_, _04831_, _04826_);
  and (_04833_, _04177_, _04623_);
  and (_04834_, _04206_, _04590_);
  or (_04835_, _04834_, _04833_);
  or (_04836_, _04835_, _04832_);
  or (_04837_, _04836_, _04825_);
  and (_04838_, _04169_, _04598_);
  and (_04839_, _04166_, _04614_);
  or (_04840_, _04839_, _04838_);
  or (_04841_, _04840_, _04837_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _04841_, _04818_);
  and (_04842_, _04161_, _04339_);
  and (_04843_, _04157_, _04337_);
  or (_04844_, _04843_, _04842_);
  and (_04845_, _04152_, _04324_);
  and (_04846_, _04146_, _04344_);
  or (_04847_, _04846_, _04845_);
  or (_04848_, _04847_, _04844_);
  and (_04849_, _04183_, _04319_);
  and (_04850_, _04177_, _04313_);
  or (_04851_, _04850_, _04849_);
  and (_04852_, _04209_, _04333_);
  and (_04853_, _04206_, _04306_);
  or (_04854_, _04853_, _04852_);
  or (_04855_, _04854_, _04851_);
  and (_04856_, _04191_, _04317_);
  and (_04857_, _04198_, _04329_);
  and (_04858_, _04142_, _04322_);
  and (_04859_, _04195_, _04327_);
  or (_04860_, _04859_, _04858_);
  or (_04861_, _04860_, _04857_);
  or (_04862_, _04861_, _04856_);
  and (_04863_, _04186_, _04308_);
  and (_04864_, _04174_, _04311_);
  or (_04865_, _04864_, _04863_);
  or (_04866_, _04865_, _04862_);
  or (_04867_, _04866_, _04855_);
  and (_04868_, _04166_, _04347_);
  and (_04869_, _04169_, _04335_);
  or (_04870_, _04869_, _04868_);
  or (_04871_, _04870_, _04867_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _04871_, _04848_);
  and (_04872_, _04152_, _04371_);
  and (_04873_, _04157_, _04384_);
  or (_04874_, _04873_, _04872_);
  and (_04875_, _04146_, _04391_);
  and (_04876_, _04161_, _04386_);
  or (_04877_, _04876_, _04875_);
  or (_04878_, _04877_, _04874_);
  and (_04879_, _04177_, _04360_);
  and (_04880_, _04183_, _04366_);
  or (_04881_, _04880_, _04879_);
  and (_04882_, _04206_, _04353_);
  and (_04883_, _04209_, _04380_);
  or (_04884_, _04883_, _04882_);
  or (_04885_, _04884_, _04881_);
  and (_04886_, _04191_, _04364_);
  and (_04887_, _04142_, _04369_);
  and (_04888_, _04195_, _04374_);
  and (_04889_, _04198_, _04376_);
  or (_04890_, _04889_, _04888_);
  or (_04891_, _04890_, _04887_);
  or (_04892_, _04891_, _04886_);
  and (_04893_, _04174_, _04358_);
  and (_04894_, _04186_, _04355_);
  or (_04895_, _04894_, _04893_);
  or (_04896_, _04895_, _04892_);
  or (_04897_, _04896_, _04885_);
  and (_04898_, _04166_, _04393_);
  and (_04899_, _04169_, _04382_);
  or (_04900_, _04899_, _04898_);
  or (_04901_, _04900_, _04897_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _04901_, _04878_);
  and (_04902_, _04142_, _04437_);
  and (_04903_, _04161_, _04432_);
  and (_04904_, _04166_, _04417_);
  or (_04905_, _04904_, _04903_);
  and (_04906_, _04169_, _04430_);
  and (_04907_, _04209_, _04426_);
  and (_04908_, _04186_, _04401_);
  or (_04909_, _04908_, _04907_);
  and (_04910_, _04183_, _04410_);
  and (_04911_, _04191_, _04412_);
  or (_04912_, _04911_, _04910_);
  or (_04913_, _04912_, _04909_);
  or (_04914_, _04913_, _04906_);
  or (_04915_, _04914_, _04905_);
  and (_04916_, _04177_, _04404_);
  and (_04917_, _04195_, _04415_);
  or (_04918_, _04917_, _04916_);
  and (_04919_, _04206_, _04406_);
  and (_04920_, _04174_, _04399_);
  or (_04921_, _04920_, _04919_);
  or (_04922_, _04921_, _04918_);
  and (_04923_, _04157_, _04428_);
  and (_04924_, _04152_, _04420_);
  or (_04925_, _04924_, _04923_);
  and (_04926_, _04146_, _04439_);
  and (_04927_, _04198_, _04422_);
  or (_04928_, _04927_, _04926_);
  or (_04929_, _04928_, _04925_);
  or (_04930_, _04929_, _04922_);
  or (_04931_, _04930_, _04915_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _04931_, _04902_);
  and (_04932_, _04142_, _04462_);
  and (_04933_, _04161_, _04479_);
  and (_04934_, _04166_, _04486_);
  or (_04935_, _04934_, _04933_);
  and (_04936_, _04169_, _04475_);
  and (_04937_, _04209_, _04473_);
  and (_04938_, _04186_, _04448_);
  or (_04939_, _04938_, _04937_);
  and (_04940_, _04183_, _04459_);
  and (_04941_, _04191_, _04457_);
  or (_04942_, _04941_, _04940_);
  or (_04943_, _04942_, _04939_);
  or (_04944_, _04943_, _04936_);
  or (_04945_, _04944_, _04935_);
  and (_04946_, _04177_, _04453_);
  and (_04947_, _04195_, _04467_);
  or (_04948_, _04947_, _04946_);
  and (_04949_, _04206_, _04446_);
  and (_04950_, _04174_, _04451_);
  or (_04951_, _04950_, _04949_);
  or (_04952_, _04951_, _04948_);
  and (_04953_, _04157_, _04477_);
  and (_04954_, _04152_, _04464_);
  or (_04955_, _04954_, _04953_);
  and (_04956_, _04146_, _04484_);
  and (_04957_, _04198_, _04469_);
  or (_04958_, _04957_, _04956_);
  or (_04959_, _04958_, _04955_);
  or (_04960_, _04959_, _04952_);
  or (_04961_, _04960_, _04945_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _04961_, _04932_);
  and (_04962_, _04152_, _04510_);
  and (_04963_, _04161_, _04525_);
  or (_04964_, _04963_, _04962_);
  and (_04965_, _04157_, _04523_);
  and (_04966_, _04146_, _04530_);
  or (_04967_, _04966_, _04965_);
  or (_04968_, _04967_, _04964_);
  and (_04969_, _04177_, _04499_);
  and (_04970_, _04183_, _04505_);
  or (_04971_, _04970_, _04969_);
  and (_04972_, _04206_, _04492_);
  and (_04973_, _04209_, _04519_);
  or (_04974_, _04973_, _04972_);
  or (_04975_, _04974_, _04971_);
  and (_04976_, _04191_, _04503_);
  and (_04977_, _04142_, _04508_);
  and (_04978_, _04195_, _04513_);
  and (_04979_, _04198_, _04515_);
  or (_04980_, _04979_, _04978_);
  or (_04981_, _04980_, _04977_);
  or (_04982_, _04981_, _04976_);
  and (_04983_, _04174_, _04497_);
  and (_04984_, _04186_, _04494_);
  or (_04985_, _04984_, _04983_);
  or (_04986_, _04985_, _04982_);
  or (_04987_, _04986_, _04975_);
  and (_04988_, _04166_, _04532_);
  and (_04989_, _04169_, _04521_);
  or (_04990_, _04989_, _04988_);
  or (_04991_, _04990_, _04987_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _04991_, _04968_);
  and (_04992_, _04152_, _04555_);
  and (_04993_, _04157_, _04570_);
  or (_04994_, _04993_, _04992_);
  and (_04995_, _04146_, _04557_);
  and (_04996_, _04161_, _04568_);
  or (_04997_, _04996_, _04995_);
  or (_04998_, _04997_, _04994_);
  and (_04999_, _04177_, _04538_);
  and (_05000_, _04183_, _04550_);
  or (_05001_, _05000_, _04999_);
  and (_05002_, _04206_, _04540_);
  and (_05003_, _04209_, _04566_);
  or (_05004_, _05003_, _05002_);
  or (_05005_, _05004_, _05001_);
  and (_05006_, _04191_, _04552_);
  and (_05007_, _04142_, _04577_);
  and (_05008_, _04195_, _04579_);
  and (_05009_, _04198_, _04560_);
  or (_05010_, _05009_, _05008_);
  or (_05011_, _05010_, _05007_);
  or (_05012_, _05011_, _05006_);
  and (_05013_, _04174_, _04544_);
  and (_05014_, _04186_, _04546_);
  or (_05015_, _05014_, _05013_);
  or (_05016_, _05015_, _05012_);
  or (_05017_, _05016_, _05005_);
  and (_05018_, _04166_, _04562_);
  and (_05019_, _04169_, _04572_);
  or (_05020_, _05019_, _05018_);
  or (_05021_, _05020_, _05017_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _05021_, _04998_);
  and (_05022_, _04142_, _04623_);
  and (_05023_, _04161_, _04614_);
  and (_05024_, _04166_, _04608_);
  or (_05025_, _05024_, _05023_);
  and (_05026_, _04169_, _04618_);
  and (_05027_, _04209_, _04612_);
  and (_05028_, _04186_, _04592_);
  or (_05029_, _05028_, _05027_);
  and (_05030_, _04183_, _04596_);
  and (_05031_, _04191_, _04598_);
  or (_05032_, _05031_, _05030_);
  or (_05033_, _05032_, _05029_);
  or (_05034_, _05033_, _05026_);
  or (_05035_, _05034_, _05025_);
  and (_05036_, _04177_, _04590_);
  and (_05037_, _04195_, _04625_);
  or (_05038_, _05037_, _05036_);
  and (_05039_, _04206_, _04585_);
  and (_05040_, _04174_, _04587_);
  or (_05041_, _05040_, _05039_);
  or (_05042_, _05041_, _05038_);
  and (_05043_, _04157_, _04616_);
  and (_05044_, _04152_, _04601_);
  or (_05045_, _05044_, _05043_);
  and (_05046_, _04146_, _04603_);
  and (_05047_, _04198_, _04606_);
  or (_05048_, _05047_, _05046_);
  or (_05049_, _05048_, _05045_);
  or (_05050_, _05049_, _05042_);
  or (_05051_, _05050_, _05035_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _05051_, _05022_);
  and (_05052_, _04157_, _04306_);
  and (_05053_, _04146_, _04324_);
  or (_05054_, _05053_, _05052_);
  and (_05055_, _04152_, _04337_);
  and (_05056_, _04161_, _04317_);
  or (_05057_, _05056_, _05055_);
  or (_05058_, _05057_, _05054_);
  and (_05059_, _04166_, _04335_);
  and (_05060_, _04169_, _04339_);
  or (_05061_, _05060_, _05059_);
  and (_05062_, _04174_, _04313_);
  and (_05063_, _04177_, _04327_);
  or (_05064_, _05063_, _05062_);
  and (_05065_, _04183_, _04308_);
  and (_05066_, _04186_, _04333_);
  or (_05067_, _05066_, _05065_);
  or (_05068_, _05067_, _05064_);
  and (_05069_, _04191_, _04319_);
  and (_05070_, _04195_, _04322_);
  and (_05071_, _04198_, _04344_);
  and (_05072_, _04142_, _04347_);
  or (_05073_, _05072_, _05071_);
  or (_05074_, _05073_, _05070_);
  or (_05075_, _05074_, _05069_);
  and (_05076_, _04206_, _04311_);
  and (_05077_, _04209_, _04329_);
  or (_05078_, _05077_, _05076_);
  or (_05079_, _05078_, _05075_);
  or (_05080_, _05079_, _05068_);
  or (_05082_, _05080_, _05061_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _05082_, _05058_);
  and (_05085_, _04157_, _04353_);
  and (_05087_, _04146_, _04371_);
  or (_05089_, _05087_, _05085_);
  and (_05091_, _04152_, _04384_);
  and (_05093_, _04161_, _04364_);
  or (_05094_, _05093_, _05091_);
  or (_05095_, _05094_, _05089_);
  and (_05096_, _04166_, _04382_);
  and (_05097_, _04169_, _04386_);
  or (_05098_, _05097_, _05096_);
  and (_05099_, _04183_, _04355_);
  and (_05101_, _04186_, _04380_);
  or (_05102_, _05101_, _05099_);
  and (_05104_, _04174_, _04360_);
  and (_05105_, _04209_, _04376_);
  or (_05106_, _05105_, _05104_);
  or (_05108_, _05106_, _05102_);
  and (_05109_, _04191_, _04366_);
  and (_05110_, _04142_, _04393_);
  and (_05112_, _04195_, _04369_);
  and (_05113_, _04198_, _04391_);
  or (_05114_, _05113_, _05112_);
  or (_05116_, _05114_, _05110_);
  or (_05117_, _05116_, _05109_);
  and (_05118_, _04177_, _04374_);
  and (_05120_, _04206_, _04358_);
  or (_05121_, _05120_, _05118_);
  or (_05122_, _05121_, _05117_);
  or (_05124_, _05122_, _05108_);
  or (_05125_, _05124_, _05098_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _05125_, _05095_);
  and (_05127_, _04146_, _04420_);
  and (_05128_, _04152_, _04428_);
  or (_05129_, _05128_, _05127_);
  and (_05131_, _04157_, _04406_);
  and (_05132_, _04161_, _04412_);
  or (_05133_, _05132_, _05131_);
  or (_05134_, _05133_, _05129_);
  and (_05135_, _04166_, _04430_);
  and (_05136_, _04169_, _04432_);
  or (_05137_, _05136_, _05135_);
  and (_05138_, _04174_, _04404_);
  and (_05139_, _04177_, _04415_);
  or (_05140_, _05139_, _05138_);
  and (_05141_, _04183_, _04401_);
  and (_05142_, _04186_, _04426_);
  or (_05143_, _05142_, _05141_);
  or (_05144_, _05143_, _05140_);
  and (_05145_, _04191_, _04410_);
  and (_05146_, _04195_, _04437_);
  and (_05147_, _04198_, _04439_);
  and (_05148_, _04142_, _04417_);
  or (_05149_, _05148_, _05147_);
  or (_05150_, _05149_, _05146_);
  or (_05151_, _05150_, _05145_);
  and (_05153_, _04206_, _04399_);
  and (_05154_, _04209_, _04422_);
  or (_05156_, _05154_, _05153_);
  or (_05157_, _05156_, _05151_);
  or (_05158_, _05157_, _05144_);
  or (_05160_, _05158_, _05137_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _05160_, _05134_);
  and (_05161_, _04157_, _04446_);
  and (_05163_, _04152_, _04477_);
  or (_05164_, _05163_, _05161_);
  and (_05165_, _04146_, _04464_);
  and (_05167_, _04161_, _04457_);
  or (_05168_, _05167_, _05165_);
  or (_05169_, _05168_, _05164_);
  and (_05171_, _04166_, _04475_);
  and (_05172_, _04169_, _04479_);
  or (_05173_, _05172_, _05171_);
  and (_05175_, _04183_, _04448_);
  and (_05176_, _04186_, _04473_);
  or (_05177_, _05176_, _05175_);
  and (_05179_, _04177_, _04467_);
  and (_05180_, _04206_, _04451_);
  or (_05181_, _05180_, _05179_);
  or (_05183_, _05181_, _05177_);
  and (_05184_, _04191_, _04459_);
  and (_05185_, _04195_, _04462_);
  and (_05186_, _04198_, _04484_);
  and (_05187_, _04142_, _04486_);
  or (_05188_, _05187_, _05186_);
  or (_05189_, _05188_, _05185_);
  or (_05190_, _05189_, _05184_);
  and (_05191_, _04174_, _04453_);
  and (_05192_, _04209_, _04469_);
  or (_05193_, _05192_, _05191_);
  or (_05194_, _05193_, _05190_);
  or (_05195_, _05194_, _05183_);
  or (_05196_, _05195_, _05173_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _05196_, _05169_);
  and (_05197_, _04146_, _04510_);
  and (_05198_, _04152_, _04523_);
  or (_05199_, _05198_, _05197_);
  and (_05200_, _04157_, _04492_);
  and (_05201_, _04161_, _04503_);
  or (_05202_, _05201_, _05200_);
  or (_05204_, _05202_, _05199_);
  and (_05205_, _04166_, _04521_);
  and (_05207_, _04169_, _04525_);
  or (_05208_, _05207_, _05205_);
  and (_05209_, _04174_, _04499_);
  and (_05211_, _04177_, _04513_);
  or (_05212_, _05211_, _05209_);
  and (_05213_, _04183_, _04494_);
  and (_05215_, _04186_, _04519_);
  or (_05216_, _05215_, _05213_);
  or (_05217_, _05216_, _05212_);
  and (_05219_, _04191_, _04505_);
  and (_05220_, _04195_, _04508_);
  and (_05221_, _04198_, _04530_);
  and (_05223_, _04142_, _04532_);
  or (_05224_, _05223_, _05221_);
  or (_05225_, _05224_, _05220_);
  or (_05227_, _05225_, _05219_);
  and (_05228_, _04206_, _04497_);
  and (_05229_, _04209_, _04515_);
  or (_05231_, _05229_, _05228_);
  or (_05232_, _05231_, _05227_);
  or (_05233_, _05232_, _05217_);
  or (_05235_, _05233_, _05208_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _05235_, _05204_);
  and (_05236_, _04152_, _04570_);
  and (_05237_, _04161_, _04552_);
  or (_05238_, _05237_, _05236_);
  and (_05239_, _04157_, _04540_);
  and (_05240_, _04146_, _04555_);
  or (_05241_, _05240_, _05239_);
  or (_05242_, _05241_, _05238_);
  and (_05243_, _04166_, _04572_);
  and (_05244_, _04169_, _04568_);
  or (_05245_, _05244_, _05243_);
  and (_05246_, _04174_, _04538_);
  and (_05247_, _04206_, _04544_);
  or (_05248_, _05247_, _05246_);
  and (_05249_, _04209_, _04560_);
  and (_05250_, _04183_, _04546_);
  or (_05251_, _05250_, _05249_);
  or (_05252_, _05251_, _05248_);
  and (_05253_, _04191_, _04550_);
  and (_05254_, _04198_, _04557_);
  and (_05256_, _04195_, _04577_);
  and (_05257_, _04142_, _04562_);
  or (_05259_, _05257_, _05256_);
  or (_05260_, _05259_, _05254_);
  or (_05261_, _05260_, _05253_);
  and (_05263_, _04177_, _04579_);
  and (_05264_, _04186_, _04566_);
  or (_05265_, _05264_, _05263_);
  or (_05267_, _05265_, _05261_);
  or (_05268_, _05267_, _05252_);
  or (_05269_, _05268_, _05245_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _05269_, _05242_);
  and (_05271_, _04157_, _04585_);
  and (_05272_, _04152_, _04616_);
  or (_05274_, _05272_, _05271_);
  and (_05275_, _04146_, _04601_);
  and (_05276_, _04161_, _04598_);
  or (_05278_, _05276_, _05275_);
  or (_05279_, _05278_, _05274_);
  and (_05280_, _04166_, _04618_);
  and (_05282_, _04169_, _04614_);
  or (_05283_, _05282_, _05280_);
  and (_05284_, _04183_, _04592_);
  and (_05286_, _04186_, _04612_);
  or (_05287_, _05286_, _05284_);
  and (_05288_, _04177_, _04625_);
  and (_05289_, _04206_, _04587_);
  or (_05290_, _05289_, _05288_);
  or (_05291_, _05290_, _05287_);
  and (_05292_, _04191_, _04596_);
  and (_05293_, _04195_, _04623_);
  and (_05294_, _04198_, _04603_);
  and (_05295_, _04142_, _04608_);
  or (_05296_, _05295_, _05294_);
  or (_05297_, _05296_, _05293_);
  or (_05298_, _05297_, _05292_);
  and (_05299_, _04174_, _04590_);
  and (_05300_, _04209_, _04606_);
  or (_05301_, _05300_, _05299_);
  or (_05302_, _05301_, _05298_);
  or (_05303_, _05302_, _05291_);
  or (_05304_, _05303_, _05283_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _05304_, _05279_);
  nand (_05305_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_05307_, \oc8051_golden_model_1.PC [3]);
  or (_05308_, \oc8051_golden_model_1.PC [2], _05307_);
  or (_05310_, _05308_, _05305_);
  or (_05311_, _05310_, _00434_);
  not (_05312_, \oc8051_golden_model_1.PC [1]);
  or (_05314_, _05312_, \oc8051_golden_model_1.PC [0]);
  or (_05315_, _05314_, _05308_);
  or (_05316_, _05315_, _00393_);
  and (_05318_, _05316_, _05311_);
  not (_05319_, \oc8051_golden_model_1.PC [2]);
  or (_05320_, _05319_, \oc8051_golden_model_1.PC [3]);
  or (_05322_, _05320_, _05305_);
  or (_05323_, _05322_, _00270_);
  or (_05324_, _05320_, _05314_);
  or (_05326_, _05324_, _00229_);
  and (_05327_, _05326_, _05323_);
  and (_05328_, _05327_, _05318_);
  nand (_05330_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_05331_, _05330_, _05305_);
  or (_05332_, _05331_, _00617_);
  or (_05334_, _05330_, _05314_);
  or (_05335_, _05334_, _00566_);
  and (_05336_, _05335_, _05332_);
  or (_05338_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_05339_, _05338_, _05305_);
  or (_05340_, _05339_, _00075_);
  or (_05341_, _05338_, _05314_);
  or (_05342_, _05341_, _00034_);
  and (_05343_, _05342_, _05340_);
  and (_05344_, _05343_, _05336_);
  and (_05345_, _05344_, _05328_);
  not (_05346_, \oc8051_golden_model_1.PC [0]);
  or (_05347_, \oc8051_golden_model_1.PC [1], _05346_);
  or (_05348_, _05347_, _05330_);
  or (_05349_, _05348_, _00516_);
  or (_05350_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_05351_, _05350_, _05330_);
  or (_05352_, _05351_, _00475_);
  and (_05353_, _05352_, _05349_);
  or (_05354_, _05338_, _05350_);
  or (_05355_, _05354_, _43762_);
  or (_05356_, _05338_, _05347_);
  or (_05357_, _05356_, _43803_);
  and (_05358_, _05357_, _05355_);
  and (_05360_, _05358_, _05353_);
  or (_05361_, _05347_, _05308_);
  or (_05363_, _05361_, _00352_);
  or (_05364_, _05350_, _05308_);
  or (_05365_, _05364_, _00311_);
  and (_05367_, _05365_, _05363_);
  or (_05368_, _05347_, _05320_);
  or (_05369_, _05368_, _00188_);
  or (_05371_, _05350_, _05320_);
  or (_05372_, _05371_, _00116_);
  and (_05373_, _05372_, _05369_);
  and (_05375_, _05373_, _05367_);
  and (_05376_, _05375_, _05360_);
  and (_05377_, _05376_, _05345_);
  or (_05379_, _05310_, _00399_);
  or (_05380_, _05315_, _00358_);
  and (_05381_, _05380_, _05379_);
  or (_05383_, _05322_, _00235_);
  or (_05384_, _05324_, _00194_);
  and (_05385_, _05384_, _05383_);
  and (_05387_, _05385_, _05381_);
  or (_05388_, _05331_, _00576_);
  or (_05389_, _05334_, _00522_);
  and (_05391_, _05389_, _05388_);
  or (_05392_, _05339_, _00040_);
  or (_05393_, _05341_, _43809_);
  and (_05394_, _05393_, _05392_);
  and (_05395_, _05394_, _05391_);
  and (_05396_, _05395_, _05387_);
  or (_05397_, _05348_, _00481_);
  or (_05398_, _05351_, _00440_);
  and (_05399_, _05398_, _05397_);
  or (_05400_, _05354_, _43727_);
  or (_05401_, _05356_, _43768_);
  and (_05402_, _05401_, _05400_);
  and (_05403_, _05402_, _05399_);
  or (_05404_, _05361_, _00317_);
  or (_05405_, _05364_, _00276_);
  and (_05406_, _05405_, _05404_);
  or (_05407_, _05368_, _00122_);
  or (_05408_, _05371_, _00081_);
  and (_05409_, _05408_, _05407_);
  and (_05410_, _05409_, _05406_);
  and (_05411_, _05410_, _05403_);
  and (_05413_, _05411_, _05396_);
  and (_05414_, _05413_, _05377_);
  or (_05416_, _05310_, _00424_);
  or (_05417_, _05315_, _00383_);
  and (_05418_, _05417_, _05416_);
  or (_05420_, _05322_, _00260_);
  or (_05421_, _05324_, _00219_);
  and (_05422_, _05421_, _05420_);
  and (_05424_, _05422_, _05418_);
  or (_05425_, _05331_, _00607_);
  or (_05426_, _05334_, _00550_);
  and (_05428_, _05426_, _05425_);
  or (_05429_, _05339_, _00065_);
  or (_05430_, _05341_, _00024_);
  and (_05432_, _05430_, _05429_);
  and (_05433_, _05432_, _05428_);
  and (_05434_, _05433_, _05424_);
  or (_05436_, _05348_, _00506_);
  or (_05437_, _05351_, _00465_);
  and (_05438_, _05437_, _05436_);
  or (_05440_, _05354_, _43752_);
  or (_05441_, _05356_, _43793_);
  and (_05442_, _05441_, _05440_);
  and (_05444_, _05442_, _05438_);
  or (_05445_, _05361_, _00342_);
  or (_05446_, _05364_, _00301_);
  and (_05447_, _05446_, _05445_);
  or (_05448_, _05368_, _00168_);
  or (_05449_, _05371_, _00106_);
  and (_05450_, _05449_, _05448_);
  and (_05451_, _05450_, _05447_);
  and (_05452_, _05451_, _05444_);
  nand (_05453_, _05452_, _05434_);
  or (_05454_, _05310_, _00429_);
  or (_05455_, _05315_, _00388_);
  and (_05456_, _05455_, _05454_);
  or (_05457_, _05322_, _00265_);
  or (_05458_, _05324_, _00224_);
  and (_05459_, _05458_, _05457_);
  and (_05460_, _05459_, _05456_);
  or (_05461_, _05331_, _00612_);
  or (_05462_, _05334_, _00558_);
  and (_05463_, _05462_, _05461_);
  or (_05464_, _05339_, _00070_);
  or (_05466_, _05341_, _00029_);
  and (_05467_, _05466_, _05464_);
  and (_05469_, _05467_, _05463_);
  and (_05470_, _05469_, _05460_);
  or (_05471_, _05348_, _00511_);
  or (_05473_, _05351_, _00470_);
  and (_05474_, _05473_, _05471_);
  or (_05475_, _05354_, _43757_);
  or (_05477_, _05356_, _43798_);
  and (_05478_, _05477_, _05475_);
  and (_05479_, _05478_, _05474_);
  or (_05481_, _05361_, _00347_);
  or (_05482_, _05364_, _00306_);
  and (_05483_, _05482_, _05481_);
  or (_05485_, _05368_, _00179_);
  or (_05486_, _05371_, _00111_);
  and (_05487_, _05486_, _05485_);
  and (_05489_, _05487_, _05483_);
  and (_05490_, _05489_, _05479_);
  and (_05491_, _05490_, _05470_);
  nand (_05493_, _05491_, _05453_);
  not (_05494_, _05493_);
  and (_05495_, _05494_, _05414_);
  or (_05497_, _05310_, _00414_);
  or (_05498_, _05315_, _00373_);
  and (_05499_, _05498_, _05497_);
  or (_05500_, _05322_, _00250_);
  or (_05501_, _05324_, _00209_);
  and (_05502_, _05501_, _05500_);
  and (_05503_, _05502_, _05499_);
  or (_05504_, _05331_, _00597_);
  or (_05505_, _05334_, _00537_);
  and (_05506_, _05505_, _05504_);
  or (_05507_, _05339_, _00055_);
  or (_05508_, _05341_, _00014_);
  and (_05509_, _05508_, _05507_);
  and (_05510_, _05509_, _05506_);
  and (_05511_, _05510_, _05503_);
  or (_05512_, _05348_, _00496_);
  or (_05513_, _05351_, _00455_);
  and (_05514_, _05513_, _05512_);
  or (_05515_, _05354_, _43742_);
  or (_05516_, _05356_, _43783_);
  and (_05517_, _05516_, _05515_);
  and (_05519_, _05517_, _05514_);
  or (_05520_, _05361_, _00332_);
  or (_05522_, _05364_, _00291_);
  and (_05523_, _05522_, _05520_);
  or (_05524_, _05368_, _00146_);
  or (_05526_, _05371_, _00096_);
  and (_05527_, _05526_, _05524_);
  and (_05528_, _05527_, _05523_);
  and (_05530_, _05528_, _05519_);
  nand (_05531_, _05530_, _05511_);
  or (_05532_, _05310_, _00419_);
  or (_05534_, _05315_, _00378_);
  and (_05535_, _05534_, _05532_);
  or (_05536_, _05322_, _00255_);
  or (_05538_, _05324_, _00214_);
  and (_05539_, _05538_, _05536_);
  and (_05540_, _05539_, _05535_);
  or (_05542_, _05331_, _00602_);
  or (_05543_, _05334_, _00542_);
  and (_05544_, _05543_, _05542_);
  or (_05546_, _05339_, _00060_);
  or (_05547_, _05341_, _00019_);
  and (_05548_, _05547_, _05546_);
  and (_05550_, _05548_, _05544_);
  and (_05551_, _05550_, _05540_);
  or (_05552_, _05348_, _00501_);
  or (_05553_, _05351_, _00460_);
  and (_05554_, _05553_, _05552_);
  or (_05555_, _05354_, _43747_);
  or (_05556_, _05356_, _43788_);
  and (_05557_, _05556_, _05555_);
  and (_05558_, _05557_, _05554_);
  or (_05559_, _05361_, _00337_);
  or (_05560_, _05364_, _00296_);
  and (_05561_, _05560_, _05559_);
  or (_05562_, _05368_, _00157_);
  or (_05563_, _05371_, _00101_);
  and (_05564_, _05563_, _05562_);
  and (_05565_, _05564_, _05561_);
  and (_05566_, _05565_, _05558_);
  nand (_05567_, _05566_, _05551_);
  or (_05568_, _05567_, _05531_);
  not (_05569_, _05568_);
  or (_05570_, _05310_, _00409_);
  or (_05572_, _05315_, _00368_);
  and (_05573_, _05572_, _05570_);
  or (_05575_, _05322_, _00245_);
  or (_05576_, _05324_, _00204_);
  and (_05577_, _05576_, _05575_);
  and (_05579_, _05577_, _05573_);
  or (_05580_, _05331_, _00592_);
  or (_05581_, _05334_, _00532_);
  and (_05583_, _05581_, _05580_);
  or (_05584_, _05339_, _00050_);
  or (_05585_, _05341_, _00009_);
  and (_05587_, _05585_, _05584_);
  and (_05588_, _05587_, _05583_);
  and (_05589_, _05588_, _05579_);
  or (_05591_, _05348_, _00491_);
  or (_05592_, _05351_, _00450_);
  and (_05593_, _05592_, _05591_);
  or (_05595_, _05354_, _43737_);
  or (_05596_, _05356_, _43778_);
  and (_05597_, _05596_, _05595_);
  and (_05599_, _05597_, _05593_);
  or (_05600_, _05361_, _00327_);
  or (_05601_, _05364_, _00286_);
  and (_05603_, _05601_, _05600_);
  or (_05604_, _05368_, _00135_);
  or (_05605_, _05371_, _00091_);
  and (_05606_, _05605_, _05604_);
  and (_05607_, _05606_, _05603_);
  and (_05608_, _05607_, _05599_);
  nand (_05609_, _05608_, _05589_);
  not (_05610_, _05609_);
  or (_05611_, _05310_, _00404_);
  or (_05612_, _05315_, _00363_);
  and (_05613_, _05612_, _05611_);
  or (_05614_, _05322_, _00240_);
  or (_05615_, _05324_, _00199_);
  and (_05616_, _05615_, _05614_);
  and (_05617_, _05616_, _05613_);
  or (_05618_, _05331_, _00584_);
  or (_05619_, _05334_, _00527_);
  and (_05620_, _05619_, _05618_);
  or (_05621_, _05339_, _00045_);
  or (_05622_, _05341_, _00004_);
  and (_05623_, _05622_, _05621_);
  and (_05625_, _05623_, _05620_);
  and (_05626_, _05625_, _05617_);
  or (_05628_, _05348_, _00486_);
  or (_05629_, _05351_, _00445_);
  and (_05630_, _05629_, _05628_);
  or (_05632_, _05354_, _43732_);
  or (_05633_, _05356_, _43773_);
  and (_05634_, _05633_, _05632_);
  and (_05636_, _05634_, _05630_);
  or (_05637_, _05361_, _00322_);
  or (_05638_, _05364_, _00281_);
  and (_05640_, _05638_, _05637_);
  or (_05641_, _05368_, _00127_);
  or (_05642_, _05371_, _00086_);
  and (_05644_, _05642_, _05641_);
  and (_05645_, _05644_, _05640_);
  and (_05646_, _05645_, _05636_);
  and (_05648_, _05646_, _05626_);
  and (_05649_, _05648_, _05610_);
  and (_05650_, _05649_, _05569_);
  and (_05652_, _05650_, _05495_);
  not (_05653_, _05652_);
  and (_05654_, _05452_, _05434_);
  nand (_05656_, _05491_, _05654_);
  nand (_05657_, _05376_, _05345_);
  or (_05658_, _05413_, _05657_);
  nor (_05659_, _05658_, _05656_);
  not (_05660_, _05659_);
  or (_05661_, _05648_, _05610_);
  or (_05662_, _05661_, _05568_);
  nor (_05663_, _05662_, _05660_);
  not (_05664_, _05663_);
  or (_05665_, _05648_, _05609_);
  not (_05666_, _05531_);
  or (_05667_, _05567_, _05666_);
  or (_05668_, _05667_, _05665_);
  or (_05669_, _05668_, _05660_);
  or (_05670_, _05665_, _05568_);
  nor (_05671_, _05658_, _05493_);
  not (_05672_, _05671_);
  or (_05673_, _05672_, _05670_);
  and (_05674_, _05673_, _05669_);
  or (_05675_, _05672_, _05662_);
  not (_05676_, _05675_);
  and (_05678_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_05679_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_05681_, _05679_, _05678_);
  nand (_05682_, _05681_, _05676_);
  or (_05683_, _05491_, _05654_);
  or (_05685_, _05683_, _05658_);
  or (_05686_, _05685_, _05670_);
  or (_05687_, _05413_, _05377_);
  or (_05689_, _05687_, _05493_);
  or (_05690_, _05689_, _05670_);
  and (_05691_, _05690_, _05686_);
  or (_05693_, _05687_, _05656_);
  or (_05694_, _05693_, _05670_);
  or (_05695_, _05491_, _05453_);
  or (_05697_, _05695_, _05687_);
  or (_05698_, _05697_, _05670_);
  and (_05699_, _05698_, _05694_);
  or (_05701_, _05695_, _05658_);
  or (_05702_, _05701_, _05670_);
  or (_05703_, _05687_, _05683_);
  or (_05705_, _05703_, _05670_);
  and (_05706_, _05705_, _05702_);
  and (_05707_, _05706_, _05699_);
  and (_05709_, _05707_, _05691_);
  and (_05710_, _05675_, _05346_);
  nand (_05711_, _05710_, _05709_);
  nand (_05712_, _05711_, _05682_);
  nand (_05713_, _05712_, _05674_);
  and (_05714_, _05709_, _05674_);
  or (_05715_, _05714_, _05346_);
  nand (_05716_, _05715_, _05713_);
  nand (_05717_, _05716_, _05664_);
  not (_05718_, _05670_);
  and (_05719_, _05718_, _05659_);
  not (_05720_, _05719_);
  not (_05721_, _05683_);
  and (_05722_, _05413_, _05657_);
  and (_05723_, _05722_, _05721_);
  and (_05724_, _05723_, _05718_);
  not (_05725_, _05695_);
  and (_05726_, _05722_, _05725_);
  and (_05727_, _05726_, _05718_);
  nor (_05728_, _05727_, _05724_);
  and (_05729_, _05728_, _05720_);
  and (_05731_, _05721_, _05414_);
  and (_05732_, _05731_, _05718_);
  not (_05734_, _05732_);
  and (_05735_, _05722_, _05494_);
  and (_05736_, _05735_, _05718_);
  not (_05738_, _05656_);
  and (_05739_, _05722_, _05738_);
  and (_05740_, _05739_, _05718_);
  nor (_05742_, _05740_, _05736_);
  and (_05743_, _05742_, _05734_);
  and (_05744_, _05743_, _05729_);
  and (_05746_, _05725_, _05414_);
  and (_05747_, _05746_, _05718_);
  not (_05748_, _05747_);
  and (_05750_, _05738_, _05414_);
  and (_05751_, _05750_, _05718_);
  and (_05752_, _05718_, _05495_);
  nor (_05754_, _05752_, _05751_);
  and (_05755_, _05754_, _05748_);
  and (_05756_, _05755_, _05744_);
  not (_05758_, \oc8051_golden_model_1.ACC [0]);
  and (_05759_, _05758_, \oc8051_golden_model_1.PC [0]);
  and (_05760_, \oc8051_golden_model_1.ACC [0], _05346_);
  or (_05762_, _05760_, _05664_);
  or (_05763_, _05762_, _05759_);
  and (_05764_, _05763_, _05756_);
  nand (_05765_, _05764_, _05717_);
  or (_05766_, _05756_, \oc8051_golden_model_1.PC [0]);
  and (_05767_, _05766_, _05765_);
  and (_05768_, _05756_, _05714_);
  or (_05769_, _05768_, _05312_);
  and (_05770_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_05771_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_05772_, _05771_, _05770_);
  and (_05773_, _05772_, _05678_);
  nor (_05774_, _05772_, _05678_);
  nor (_05775_, _05774_, _05773_);
  or (_05776_, _05775_, _05675_);
  and (_05777_, _05347_, _05314_);
  and (_05778_, _05777_, _05675_);
  nand (_05779_, _05778_, _05709_);
  nand (_05780_, _05779_, _05776_);
  and (_05781_, _05674_, _05664_);
  and (_05782_, _05781_, _05780_);
  not (_05784_, \oc8051_golden_model_1.ACC [1]);
  nor (_05785_, _05777_, _05784_);
  and (_05787_, _05777_, _05784_);
  nor (_05788_, _05787_, _05785_);
  and (_05789_, _05788_, _05760_);
  nor (_05791_, _05788_, _05760_);
  nor (_05792_, _05791_, _05789_);
  nor (_05793_, _05792_, _05664_);
  or (_05795_, _05793_, _05782_);
  nand (_05796_, _05795_, _05756_);
  nand (_05797_, _05796_, _05769_);
  or (_05799_, _05797_, _05767_);
  and (_05800_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_05801_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_05803_, _05801_, _05800_);
  not (_05804_, _05803_);
  nor (_05805_, _05804_, _05755_);
  not (_05807_, _05805_);
  nor (_05808_, _05773_, _05770_);
  and (_05809_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_05811_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_05812_, _05811_, _05809_);
  not (_05813_, _05812_);
  nor (_05815_, _05813_, _05808_);
  and (_05816_, _05813_, _05808_);
  nor (_05817_, _05816_, _05815_);
  not (_05818_, _05817_);
  or (_05819_, _05818_, _05675_);
  and (_05820_, _05819_, _05674_);
  nor (_05821_, _05305_, _05319_);
  and (_05822_, _05305_, _05319_);
  nor (_05823_, _05822_, _05821_);
  not (_05824_, _05823_);
  nand (_05825_, _05824_, _05709_);
  nand (_05826_, _05825_, _05675_);
  nand (_05827_, _05826_, _05820_);
  or (_05828_, _05803_, _05714_);
  and (_05829_, _05828_, _05664_);
  nand (_05830_, _05829_, _05827_);
  nor (_05831_, _05789_, _05785_);
  and (_05832_, _05823_, \oc8051_golden_model_1.ACC [2]);
  nor (_05833_, _05823_, \oc8051_golden_model_1.ACC [2]);
  nor (_05834_, _05833_, _05832_);
  not (_05835_, _05834_);
  and (_05837_, _05835_, _05831_);
  nor (_05838_, _05835_, _05831_);
  nor (_05840_, _05838_, _05837_);
  and (_05841_, _05840_, _05663_);
  not (_05842_, _05841_);
  and (_05844_, _05842_, _05744_);
  nand (_05845_, _05844_, _05830_);
  or (_05846_, _05803_, _05756_);
  nand (_05848_, _05846_, _05845_);
  and (_05849_, _05848_, _05807_);
  nor (_05850_, _05330_, _05312_);
  nor (_05852_, _05800_, \oc8051_golden_model_1.PC [3]);
  nor (_05853_, _05852_, _05850_);
  or (_05854_, _05853_, _05768_);
  nor (_05856_, _05815_, _05809_);
  and (_05857_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_05858_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_05860_, _05858_, _05857_);
  not (_05861_, _05860_);
  nor (_05862_, _05861_, _05856_);
  and (_05864_, _05861_, _05856_);
  nor (_05865_, _05864_, _05862_);
  or (_05866_, _05865_, _05675_);
  not (_05868_, _05322_);
  nor (_05869_, _05821_, _05307_);
  nor (_05870_, _05869_, _05868_);
  and (_05871_, _05675_, _05870_);
  nand (_05872_, _05871_, _05709_);
  nand (_05873_, _05872_, _05866_);
  and (_05874_, _05873_, _05781_);
  nor (_05875_, _05838_, _05832_);
  nor (_05876_, _05870_, \oc8051_golden_model_1.ACC [3]);
  and (_05877_, _05870_, \oc8051_golden_model_1.ACC [3]);
  nor (_05878_, _05877_, _05876_);
  and (_05879_, _05878_, _05875_);
  nor (_05880_, _05878_, _05875_);
  nor (_05881_, _05880_, _05879_);
  nor (_05882_, _05881_, _05664_);
  or (_05883_, _05882_, _05874_);
  nand (_05884_, _05883_, _05756_);
  and (_05885_, _05884_, _05854_);
  or (_05886_, _05885_, _05849_);
  or (_05887_, _05886_, _05799_);
  or (_05888_, _05887_, _00194_);
  nand (_05890_, _05766_, _05765_);
  and (_05891_, _05796_, _05769_);
  or (_05893_, _05891_, _05890_);
  or (_05894_, _05893_, _05886_);
  or (_05895_, _05894_, _00122_);
  and (_05897_, _05895_, _05888_);
  nand (_05898_, _05884_, _05854_);
  or (_05899_, _05898_, _05849_);
  or (_05901_, _05797_, _05890_);
  or (_05902_, _05901_, _05899_);
  or (_05903_, _05902_, _00576_);
  nand (_05905_, _05848_, _05807_);
  or (_05906_, _05898_, _05905_);
  or (_05907_, _05906_, _05901_);
  or (_05909_, _05907_, _00399_);
  and (_05910_, _05909_, _05903_);
  and (_05911_, _05910_, _05897_);
  or (_05913_, _05906_, _05799_);
  or (_05914_, _05913_, _00358_);
  or (_05915_, _05906_, _05893_);
  or (_05917_, _05915_, _00317_);
  and (_05918_, _05917_, _05914_);
  or (_05919_, _05899_, _05893_);
  or (_05921_, _05919_, _00481_);
  or (_05922_, _05891_, _05767_);
  or (_05923_, _05922_, _05899_);
  or (_05924_, _05923_, _00440_);
  and (_05925_, _05924_, _05921_);
  and (_05926_, _05925_, _05918_);
  and (_05927_, _05926_, _05911_);
  or (_05928_, _05885_, _05905_);
  or (_05929_, _05928_, _05922_);
  or (_05930_, _05929_, _43727_);
  or (_05931_, _05928_, _05799_);
  or (_05932_, _05931_, _43809_);
  and (_05933_, _05932_, _05930_);
  or (_05934_, _05901_, _05886_);
  or (_05935_, _05934_, _00235_);
  or (_05936_, _05922_, _05886_);
  or (_05937_, _05936_, _00081_);
  and (_05938_, _05937_, _05935_);
  and (_05939_, _05938_, _05933_);
  or (_05940_, _05899_, _05799_);
  or (_05941_, _05940_, _00522_);
  or (_05942_, _05906_, _05922_);
  or (_05943_, _05942_, _00276_);
  and (_05944_, _05943_, _05941_);
  or (_05945_, _05928_, _05901_);
  or (_05946_, _05945_, _00040_);
  or (_05947_, _05928_, _05893_);
  or (_05948_, _05947_, _43768_);
  and (_05949_, _05948_, _05946_);
  and (_05950_, _05949_, _05944_);
  and (_05951_, _05950_, _05939_);
  nand (_05952_, _05951_, _05927_);
  or (_05953_, _05907_, _00419_);
  or (_05954_, _05929_, _43747_);
  and (_05955_, _05954_, _05953_);
  or (_05956_, _05919_, _00501_);
  or (_05957_, _05887_, _00214_);
  and (_05958_, _05957_, _05956_);
  and (_05959_, _05958_, _05955_);
  or (_05960_, _05913_, _00378_);
  or (_05961_, _05915_, _00337_);
  and (_05962_, _05961_, _05960_);
  or (_05963_, _05940_, _00542_);
  or (_05964_, _05945_, _00060_);
  and (_05965_, _05964_, _05963_);
  and (_05966_, _05965_, _05962_);
  and (_05967_, _05966_, _05959_);
  or (_05968_, _05936_, _00101_);
  or (_05969_, _05947_, _43788_);
  and (_05970_, _05969_, _05968_);
  or (_05971_, _05934_, _00255_);
  or (_05972_, _05894_, _00157_);
  and (_05973_, _05972_, _05971_);
  and (_05974_, _05973_, _05970_);
  or (_05975_, _05942_, _00296_);
  or (_05976_, _05931_, _00019_);
  and (_05977_, _05976_, _05975_);
  or (_05978_, _05902_, _00602_);
  or (_05979_, _05923_, _00460_);
  and (_05980_, _05979_, _05978_);
  and (_05981_, _05980_, _05977_);
  and (_05982_, _05981_, _05974_);
  and (_05983_, _05982_, _05967_);
  or (_05984_, _05983_, _05952_);
  nor (_05985_, _05984_, _05653_);
  or (_05986_, _05945_, _00045_);
  or (_05987_, _05929_, _43732_);
  and (_05988_, _05987_, _05986_);
  or (_05989_, _05942_, _00281_);
  or (_05990_, _05931_, _00004_);
  and (_05991_, _05990_, _05989_);
  and (_05992_, _05991_, _05988_);
  or (_05993_, _05934_, _00240_);
  or (_05994_, _05887_, _00199_);
  and (_05995_, _05994_, _05993_);
  or (_05996_, _05902_, _00584_);
  or (_05997_, _05923_, _00445_);
  and (_05998_, _05997_, _05996_);
  and (_05999_, _05998_, _05995_);
  and (_06000_, _05999_, _05992_);
  or (_06001_, _05936_, _00086_);
  or (_06002_, _05947_, _43773_);
  and (_06003_, _06002_, _06001_);
  or (_06004_, _05907_, _00404_);
  or (_06005_, _05913_, _00363_);
  and (_06006_, _06005_, _06004_);
  and (_06007_, _06006_, _06003_);
  or (_06008_, _05940_, _00527_);
  or (_06009_, _05919_, _00486_);
  and (_06010_, _06009_, _06008_);
  or (_06011_, _05915_, _00322_);
  or (_06012_, _05894_, _00127_);
  and (_06013_, _06012_, _06011_);
  and (_06014_, _06013_, _06010_);
  and (_06015_, _06014_, _06007_);
  and (_06016_, _06015_, _06000_);
  not (_06017_, _06016_);
  not (_06018_, _05668_);
  and (_06019_, _05723_, _06018_);
  not (_06020_, _06019_);
  nor (_06021_, _06020_, _05952_);
  and (_06022_, _06021_, _06017_);
  not (_06023_, _05673_);
  and (_06024_, _05648_, _05609_);
  and (_06025_, _06024_, _05569_);
  and (_06026_, _06025_, _05671_);
  not (_06027_, _06026_);
  nor (_06028_, _06027_, _05984_);
  not (_06029_, \oc8051_golden_model_1.SP [0]);
  nor (_06030_, _05686_, _06029_);
  not (_06031_, _05685_);
  and (_06032_, _06025_, _06031_);
  not (_06033_, _06032_);
  nor (_06034_, _06033_, _05984_);
  nor (_06035_, _06033_, _05952_);
  not (_06036_, _06035_);
  not (_06037_, _05693_);
  and (_06038_, _06037_, _05650_);
  and (_06039_, _06025_, _06037_);
  not (_06040_, _06039_);
  nor (_06041_, _06040_, _05984_);
  not (_06042_, _05689_);
  and (_06043_, _06025_, _06042_);
  not (_06044_, _06043_);
  or (_06045_, _06044_, _05984_);
  not (_06046_, _05705_);
  and (_06047_, _05750_, _06018_);
  not (_06048_, _06047_);
  and (_06049_, _06025_, _05746_);
  not (_06050_, _06049_);
  and (_06051_, _05746_, _06018_);
  not (_06052_, _06051_);
  not (_06053_, _05952_);
  nor (_06054_, _05907_, _00434_);
  nor (_06055_, _05934_, _00270_);
  nor (_06056_, _06055_, _06054_);
  nor (_06057_, _05887_, _00229_);
  nor (_06058_, _05929_, _43762_);
  nor (_06059_, _06058_, _06057_);
  and (_06060_, _06059_, _06056_);
  nor (_06061_, _05919_, _00516_);
  nor (_06062_, _05940_, _00566_);
  nor (_06063_, _06062_, _06061_);
  nor (_06064_, _05902_, _00617_);
  nor (_06065_, _05945_, _00075_);
  nor (_06066_, _06065_, _06064_);
  and (_06067_, _06066_, _06063_);
  and (_06068_, _06067_, _06060_);
  nor (_06069_, _05894_, _00188_);
  nor (_06070_, _05936_, _00116_);
  nor (_06071_, _06070_, _06069_);
  nor (_06072_, _05923_, _00475_);
  nor (_06073_, _05947_, _43803_);
  nor (_06074_, _06073_, _06072_);
  and (_06075_, _06074_, _06071_);
  nor (_06076_, _05913_, _00393_);
  nor (_06077_, _05931_, _00034_);
  nor (_06078_, _06077_, _06076_);
  nor (_06079_, _05915_, _00352_);
  nor (_06080_, _05942_, _00311_);
  nor (_06081_, _06080_, _06079_);
  and (_06082_, _06081_, _06078_);
  and (_06083_, _06082_, _06075_);
  and (_06084_, _06083_, _06068_);
  and (_06085_, _06084_, _06053_);
  and (_06086_, _05983_, _05952_);
  nor (_06087_, _06086_, _06085_);
  and (_06088_, _06025_, _05723_);
  and (_06089_, _06025_, _05659_);
  nor (_06090_, _06089_, _06088_);
  nor (_06091_, _06090_, _06087_);
  not (_06092_, _05661_);
  and (_06093_, _05567_, _05531_);
  and (_06094_, _06093_, _06092_);
  and (_06095_, _05567_, _05666_);
  and (_06096_, _06095_, _05649_);
  not (_06097_, _05665_);
  and (_06098_, _06093_, _06097_);
  or (_06099_, _06098_, _06096_);
  nor (_06100_, _06099_, _06094_);
  or (_06101_, _06100_, _05685_);
  nor (_06102_, _05689_, _05668_);
  nor (_06103_, _05667_, _05610_);
  and (_06104_, _06103_, _06031_);
  nor (_06105_, _06104_, _06102_);
  and (_06106_, _06105_, _06101_);
  not (_06107_, _05662_);
  and (_06108_, _05735_, _06107_);
  nor (_06109_, _06108_, _06019_);
  and (_06110_, _05671_, _05650_);
  not (_06111_, _06110_);
  and (_06112_, _05726_, _06107_);
  not (_06113_, _05667_);
  and (_06114_, _06113_, _05649_);
  and (_06115_, _06114_, _06031_);
  nor (_06116_, _06115_, _06112_);
  and (_06117_, _06116_, _06111_);
  and (_06118_, _06117_, _06109_);
  and (_06119_, _06025_, _05750_);
  nor (_06120_, _06119_, _05652_);
  nor (_06121_, _05685_, _05668_);
  and (_06122_, _06093_, _06024_);
  and (_06123_, _06122_, _06031_);
  nor (_06124_, _06123_, _06121_);
  and (_06125_, _06124_, _06120_);
  and (_06126_, _05746_, _05650_);
  and (_06127_, _06025_, _05495_);
  nor (_06128_, _06127_, _06126_);
  and (_06129_, _05731_, _05650_);
  and (_06130_, _05739_, _06107_);
  nor (_06131_, _06130_, _06129_);
  and (_06132_, _06131_, _06128_);
  and (_06133_, _06095_, _06097_);
  and (_06134_, _06133_, _06031_);
  and (_06135_, _06095_, _05609_);
  and (_06136_, _06093_, _05649_);
  nor (_06137_, _06136_, _06135_);
  nor (_06138_, _06137_, _05685_);
  or (_06139_, _06138_, _06134_);
  not (_06140_, _06139_);
  and (_06141_, _06140_, _06132_);
  and (_06142_, _06141_, _06125_);
  and (_06143_, _06142_, _06118_);
  and (_06144_, _06143_, _06106_);
  nor (_06145_, _06144_, _05803_);
  and (_06146_, _06144_, _05824_);
  nor (_06147_, _06146_, _06145_);
  not (_06148_, _05853_);
  nor (_06149_, _06144_, _06148_);
  not (_06150_, _05870_);
  and (_06151_, _06144_, _06150_);
  nor (_06152_, _06151_, _06149_);
  nor (_06153_, _06152_, _06147_);
  and (_06154_, _06144_, _05346_);
  nor (_06155_, _06154_, \oc8051_golden_model_1.PC [1]);
  and (_06156_, _06154_, \oc8051_golden_model_1.PC [1]);
  nor (_06157_, _06156_, _06155_);
  nor (_06158_, _06144_, _05346_);
  nor (_06159_, _06158_, _06154_);
  nor (_06160_, _06159_, _06157_);
  and (_06161_, _06160_, _06153_);
  and (_06162_, _06161_, _04446_);
  and (_06163_, _06159_, _06157_);
  not (_06164_, _06152_);
  nor (_06165_, _06164_, _06147_);
  and (_06166_, _06165_, _06163_);
  and (_06167_, _06166_, _04486_);
  nor (_06168_, _06167_, _06162_);
  and (_06169_, _06164_, _06147_);
  and (_06170_, _06169_, _06160_);
  and (_06171_, _06170_, _04462_);
  not (_06172_, _06159_);
  nor (_06173_, _06172_, _06157_);
  and (_06174_, _06152_, _06147_);
  and (_06175_, _06174_, _06173_);
  and (_06176_, _06175_, _04473_);
  nor (_06177_, _06176_, _06171_);
  and (_06178_, _06177_, _06168_);
  and (_06179_, _06173_, _06153_);
  and (_06180_, _06179_, _04477_);
  and (_06181_, _06172_, _06157_);
  and (_06182_, _06181_, _06153_);
  and (_06183_, _06182_, _04464_);
  nor (_06184_, _06183_, _06180_);
  and (_06185_, _06173_, _06169_);
  and (_06186_, _06185_, _04467_);
  and (_06187_, _06165_, _06160_);
  and (_06188_, _06187_, _04457_);
  nor (_06189_, _06188_, _06186_);
  and (_06190_, _06189_, _06184_);
  and (_06191_, _06190_, _06178_);
  and (_06192_, _06174_, _06163_);
  and (_06193_, _06192_, _04459_);
  and (_06194_, _06181_, _06165_);
  and (_06195_, _06194_, _04475_);
  nor (_06196_, _06195_, _06193_);
  and (_06197_, _06174_, _06160_);
  and (_06198_, _06197_, _04469_);
  and (_06199_, _06174_, _06181_);
  and (_06200_, _06199_, _04448_);
  nor (_06201_, _06200_, _06198_);
  and (_06202_, _06201_, _06196_);
  and (_06203_, _06163_, _06153_);
  and (_06204_, _06203_, _04484_);
  and (_06205_, _06173_, _06165_);
  and (_06206_, _06205_, _04479_);
  nor (_06207_, _06206_, _06204_);
  and (_06208_, _06181_, _06169_);
  and (_06209_, _06208_, _04453_);
  and (_06210_, _06169_, _06163_);
  and (_06211_, _06210_, _04451_);
  nor (_06212_, _06211_, _06209_);
  and (_06213_, _06212_, _06207_);
  and (_06214_, _06213_, _06202_);
  and (_06215_, _06214_, _06191_);
  nor (_06216_, _06215_, _05669_);
  not (_06217_, _06090_);
  nor (_06218_, _06121_, _06038_);
  nor (_06219_, _05693_, _05668_);
  not (_06220_, _06219_);
  not (_06221_, _05701_);
  and (_06222_, _06093_, _06221_);
  not (_06223_, _06222_);
  and (_06224_, _06096_, _06221_);
  and (_06225_, _06133_, _06221_);
  nor (_06226_, _06225_, _06224_);
  and (_06227_, _06095_, _06024_);
  and (_06228_, _06227_, _06221_);
  and (_06229_, _06095_, _06092_);
  and (_06230_, _06229_, _06221_);
  nor (_06231_, _06230_, _06228_);
  and (_06232_, _06231_, _06226_);
  and (_06233_, _06232_, _06223_);
  and (_06234_, _06233_, _06220_);
  and (_06235_, _06234_, _06218_);
  or (_06236_, _06235_, _05983_);
  nor (_06237_, _06044_, _06087_);
  not (_06238_, \oc8051_golden_model_1.SP [3]);
  and (_06239_, _06042_, _05650_);
  and (_06240_, _06239_, _06238_);
  nor (_06241_, _05697_, _05668_);
  nor (_06242_, _06241_, _06102_);
  or (_06243_, _06242_, _05983_);
  nor (_06244_, _06239_, _06043_);
  nand (_06245_, _06242_, \oc8051_golden_model_1.PSW [3]);
  and (_06246_, _06245_, _06244_);
  or (_06247_, _06246_, _06219_);
  and (_06248_, _06247_, _06243_);
  or (_06249_, _06248_, _06240_);
  and (_06250_, _06221_, _05650_);
  and (_06251_, _06025_, _06221_);
  nor (_06252_, _06251_, _06250_);
  and (_06253_, _06031_, _05650_);
  nor (_06254_, _06032_, _06253_);
  and (_06255_, _06254_, _06040_);
  and (_06256_, _06255_, _06252_);
  and (_06257_, _06256_, _06249_);
  or (_06258_, _06257_, _06237_);
  and (_06259_, _06258_, _06236_);
  nor (_06260_, _06256_, _06087_);
  nor (_06261_, _05672_, _05668_);
  nand (_06262_, _06233_, _06218_);
  and (_06263_, _06262_, _05983_);
  or (_06264_, _06263_, _06261_);
  or (_06265_, _06264_, _06260_);
  nor (_06266_, _06265_, _06259_);
  not (_06267_, _06261_);
  nor (_06268_, _06267_, _05983_);
  or (_06269_, _06268_, _06266_);
  and (_06270_, _06269_, _06027_);
  and (_06271_, _06087_, _06026_);
  or (_06272_, _06271_, _06270_);
  and (_06273_, _06272_, _05669_);
  or (_06274_, _06273_, _06217_);
  nor (_06275_, _06274_, _06216_);
  or (_06276_, _06275_, _06091_);
  and (_06277_, _06025_, _05735_);
  not (_06278_, _06277_);
  and (_06279_, _05735_, _06018_);
  nor (_06280_, _06279_, _06108_);
  and (_06281_, _06280_, _06278_);
  and (_06282_, _05726_, _06018_);
  not (_06283_, _06282_);
  and (_06284_, _06025_, _05726_);
  nor (_06285_, _06284_, _06112_);
  and (_06286_, _06285_, _06283_);
  and (_06287_, _06286_, _06281_);
  and (_06288_, _05731_, _06018_);
  not (_06289_, _06288_);
  and (_06290_, _05739_, _06018_);
  not (_06291_, _06290_);
  and (_06292_, _06025_, _05739_);
  nor (_06293_, _06292_, _06130_);
  and (_06294_, _06293_, _06291_);
  and (_06295_, _06294_, _06289_);
  and (_06296_, _06295_, _06287_);
  nand (_06297_, _06296_, _06276_);
  and (_06298_, _06025_, _05731_);
  not (_06299_, _05983_);
  nor (_06300_, _06296_, _06299_);
  nor (_06301_, _06300_, _06298_);
  and (_06302_, _06301_, _06297_);
  and (_06303_, _06298_, \oc8051_golden_model_1.SP [3]);
  or (_06304_, _06303_, _06129_);
  nor (_06305_, _06304_, _06302_);
  not (_06306_, _06129_);
  nor (_06307_, _06087_, _06306_);
  or (_06308_, _06307_, _06305_);
  and (_06309_, _06308_, _06052_);
  and (_06310_, _06051_, _05983_);
  or (_06311_, _06310_, _06309_);
  nand (_06312_, _06311_, _06050_);
  and (_06313_, _06049_, _06238_);
  nor (_06314_, _06313_, _06126_);
  nand (_06315_, _06314_, _06312_);
  and (_06316_, _06018_, _05495_);
  and (_06317_, _06126_, _06087_);
  nor (_06318_, _06317_, _06316_);
  nand (_06319_, _06318_, _06315_);
  and (_06320_, _06316_, _05983_);
  nor (_06321_, _06320_, _05652_);
  and (_06322_, _06321_, _06319_);
  and (_06323_, _06087_, _05652_);
  or (_06324_, _06323_, _06322_);
  nand (_06325_, _06324_, _06048_);
  nor (_06326_, _06048_, _05983_);
  not (_06327_, _06326_);
  and (_06328_, _06327_, _06325_);
  nor (_06329_, _05902_, _00612_);
  nor (_06330_, _05915_, _00347_);
  nor (_06331_, _06330_, _06329_);
  nor (_06332_, _05913_, _00388_);
  nor (_06333_, _05945_, _00070_);
  nor (_06334_, _06333_, _06332_);
  and (_06335_, _06334_, _06331_);
  nor (_06336_, _05934_, _00265_);
  nor (_06337_, _05894_, _00179_);
  nor (_06338_, _06337_, _06336_);
  nor (_06339_, _05940_, _00558_);
  nor (_06340_, _05923_, _00470_);
  nor (_06341_, _06340_, _06339_);
  and (_06342_, _06341_, _06338_);
  and (_06343_, _06342_, _06335_);
  nor (_06344_, _05936_, _00111_);
  nor (_06345_, _05931_, _00029_);
  nor (_06346_, _06345_, _06344_);
  nor (_06347_, _05929_, _43757_);
  nor (_06348_, _05947_, _43798_);
  nor (_06349_, _06348_, _06347_);
  and (_06350_, _06349_, _06346_);
  nor (_06351_, _05919_, _00511_);
  nor (_06352_, _05887_, _00224_);
  nor (_06353_, _06352_, _06351_);
  nor (_06354_, _05907_, _00429_);
  nor (_06355_, _05942_, _00306_);
  nor (_06356_, _06355_, _06354_);
  and (_06357_, _06356_, _06353_);
  and (_06358_, _06357_, _06350_);
  and (_06359_, _06358_, _06343_);
  nor (_06360_, _06359_, _05952_);
  not (_06361_, _06360_);
  and (_06362_, _06254_, _06252_);
  nor (_06363_, _06126_, _06043_);
  and (_06364_, _06363_, _06306_);
  nor (_06365_, _06026_, _05652_);
  and (_06366_, _06365_, _06090_);
  and (_06367_, _06366_, _06364_);
  and (_06368_, _06367_, _06362_);
  nor (_06369_, _06368_, _06361_);
  not (_06370_, _06369_);
  and (_06371_, _06360_, _06039_);
  not (_06372_, _06371_);
  nor (_06373_, _05915_, _00332_);
  nor (_06374_, _05936_, _00096_);
  nor (_06375_, _06374_, _06373_);
  nor (_06376_, _05902_, _00597_);
  nor (_06377_, _05934_, _00250_);
  nor (_06378_, _06377_, _06376_);
  and (_06379_, _06378_, _06375_);
  nor (_06380_, _05942_, _00291_);
  nor (_06381_, _05894_, _00146_);
  nor (_06382_, _06381_, _06380_);
  nor (_06383_, _05929_, _43742_);
  nor (_06384_, _05947_, _43783_);
  nor (_06385_, _06384_, _06383_);
  and (_06386_, _06385_, _06382_);
  and (_06387_, _06386_, _06379_);
  nor (_06388_, _05919_, _00496_);
  nor (_06389_, _05913_, _00373_);
  nor (_06390_, _06389_, _06388_);
  nor (_06391_, _05887_, _00209_);
  nor (_06392_, _05931_, _00014_);
  nor (_06393_, _06392_, _06391_);
  and (_06394_, _06393_, _06390_);
  nor (_06395_, _05907_, _00414_);
  nor (_06396_, _05923_, _00455_);
  nor (_06397_, _06396_, _06395_);
  nor (_06398_, _05940_, _00537_);
  nor (_06399_, _05945_, _00055_);
  nor (_06400_, _06399_, _06398_);
  and (_06401_, _06400_, _06397_);
  and (_06402_, _06401_, _06394_);
  and (_06403_, _06402_, _06387_);
  nor (_06404_, _06288_, _06261_);
  and (_06405_, _06404_, _06218_);
  and (_06406_, _06405_, _06242_);
  and (_06407_, _06406_, _06234_);
  nor (_06408_, _06316_, _06047_);
  and (_06409_, _06408_, _06052_);
  and (_06410_, _06409_, _06294_);
  and (_06411_, _06410_, _06287_);
  and (_06412_, _06411_, _06407_);
  nor (_06413_, _06412_, _06403_);
  not (_06414_, _06413_);
  and (_06415_, _06170_, _04437_);
  and (_06416_, _06161_, _04406_);
  nor (_06417_, _06416_, _06415_);
  and (_06418_, _06192_, _04410_);
  and (_06419_, _06166_, _04417_);
  nor (_06420_, _06419_, _06418_);
  and (_06421_, _06420_, _06417_);
  and (_06422_, _06185_, _04415_);
  and (_06423_, _06210_, _04399_);
  nor (_06424_, _06423_, _06422_);
  and (_06425_, _06179_, _04428_);
  and (_06426_, _06203_, _04439_);
  nor (_06427_, _06426_, _06425_);
  and (_06428_, _06427_, _06424_);
  and (_06429_, _06428_, _06421_);
  and (_06430_, _06197_, _04422_);
  and (_06431_, _06175_, _04426_);
  nor (_06432_, _06431_, _06430_);
  and (_06433_, _06199_, _04401_);
  and (_06434_, _06187_, _04412_);
  nor (_06435_, _06434_, _06433_);
  and (_06436_, _06435_, _06432_);
  and (_06437_, _06205_, _04432_);
  and (_06438_, _06194_, _04430_);
  nor (_06439_, _06438_, _06437_);
  and (_06440_, _06208_, _04404_);
  and (_06441_, _06182_, _04420_);
  nor (_06442_, _06441_, _06440_);
  and (_06443_, _06442_, _06439_);
  and (_06444_, _06443_, _06436_);
  and (_06445_, _06444_, _06429_);
  nor (_06446_, _06445_, _05669_);
  not (_06447_, \oc8051_golden_model_1.SP [2]);
  nor (_06448_, _06298_, _06049_);
  nor (_06449_, _06448_, _06447_);
  and (_06450_, _06093_, _05609_);
  not (_06451_, _06450_);
  and (_06452_, _05453_, _05414_);
  or (_06453_, _06037_, _05659_);
  nor (_06454_, _06453_, _06452_);
  nor (_06455_, _06454_, _06451_);
  nor (_06456_, _06455_, _06449_);
  and (_06457_, _06136_, _05495_);
  and (_06458_, _06098_, _05495_);
  nor (_06459_, _06458_, _06457_);
  and (_06460_, _06093_, _05610_);
  and (_06461_, _06460_, _06042_);
  not (_06462_, _06461_);
  and (_06463_, _06460_, _06037_);
  and (_06464_, _06093_, _05750_);
  nor (_06465_, _06464_, _06463_);
  and (_06466_, _06465_, _06462_);
  and (_06467_, _06466_, _06459_);
  and (_06468_, _06467_, _06456_);
  not (_06469_, _06460_);
  nor (_06470_, _05731_, _05659_);
  and (_06471_, _05697_, _05685_);
  nor (_06472_, _05726_, _05671_);
  and (_06473_, _06472_, _06471_);
  and (_06474_, _06473_, _06470_);
  nor (_06475_, _06474_, _06469_);
  not (_06476_, _06475_);
  and (_06477_, _06093_, _05739_);
  not (_06478_, _06477_);
  and (_06479_, _06239_, \oc8051_golden_model_1.SP [2]);
  not (_06480_, _06479_);
  and (_06481_, _06450_, _05746_);
  and (_06482_, _06450_, _05735_);
  nor (_06483_, _06482_, _06481_);
  and (_06484_, _06483_, _06480_);
  and (_06485_, _06484_, _06478_);
  and (_06486_, _06471_, _05689_);
  nor (_06487_, _06486_, _06451_);
  not (_06488_, _06487_);
  and (_06489_, _06450_, _05726_);
  and (_06490_, _06460_, _05735_);
  nor (_06491_, _06490_, _06489_);
  and (_06492_, _06450_, _05671_);
  and (_06493_, _06460_, _05746_);
  nor (_06494_, _06493_, _06492_);
  and (_06495_, _06494_, _06491_);
  and (_06496_, _06495_, _06488_);
  and (_06497_, _06496_, _06485_);
  and (_06498_, _06497_, _06476_);
  and (_06499_, _06498_, _06468_);
  not (_06500_, _06499_);
  nor (_06501_, _06500_, _06446_);
  and (_06502_, _06501_, _06414_);
  and (_06503_, _06502_, _06372_);
  and (_06504_, _06503_, _06370_);
  not (_06505_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_06506_, _06048_, _06016_);
  not (_06507_, _06506_);
  nor (_06508_, _06267_, _06016_);
  not (_06509_, _06121_);
  nor (_06510_, _06509_, _06016_);
  or (_06511_, _06220_, _06016_);
  nor (_06512_, _06242_, _06016_);
  and (_06513_, _06024_, _06113_);
  and (_06514_, _06513_, _06042_);
  not (_06515_, _06514_);
  and (_06516_, _06122_, _06042_);
  not (_06517_, _06096_);
  nor (_06518_, _06136_, _06227_);
  nand (_06519_, _06518_, _06517_);
  and (_06520_, _06519_, _06042_);
  nor (_06521_, _06520_, _06516_);
  and (_06522_, _06521_, _06515_);
  not (_06523_, _05697_);
  and (_06524_, _06227_, _06523_);
  and (_06525_, _06096_, _06523_);
  nor (_06526_, _06525_, _06524_);
  and (_06527_, _06513_, _06523_);
  or (_06528_, _06527_, _06241_);
  not (_06529_, _06528_);
  and (_06530_, _06122_, _06523_);
  nor (_06531_, _06530_, _06102_);
  and (_06532_, _06136_, _06523_);
  not (_06533_, _05703_);
  and (_06534_, _06513_, _06533_);
  nor (_06535_, _06534_, _06532_);
  and (_06536_, _06535_, _06531_);
  and (_06537_, _06536_, _06529_);
  and (_06538_, _06537_, _06526_);
  and (_06539_, _06538_, _06522_);
  or (_06540_, _06539_, _06512_);
  nand (_06541_, _06540_, _06044_);
  nand (_06542_, _06045_, _06541_);
  and (_06543_, _06239_, _06029_);
  nor (_06544_, _06543_, _06219_);
  not (_06545_, _05648_);
  and (_06546_, _06450_, _06037_);
  and (_06547_, _06135_, _06037_);
  nor (_06548_, _06547_, _06546_);
  nor (_06549_, _06548_, _06545_);
  not (_06550_, _06549_);
  and (_06551_, _06136_, _06037_);
  not (_06552_, _06551_);
  and (_06553_, _06513_, _06037_);
  and (_06554_, _06096_, _06037_);
  nor (_06555_, _06554_, _06553_);
  and (_06556_, _06555_, _06552_);
  and (_06557_, _06556_, _06550_);
  and (_06558_, _06557_, _06544_);
  nand (_06559_, _06558_, _06542_);
  nand (_06560_, _06559_, _06511_);
  and (_06561_, _06560_, _06040_);
  or (_06562_, _06041_, _06561_);
  and (_06563_, _06038_, _06016_);
  nor (_06564_, _06122_, _06018_);
  nor (_06565_, _06513_, _06096_);
  and (_06566_, _06565_, _06564_);
  and (_06567_, _06566_, _06518_);
  nor (_06568_, _06567_, _05685_);
  nor (_06569_, _06568_, _06563_);
  and (_06570_, _06569_, _06562_);
  or (_06571_, _06570_, _06510_);
  nand (_06572_, _06571_, _06254_);
  not (_06573_, _06233_);
  nor (_06574_, _06254_, _05984_);
  nor (_06575_, _06574_, _06573_);
  nand (_06576_, _06575_, _06572_);
  and (_06577_, _06573_, _06016_);
  not (_06578_, _06252_);
  and (_06579_, _06513_, _06221_);
  nor (_06580_, _06579_, _06578_);
  not (_06581_, _06580_);
  nor (_06582_, _06581_, _06577_);
  and (_06583_, _06582_, _06576_);
  nor (_06584_, _06252_, _05984_);
  or (_06585_, _06584_, _06583_);
  nor (_06586_, _06096_, _06018_);
  and (_06587_, _06093_, _05648_);
  not (_06588_, _06587_);
  and (_06589_, _06588_, _06586_);
  nor (_06590_, _06589_, _05672_);
  and (_06591_, _06513_, _05671_);
  and (_06592_, _06135_, _05671_);
  and (_06593_, _06592_, _05648_);
  nor (_06594_, _06593_, _06591_);
  not (_06595_, _06594_);
  nor (_06596_, _06595_, _06590_);
  and (_06597_, _06596_, _06585_);
  or (_06598_, _06597_, _06508_);
  and (_06599_, _06598_, _06027_);
  nor (_06600_, _06599_, _06028_);
  nor (_06601_, _06567_, _05660_);
  nor (_06602_, _06601_, _06600_);
  and (_06603_, _06161_, _04306_);
  and (_06604_, _06194_, _04335_);
  nor (_06605_, _06604_, _06603_);
  and (_06606_, _06170_, _04322_);
  and (_06607_, _06175_, _04333_);
  nor (_06608_, _06607_, _06606_);
  and (_06609_, _06608_, _06605_);
  and (_06610_, _06179_, _04337_);
  and (_06611_, _06182_, _04324_);
  nor (_06612_, _06611_, _06610_);
  and (_06613_, _06185_, _04327_);
  and (_06614_, _06187_, _04317_);
  nor (_06615_, _06614_, _06613_);
  and (_06616_, _06615_, _06612_);
  and (_06617_, _06616_, _06609_);
  and (_06618_, _06192_, _04319_);
  and (_06619_, _06166_, _04347_);
  nor (_06620_, _06619_, _06618_);
  and (_06621_, _06197_, _04329_);
  and (_06622_, _06199_, _04308_);
  nor (_06623_, _06622_, _06621_);
  and (_06624_, _06623_, _06620_);
  and (_06625_, _06203_, _04344_);
  and (_06626_, _06205_, _04339_);
  nor (_06627_, _06626_, _06625_);
  and (_06628_, _06208_, _04313_);
  and (_06629_, _06210_, _04311_);
  nor (_06630_, _06629_, _06628_);
  and (_06631_, _06630_, _06627_);
  and (_06632_, _06631_, _06624_);
  and (_06633_, _06632_, _06617_);
  nor (_06634_, _06633_, _05669_);
  or (_06635_, _06634_, _06602_);
  not (_06636_, _06088_);
  and (_06637_, _06089_, _05984_);
  and (_06638_, _06513_, _05723_);
  nor (_06639_, _06638_, _06637_);
  and (_06640_, _06639_, _06636_);
  and (_06641_, _06640_, _06635_);
  nor (_06642_, _06636_, _05984_);
  or (_06643_, _06642_, _06641_);
  not (_06644_, _05726_);
  nor (_06645_, _06518_, _06644_);
  not (_06646_, _06645_);
  and (_06647_, _06513_, _05726_);
  not (_06648_, _06647_);
  and (_06649_, _06122_, _05726_);
  and (_06650_, _06096_, _05726_);
  nor (_06651_, _06650_, _06649_);
  and (_06652_, _06651_, _06648_);
  and (_06653_, _06652_, _06646_);
  and (_06654_, _06653_, _06643_);
  nor (_06655_, _06286_, _06017_);
  not (_06656_, _05735_);
  not (_06657_, _06227_);
  and (_06658_, _06565_, _06657_);
  and (_06659_, _06588_, _06658_);
  nor (_06660_, _06659_, _06656_);
  nor (_06661_, _06660_, _06655_);
  and (_06663_, _06661_, _06654_);
  nor (_06664_, _06281_, _06017_);
  and (_06665_, _06227_, _05739_);
  not (_06666_, _06665_);
  and (_06667_, _06096_, _05739_);
  not (_06668_, _06667_);
  and (_06669_, _06513_, _05739_);
  and (_06670_, _06587_, _05739_);
  nor (_06671_, _06670_, _06669_);
  and (_06672_, _06671_, _06668_);
  and (_06673_, _06672_, _06666_);
  not (_06674_, _06673_);
  nor (_06675_, _06674_, _06664_);
  and (_06676_, _06675_, _06663_);
  nor (_06677_, _06294_, _06017_);
  not (_06678_, _05731_);
  nor (_06679_, _06567_, _06678_);
  nor (_06680_, _06679_, _06677_);
  and (_06681_, _06680_, _06676_);
  nor (_06682_, _06289_, _06016_);
  or (_06683_, _06682_, _06681_);
  and (_06684_, _06298_, _06029_);
  nor (_06685_, _06684_, _06129_);
  and (_06686_, _06685_, _06683_);
  nor (_06687_, _06306_, _05984_);
  or (_06688_, _06687_, _06686_);
  nor (_06689_, _06493_, _06481_);
  or (_06690_, _06689_, _06545_);
  and (_06691_, _06227_, _05746_);
  and (_06692_, _06513_, _05746_);
  and (_06693_, _06096_, _05746_);
  or (_06694_, _06693_, _06051_);
  or (_06695_, _06694_, _06692_);
  nor (_06696_, _06695_, _06691_);
  and (_06697_, _06696_, _06690_);
  and (_06698_, _06697_, _06688_);
  nor (_06699_, _06052_, _06016_);
  or (_06700_, _06699_, _06698_);
  and (_06701_, _06049_, _06029_);
  nor (_06702_, _06701_, _06126_);
  and (_06703_, _06702_, _06700_);
  not (_06704_, _06126_);
  nor (_06705_, _06704_, _05984_);
  or (_06706_, _06705_, _06703_);
  and (_06707_, _06227_, _05495_);
  and (_06708_, _06096_, _05495_);
  or (_06709_, _06708_, _06707_);
  not (_06710_, _06709_);
  and (_06711_, _06122_, _05495_);
  and (_06712_, _06513_, _05495_);
  nor (_06713_, _06712_, _06711_);
  nor (_06714_, _06457_, _06316_);
  and (_06715_, _06714_, _06713_);
  and (_06716_, _06715_, _06710_);
  and (_06717_, _06716_, _06706_);
  not (_06718_, _06316_);
  nor (_06719_, _06718_, _06016_);
  or (_06720_, _06719_, _06717_);
  and (_06721_, _06720_, _05653_);
  nor (_06722_, _06721_, _05985_);
  not (_06723_, _05750_);
  nor (_06724_, _06567_, _06723_);
  or (_06725_, _06724_, _06722_);
  nand (_06726_, _06725_, _06507_);
  or (_06727_, _06726_, _06505_);
  nor (_06728_, _05934_, _00260_);
  nor (_06729_, _05887_, _00219_);
  nor (_06730_, _06729_, _06728_);
  nor (_06731_, _05894_, _00168_);
  nor (_06732_, _05945_, _00065_);
  nor (_06733_, _06732_, _06731_);
  and (_06734_, _06733_, _06730_);
  nor (_06735_, _05902_, _00607_);
  nor (_06736_, _05940_, _00550_);
  nor (_06737_, _06736_, _06735_);
  nor (_06738_, _05919_, _00506_);
  nor (_06739_, _05913_, _00383_);
  nor (_06740_, _06739_, _06738_);
  and (_06741_, _06740_, _06737_);
  and (_06742_, _06741_, _06734_);
  nor (_06743_, _05915_, _00342_);
  nor (_06744_, _05929_, _43752_);
  nor (_06745_, _06744_, _06743_);
  nor (_06746_, _05907_, _00424_);
  nor (_06747_, _05947_, _43793_);
  nor (_06748_, _06747_, _06746_);
  and (_06749_, _06748_, _06745_);
  nor (_06750_, _05942_, _00301_);
  nor (_06751_, _05931_, _00024_);
  nor (_06752_, _06751_, _06750_);
  nor (_06753_, _05923_, _00465_);
  nor (_06754_, _05936_, _00106_);
  nor (_06755_, _06754_, _06753_);
  and (_06756_, _06755_, _06752_);
  and (_06757_, _06756_, _06749_);
  and (_06758_, _06757_, _06742_);
  nor (_06759_, _06758_, _05952_);
  nor (_06760_, _06039_, _05652_);
  and (_06761_, _06760_, _06090_);
  and (_06762_, _06761_, _06364_);
  and (_06763_, _06762_, _06362_);
  not (_06764_, _06763_);
  and (_06765_, _06764_, _06759_);
  not (_06766_, _06765_);
  and (_06767_, _06759_, _06026_);
  not (_06768_, _06767_);
  nor (_06769_, _05907_, _00409_);
  nor (_06770_, _05934_, _00245_);
  nor (_06771_, _06770_, _06769_);
  nor (_06772_, _05887_, _00204_);
  nor (_06773_, _05947_, _43778_);
  nor (_06774_, _06773_, _06772_);
  and (_06775_, _06774_, _06771_);
  nor (_06776_, _05902_, _00592_);
  nor (_06777_, _05945_, _00050_);
  nor (_06778_, _06777_, _06776_);
  nor (_06779_, _05940_, _00532_);
  nor (_06780_, _05942_, _00286_);
  nor (_06781_, _06780_, _06779_);
  and (_06782_, _06781_, _06778_);
  and (_06783_, _06782_, _06775_);
  nor (_06784_, _05894_, _00135_);
  nor (_06785_, _05936_, _00091_);
  nor (_06786_, _06785_, _06784_);
  nor (_06787_, _05913_, _00368_);
  nor (_06788_, _05929_, _43737_);
  nor (_06789_, _06788_, _06787_);
  and (_06790_, _06789_, _06786_);
  nor (_06791_, _05919_, _00491_);
  nor (_06792_, _05931_, _00009_);
  nor (_06793_, _06792_, _06791_);
  nor (_06794_, _05923_, _00450_);
  nor (_06795_, _05915_, _00327_);
  nor (_06796_, _06795_, _06794_);
  and (_06797_, _06796_, _06793_);
  and (_06798_, _06797_, _06790_);
  and (_06799_, _06798_, _06783_);
  nor (_06800_, _06799_, _06412_);
  not (_06801_, _06800_);
  and (_06802_, _06194_, _04382_);
  and (_06803_, _06205_, _04386_);
  nor (_06804_, _06803_, _06802_);
  and (_06805_, _06185_, _04374_);
  and (_06806_, _06175_, _04380_);
  nor (_06807_, _06806_, _06805_);
  and (_06808_, _06807_, _06804_);
  and (_06809_, _06161_, _04353_);
  and (_06810_, _06203_, _04391_);
  nor (_06811_, _06810_, _06809_);
  and (_06812_, _06192_, _04366_);
  and (_06813_, _06166_, _04393_);
  nor (_06814_, _06813_, _06812_);
  and (_06815_, _06814_, _06811_);
  and (_06816_, _06815_, _06808_);
  and (_06817_, _06210_, _04358_);
  and (_06818_, _06182_, _04371_);
  nor (_06819_, _06818_, _06817_);
  and (_06820_, _06170_, _04369_);
  and (_06821_, _06208_, _04360_);
  nor (_06822_, _06821_, _06820_);
  and (_06823_, _06822_, _06819_);
  and (_06824_, _06179_, _04384_);
  and (_06825_, _06187_, _04364_);
  nor (_06826_, _06825_, _06824_);
  and (_06827_, _06197_, _04376_);
  and (_06828_, _06199_, _04355_);
  nor (_06829_, _06828_, _06827_);
  and (_06830_, _06829_, _06826_);
  and (_06831_, _06830_, _06823_);
  and (_06832_, _06831_, _06816_);
  nor (_06833_, _06832_, _05669_);
  and (_06834_, _06135_, _05739_);
  and (_06835_, _06135_, _05735_);
  nor (_06836_, _06835_, _06834_);
  and (_06837_, _06135_, _06031_);
  nor (_06838_, _06592_, _06837_);
  and (_06839_, _06838_, _06836_);
  and (_06840_, _06839_, _06488_);
  not (_06841_, _05746_);
  nor (_06842_, _05739_, _05735_);
  and (_06843_, _06842_, _06841_);
  nor (_06844_, _06843_, _06451_);
  nor (_06845_, _06844_, _06455_);
  and (_06846_, _06845_, _06840_);
  not (_06847_, \oc8051_golden_model_1.SP [1]);
  not (_06848_, _06239_);
  and (_06849_, _06448_, _06848_);
  nor (_06850_, _06849_, _06847_);
  not (_06851_, _06850_);
  not (_06852_, _06229_);
  nor (_06853_, _05746_, _06523_);
  nor (_06854_, _06853_, _06852_);
  not (_06855_, _06854_);
  nor (_06856_, _06450_, _06135_);
  nor (_06857_, _05750_, _05726_);
  nor (_06858_, _06857_, _06856_);
  not (_06859_, _06135_);
  nor (_06860_, _06470_, _06859_);
  nor (_06861_, _06860_, _06858_);
  and (_06862_, _06861_, _06855_);
  and (_06863_, _06135_, _06042_);
  not (_06864_, _06863_);
  and (_06865_, _06229_, _05495_);
  nor (_06866_, _06865_, _06707_);
  and (_06867_, _06866_, _06864_);
  nor (_06868_, _06547_, _06492_);
  and (_06869_, _06868_, _06867_);
  nor (_06870_, _06691_, _06524_);
  and (_06871_, _06870_, _06869_);
  and (_06872_, _06871_, _06862_);
  and (_06873_, _06872_, _06851_);
  and (_06874_, _06873_, _06846_);
  not (_06875_, _06874_);
  nor (_06876_, _06875_, _06833_);
  and (_06877_, _06876_, _06801_);
  and (_06878_, _06877_, _06768_);
  and (_06879_, _06878_, _06766_);
  not (_06880_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_06881_, _06725_, _06507_);
  or (_06882_, _06881_, _06880_);
  and (_06883_, _06882_, _06879_);
  nand (_06884_, _06883_, _06727_);
  not (_06885_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_06886_, _06881_, _06885_);
  not (_06887_, _06879_);
  not (_06888_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_06889_, _06726_, _06888_);
  and (_06890_, _06889_, _06887_);
  nand (_06891_, _06890_, _06886_);
  nand (_06892_, _06891_, _06884_);
  nand (_06893_, _06892_, _06504_);
  not (_06894_, _06504_);
  not (_06895_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_06896_, _06881_, _06895_);
  nand (_06897_, _06881_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_06898_, _06897_, _06887_);
  nand (_06899_, _06898_, _06896_);
  nand (_06900_, _06881_, \oc8051_golden_model_1.IRAM[4] [0]);
  nand (_06901_, _06726_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_06902_, _06901_, _06879_);
  nand (_06903_, _06902_, _06900_);
  nand (_06904_, _06903_, _06899_);
  nand (_06905_, _06904_, _06894_);
  nand (_06906_, _06905_, _06893_);
  nand (_06907_, _06906_, _06328_);
  not (_06908_, _06328_);
  nand (_06909_, _06726_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_06910_, _06881_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_06911_, _06910_, _06887_);
  nand (_06912_, _06911_, _06909_);
  nand (_06913_, _06881_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand (_06914_, _06726_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_06915_, _06914_, _06879_);
  nand (_06916_, _06915_, _06913_);
  nand (_06917_, _06916_, _06912_);
  nand (_06918_, _06917_, _06504_);
  nand (_06919_, _06726_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_06920_, _06881_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_06921_, _06920_, _06887_);
  nand (_06922_, _06921_, _06919_);
  nand (_06923_, _06881_, \oc8051_golden_model_1.IRAM[12] [0]);
  nand (_06924_, _06726_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_06925_, _06924_, _06879_);
  nand (_06926_, _06925_, _06923_);
  nand (_06927_, _06926_, _06922_);
  nand (_06928_, _06927_, _06894_);
  nand (_06929_, _06928_, _06918_);
  nand (_06930_, _06929_, _06908_);
  and (_06931_, _06930_, _06907_);
  and (_06932_, _06931_, _06046_);
  nor (_06933_, _06114_, _05718_);
  and (_06934_, _06933_, _06565_);
  nor (_06935_, _06934_, _05703_);
  not (_06936_, _06935_);
  nor (_06937_, _06936_, _06932_);
  and (_06938_, _06094_, _06523_);
  not (_06939_, _06938_);
  nor (_06940_, _06939_, _05952_);
  and (_06941_, _06940_, _06016_);
  nor (_06942_, _06941_, _06937_);
  and (_06943_, _06098_, _06523_);
  and (_06944_, _06943_, \oc8051_golden_model_1.SP [0]);
  not (_06945_, _06944_);
  and (_06946_, _06945_, _06521_);
  and (_06947_, _06946_, _06942_);
  and (_06948_, _06103_, _06042_);
  not (_06949_, _06948_);
  nor (_06950_, _06949_, _06931_);
  not (_06951_, _06950_);
  and (_06952_, _06951_, _06947_);
  nor (_06953_, _06044_, _05952_);
  not (_06954_, _06102_);
  nor (_06955_, _06954_, _05952_);
  and (_06956_, _06955_, _06016_);
  nor (_06957_, _06956_, _06953_);
  and (_06958_, _06957_, _06952_);
  not (_06959_, _06958_);
  and (_06960_, _06959_, _06045_);
  nor (_06961_, _05690_, _06029_);
  nor (_06962_, _06961_, _06960_);
  nor (_06963_, _06848_, _05952_);
  and (_06964_, _06963_, _06016_);
  or (_06965_, _06554_, _06551_);
  nor (_06966_, _06965_, _06549_);
  not (_06967_, _06966_);
  nor (_06968_, _06967_, _06964_);
  and (_06969_, _06968_, _06962_);
  and (_06970_, _06103_, _06037_);
  not (_06971_, _06970_);
  nor (_06972_, _06971_, _06931_);
  not (_06973_, _06972_);
  and (_06974_, _06973_, _06969_);
  nor (_06975_, _06040_, _05952_);
  nor (_06976_, _06220_, _05952_);
  and (_06977_, _06976_, _06016_);
  nor (_06978_, _06977_, _06975_);
  and (_06979_, _06978_, _06974_);
  nor (_06980_, _06979_, _06041_);
  or (_06981_, _06980_, _06038_);
  nand (_06982_, _06038_, _06029_);
  nand (_06983_, _06982_, _06981_);
  and (_06984_, _06983_, _06036_);
  nor (_06985_, _06984_, _06034_);
  or (_06986_, _06228_, _06224_);
  and (_06987_, _06587_, _06221_);
  or (_06988_, _06987_, _06986_);
  or (_06989_, _06988_, _06985_);
  nor (_06990_, _06989_, _06030_);
  nor (_06991_, _06027_, _05952_);
  and (_06992_, _06103_, _06221_);
  not (_06993_, _06992_);
  nor (_06994_, _06993_, _06931_);
  nor (_06995_, _06994_, _06991_);
  and (_06996_, _06995_, _06990_);
  nor (_06997_, _06996_, _06028_);
  nor (_06998_, _06997_, _06023_);
  nor (_06999_, _05673_, \oc8051_golden_model_1.SP [0]);
  nor (_07000_, _06999_, _06998_);
  nor (_07001_, _05952_, _05660_);
  and (_07002_, _06095_, _05610_);
  or (_07003_, _07002_, _06136_);
  and (_07004_, _07003_, _07001_);
  or (_07005_, _06450_, _06098_);
  nor (_07006_, _07005_, _06135_);
  not (_07007_, _07006_);
  and (_07008_, _07007_, _07001_);
  nor (_07009_, _07008_, _07004_);
  nor (_07010_, _05952_, _05669_);
  and (_07011_, _06103_, _05659_);
  not (_07012_, _07011_);
  nor (_07013_, _07012_, _05952_);
  nor (_07014_, _07013_, _07010_);
  and (_07015_, _07014_, _07009_);
  nor (_07016_, _07015_, _06017_);
  and (_07017_, _05648_, _05567_);
  and (_07018_, _07017_, _05723_);
  nor (_07019_, _07018_, _07016_);
  not (_07020_, _07019_);
  nor (_07021_, _07020_, _07000_);
  not (_07022_, _06931_);
  and (_07023_, _06103_, _05723_);
  and (_07024_, _07023_, _07022_);
  nor (_07025_, _07024_, _06021_);
  and (_07026_, _07025_, _07021_);
  nor (_07027_, _07026_, _06022_);
  nor (_07028_, _07027_, _05724_);
  and (_07029_, _05724_, _06029_);
  nor (_07030_, _07029_, _07028_);
  nor (_07031_, _06278_, _05952_);
  not (_07032_, _06108_);
  and (_07033_, _06285_, _07032_);
  nor (_07034_, _07033_, _05952_);
  nor (_07035_, _07034_, _07031_);
  nor (_07036_, _07035_, _06017_);
  nor (_07037_, _07036_, _05736_);
  not (_07038_, _07037_);
  nor (_07039_, _07038_, _07030_);
  and (_07040_, _05736_, _06029_);
  nor (_07041_, _07040_, _07039_);
  nor (_07042_, _06293_, _05952_);
  and (_07043_, _07042_, _06016_);
  nor (_07044_, _07043_, _07041_);
  and (_07045_, _05732_, \oc8051_golden_model_1.SP [0]);
  and (_07046_, _06587_, _05495_);
  nor (_07047_, _07046_, _07045_);
  and (_07048_, _07047_, _06710_);
  and (_07049_, _07048_, _07044_);
  nor (_07050_, _06718_, _05952_);
  and (_07051_, _06103_, _05495_);
  not (_07052_, _07051_);
  nor (_07053_, _07052_, _06931_);
  nor (_07054_, _07053_, _07050_);
  and (_07055_, _07054_, _07049_);
  and (_07056_, _07050_, _06017_);
  nor (_07057_, _07056_, _07055_);
  nor (_07058_, _05952_, _05653_);
  nor (_07059_, _06127_, _05752_);
  nor (_07060_, _07059_, _06029_);
  nor (_07061_, _07060_, _07058_);
  not (_07062_, _07061_);
  nor (_07063_, _07062_, _07057_);
  nor (_07064_, _07063_, _05985_);
  and (_07065_, _07017_, _05750_);
  nor (_07066_, _07065_, _07064_);
  nor (_07067_, _06048_, _05952_);
  and (_07068_, _06103_, _05750_);
  not (_07069_, _07068_);
  nor (_07070_, _07069_, _06931_);
  nor (_07071_, _07070_, _07067_);
  and (_07072_, _07071_, _07066_);
  and (_07073_, _07067_, _06017_);
  nor (_07074_, _07073_, _07072_);
  not (_07075_, _07074_);
  not (_07076_, _06799_);
  and (_07077_, _07067_, _07076_);
  and (_07078_, _06460_, _05750_);
  and (_07079_, _06759_, _05652_);
  and (_07080_, _06847_, \oc8051_golden_model_1.SP [0]);
  and (_07081_, \oc8051_golden_model_1.SP [1], _06029_);
  nor (_07082_, _07081_, _07080_);
  not (_07083_, _07082_);
  nor (_07084_, _07083_, _07059_);
  and (_07085_, _07083_, _05732_);
  and (_07086_, _07076_, _06021_);
  and (_07087_, _06103_, _06533_);
  nand (_07088_, _06881_, \oc8051_golden_model_1.IRAM[0] [1]);
  nand (_07089_, _06726_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_07090_, _07089_, _06879_);
  nand (_07091_, _07090_, _07088_);
  nand (_07092_, _06726_, \oc8051_golden_model_1.IRAM[3] [1]);
  nand (_07093_, _06881_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_07094_, _07093_, _06887_);
  nand (_07095_, _07094_, _07092_);
  nand (_07096_, _07095_, _07091_);
  nand (_07097_, _07096_, _06504_);
  nand (_07098_, _06726_, \oc8051_golden_model_1.IRAM[7] [1]);
  nand (_07099_, _06881_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_07100_, _07099_, _06887_);
  nand (_07101_, _07100_, _07098_);
  nand (_07102_, _06881_, \oc8051_golden_model_1.IRAM[4] [1]);
  nand (_07103_, _06726_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_07104_, _07103_, _06879_);
  nand (_07105_, _07104_, _07102_);
  nand (_07106_, _07105_, _07101_);
  nand (_07107_, _07106_, _06894_);
  nand (_07108_, _07107_, _07097_);
  nand (_07109_, _07108_, _06328_);
  nand (_07110_, _06726_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_07111_, _06881_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_07112_, _07111_, _06887_);
  nand (_07113_, _07112_, _07110_);
  nand (_07114_, _06881_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_07115_, _06726_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_07116_, _07115_, _06879_);
  nand (_07117_, _07116_, _07114_);
  nand (_07118_, _07117_, _07113_);
  nand (_07119_, _07118_, _06504_);
  nand (_07120_, _06726_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_07121_, _06881_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_07122_, _07121_, _06887_);
  nand (_07123_, _07122_, _07120_);
  nand (_07124_, _06881_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand (_07125_, _06726_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_07126_, _07125_, _06879_);
  nand (_07127_, _07126_, _07124_);
  nand (_07128_, _07127_, _07123_);
  nand (_07129_, _07128_, _06894_);
  nand (_07130_, _07129_, _07119_);
  nand (_07131_, _07130_, _06908_);
  nand (_07132_, _07131_, _07109_);
  and (_07133_, _07132_, _06046_);
  or (_07134_, _07133_, _07087_);
  and (_07135_, _06940_, _06799_);
  or (_07136_, _07135_, _07134_);
  and (_07137_, _07082_, _06943_);
  not (_07138_, _07137_);
  and (_07139_, _07002_, _06042_);
  nor (_07140_, _07139_, _06461_);
  and (_07141_, _07140_, _07138_);
  not (_07142_, _07141_);
  nor (_07143_, _07142_, _07136_);
  and (_07144_, _07132_, _06948_);
  nor (_07145_, _07144_, _06955_);
  and (_07146_, _07145_, _07143_);
  and (_07147_, _06955_, _07076_);
  nor (_07148_, _07147_, _07146_);
  and (_07149_, _06758_, _06953_);
  nor (_07150_, _07149_, _07148_);
  or (_07151_, _07083_, _05690_);
  nand (_07152_, _07151_, _07150_);
  and (_07153_, _06963_, _06799_);
  and (_07154_, _07002_, _06037_);
  nor (_07155_, _07154_, _06463_);
  not (_07156_, _07155_);
  nor (_07157_, _07156_, _07153_);
  not (_07158_, _07157_);
  nor (_07159_, _07158_, _07152_);
  and (_07160_, _07132_, _06970_);
  nor (_07161_, _07160_, _06976_);
  and (_07162_, _07161_, _07159_);
  and (_07163_, _06976_, _07076_);
  nor (_07164_, _07163_, _07162_);
  and (_07165_, _06758_, _06975_);
  nor (_07166_, _07165_, _06038_);
  not (_07167_, _07166_);
  nor (_07168_, _07167_, _07164_);
  and (_07169_, _07083_, _06038_);
  nor (_07170_, _07169_, _07168_);
  and (_07171_, _06035_, _06758_);
  nor (_07172_, _07171_, _07170_);
  nand (_07173_, _06222_, _05610_);
  and (_07174_, _07002_, _06221_);
  nor (_07175_, _07083_, _05686_);
  nor (_07176_, _07175_, _07174_);
  and (_07177_, _07176_, _07173_);
  and (_07178_, _07177_, _07172_);
  and (_07179_, _07132_, _06992_);
  nor (_07180_, _07179_, _06991_);
  and (_07181_, _07180_, _07178_);
  nor (_07182_, _07181_, _06767_);
  nor (_07183_, _07182_, _06023_);
  nor (_07184_, _07082_, _05673_);
  nor (_07185_, _07184_, _07183_);
  nor (_07186_, _07015_, _07076_);
  and (_07187_, _05723_, _05610_);
  and (_07188_, _07187_, _05567_);
  nor (_07189_, _07188_, _07186_);
  not (_07190_, _07189_);
  nor (_07191_, _07190_, _07185_);
  and (_07192_, _07132_, _07023_);
  nor (_07193_, _07192_, _06021_);
  and (_07194_, _07193_, _07191_);
  nor (_07195_, _07194_, _07086_);
  nor (_07196_, _07195_, _05724_);
  and (_07197_, _07083_, _05724_);
  nor (_07198_, _07197_, _07196_);
  nor (_07199_, _07035_, _07076_);
  nor (_07200_, _07199_, _05736_);
  not (_07201_, _07200_);
  nor (_07202_, _07201_, _07198_);
  and (_07203_, _07083_, _05736_);
  nor (_07204_, _07203_, _07202_);
  and (_07205_, _07042_, _06799_);
  nor (_07206_, _07205_, _05732_);
  not (_07207_, _07206_);
  nor (_07208_, _07207_, _07204_);
  nor (_07209_, _07208_, _07085_);
  and (_07210_, _07002_, _05495_);
  not (_07211_, _07210_);
  and (_07212_, _07211_, _06459_);
  not (_07213_, _07212_);
  nor (_07214_, _07213_, _07209_);
  and (_07215_, _07132_, _07051_);
  nor (_07216_, _07215_, _07050_);
  and (_07217_, _07216_, _07214_);
  and (_07218_, _07050_, _07076_);
  nor (_07219_, _07218_, _07217_);
  or (_07220_, _07219_, _07058_);
  nor (_07221_, _07220_, _07084_);
  nor (_07222_, _07221_, _07079_);
  and (_07223_, _07002_, _05750_);
  or (_07224_, _07223_, _07222_);
  nor (_07225_, _07224_, _07078_);
  and (_07226_, _07132_, _07068_);
  nor (_07227_, _07226_, _07067_);
  and (_07228_, _07227_, _07225_);
  nor (_07229_, _07228_, _07077_);
  not (_07230_, _00000_);
  not (_07231_, _07013_);
  not (_07232_, _07067_);
  not (_07233_, _06943_);
  and (_07234_, _07059_, _07233_);
  nor (_07235_, _05736_, _05732_);
  and (_07236_, _06867_, _07235_);
  and (_07237_, _07236_, _07234_);
  and (_07238_, _06450_, _06042_);
  nor (_07239_, _06948_, _07238_);
  and (_07240_, _07239_, _06548_);
  nor (_07241_, _06554_, _06038_);
  nor (_07242_, _07051_, _06992_);
  and (_07243_, _07242_, _07241_);
  and (_07244_, _07243_, _07240_);
  and (_07245_, _07244_, _07237_);
  nand (_07246_, _06933_, _05668_);
  and (_07247_, _07246_, _06533_);
  nor (_07248_, _07002_, _06103_);
  nor (_07249_, _07248_, _05703_);
  or (_07250_, _07249_, _07247_);
  not (_07251_, _07250_);
  and (_07252_, _06095_, _05723_);
  not (_07253_, _07252_);
  and (_07254_, _06094_, _05723_);
  and (_07255_, _06222_, _06545_);
  nor (_07256_, _07255_, _07254_);
  and (_07257_, _07256_, _07253_);
  and (_07258_, _07257_, _07251_);
  and (_07259_, _07258_, _07245_);
  and (_07260_, _07069_, _06467_);
  and (_07261_, _06133_, _06037_);
  nor (_07262_, _07261_, _07139_);
  nor (_07263_, _07210_, _07174_);
  and (_07264_, _07263_, _07262_);
  nor (_07265_, _06987_, _06970_);
  and (_07266_, _06093_, _05661_);
  and (_07267_, _07266_, _05723_);
  nor (_07268_, _07267_, _07023_);
  and (_07269_, _07268_, _07265_);
  and (_07270_, _07269_, _07264_);
  and (_07271_, _05686_, _05673_);
  not (_07272_, _05690_);
  nor (_07273_, _05724_, _07272_);
  and (_07274_, _07273_, _07271_);
  and (_07275_, _06135_, _06221_);
  and (_07276_, _06135_, _05750_);
  nor (_07277_, _07276_, _07275_);
  and (_07278_, _06450_, _05495_);
  nor (_07279_, _07223_, _07278_);
  and (_07280_, _07279_, _07277_);
  and (_07281_, _07280_, _07274_);
  and (_07282_, _07281_, _07270_);
  and (_07283_, _07282_, _07260_);
  and (_07284_, _07283_, _07259_);
  and (_07285_, _07284_, _07232_);
  and (_07286_, _07285_, _07231_);
  and (_07287_, _07286_, _07009_);
  nor (_07288_, _06976_, _06963_);
  nor (_07289_, _06955_, _06940_);
  and (_07290_, _07289_, _07288_);
  nor (_07291_, _07042_, _06021_);
  nor (_07292_, _07010_, _06975_);
  and (_07293_, _07292_, _07291_);
  and (_07294_, _07293_, _07290_);
  not (_07295_, _07058_);
  nor (_07296_, _07050_, _07034_);
  and (_07297_, _07296_, _07295_);
  nor (_07298_, _06035_, _06953_);
  nor (_07299_, _07031_, _06991_);
  and (_07300_, _07299_, _07298_);
  and (_07301_, _07300_, _07297_);
  and (_07302_, _07301_, _07294_);
  and (_07303_, _07302_, _07287_);
  nor (_07304_, _07303_, _07230_);
  not (_07305_, _07304_);
  nor (_07306_, _07305_, _07229_);
  and (_07307_, _07306_, _07075_);
  not (_07308_, _06991_);
  nand (_07309_, _06881_, \oc8051_golden_model_1.IRAM[0] [3]);
  nand (_07310_, _06726_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_07311_, _07310_, _06879_);
  nand (_07312_, _07311_, _07309_);
  nand (_07313_, _06726_, \oc8051_golden_model_1.IRAM[3] [3]);
  nand (_07314_, _06881_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_07315_, _07314_, _06887_);
  nand (_07316_, _07315_, _07313_);
  nand (_07317_, _07316_, _07312_);
  nand (_07318_, _07317_, _06504_);
  nand (_07319_, _06726_, \oc8051_golden_model_1.IRAM[7] [3]);
  nand (_07320_, _06881_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_07321_, _07320_, _06887_);
  nand (_07322_, _07321_, _07319_);
  nand (_07323_, _06881_, \oc8051_golden_model_1.IRAM[4] [3]);
  nand (_07324_, _06726_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_07325_, _07324_, _06879_);
  nand (_07326_, _07325_, _07323_);
  nand (_07327_, _07326_, _07322_);
  nand (_07328_, _07327_, _06894_);
  nand (_07329_, _07328_, _07318_);
  nand (_07330_, _07329_, _06328_);
  nand (_07331_, _06726_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_07332_, _06881_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_07333_, _07332_, _06887_);
  nand (_07334_, _07333_, _07331_);
  nand (_07335_, _06881_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_07336_, _06726_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_07337_, _07336_, _06879_);
  nand (_07338_, _07337_, _07335_);
  nand (_07339_, _07338_, _07334_);
  nand (_07340_, _07339_, _06504_);
  nand (_07341_, _06726_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_07342_, _06881_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_07343_, _07342_, _06887_);
  nand (_07344_, _07343_, _07341_);
  nand (_07345_, _06881_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_07346_, _06726_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_07347_, _07346_, _06879_);
  nand (_07348_, _07347_, _07345_);
  nand (_07349_, _07348_, _07344_);
  nand (_07350_, _07349_, _06894_);
  nand (_07351_, _07350_, _07340_);
  nand (_07352_, _07351_, _06908_);
  nand (_07353_, _07352_, _07330_);
  and (_07354_, _07353_, _06992_);
  not (_07355_, _05686_);
  and (_07356_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_07357_, _07356_, \oc8051_golden_model_1.SP [2]);
  nor (_07358_, _07357_, \oc8051_golden_model_1.SP [3]);
  and (_07359_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_07360_, _07359_, \oc8051_golden_model_1.SP [3]);
  and (_07361_, _07360_, \oc8051_golden_model_1.SP [0]);
  nor (_07362_, _07361_, _07358_);
  and (_07363_, _07362_, _07355_);
  not (_07364_, _06038_);
  and (_07365_, _06953_, _06084_);
  and (_07366_, _07353_, _06948_);
  and (_07367_, _07362_, _06943_);
  and (_07368_, _07353_, _06046_);
  not (_07369_, \oc8051_golden_model_1.PSW [3]);
  and (_07370_, _05705_, _07369_);
  nor (_07371_, _07370_, _06940_);
  not (_07372_, _07371_);
  nor (_07373_, _07372_, _07368_);
  and (_07374_, _06940_, _06299_);
  nor (_07375_, _07374_, _07373_);
  nor (_07376_, _07375_, _06943_);
  or (_07377_, _07376_, _06948_);
  nor (_07378_, _07377_, _07367_);
  or (_07379_, _07378_, _06955_);
  nor (_07380_, _07379_, _07366_);
  and (_07381_, _06955_, _06299_);
  or (_07382_, _07381_, _06953_);
  nor (_07383_, _07382_, _07380_);
  nor (_07384_, _07383_, _07365_);
  nor (_07385_, _07384_, _07272_);
  nor (_07386_, _07362_, _05690_);
  nor (_07387_, _07386_, _06963_);
  not (_07388_, _07387_);
  nor (_07389_, _07388_, _07385_);
  and (_07390_, _06963_, _06299_);
  nor (_07391_, _07390_, _06970_);
  not (_07392_, _07391_);
  nor (_07393_, _07392_, _07389_);
  and (_07394_, _07353_, _06970_);
  nor (_07395_, _07394_, _06976_);
  not (_07396_, _07395_);
  nor (_07397_, _07396_, _07393_);
  and (_07398_, _06976_, _06299_);
  or (_07399_, _07398_, _06975_);
  nor (_07400_, _07399_, _07397_);
  and (_07401_, _06084_, _06975_);
  nor (_07402_, _07401_, _07400_);
  and (_07403_, _07402_, _07364_);
  and (_07404_, _07362_, _06038_);
  or (_07405_, _07404_, _06035_);
  nor (_07406_, _07405_, _07403_);
  and (_07407_, _06032_, _06085_);
  or (_07408_, _07407_, _07355_);
  nor (_07409_, _07408_, _07406_);
  or (_07410_, _07409_, _06992_);
  nor (_07411_, _07410_, _07363_);
  nor (_07412_, _07411_, _07354_);
  and (_07413_, _07412_, _07308_);
  not (_07414_, _06084_);
  and (_07415_, _06991_, _07414_);
  or (_07416_, _07415_, _07413_);
  and (_07417_, _07416_, _05673_);
  and (_07418_, _07362_, _06023_);
  not (_07419_, _07418_);
  and (_07420_, _07419_, _07015_);
  not (_07421_, _07420_);
  nor (_07422_, _07421_, _07417_);
  nor (_07423_, _07015_, _06299_);
  nor (_07424_, _07423_, _07422_);
  nor (_07425_, _07424_, _07023_);
  and (_07426_, _07353_, _07023_);
  nor (_07427_, _07426_, _06021_);
  not (_07428_, _07427_);
  nor (_07429_, _07428_, _07425_);
  nor (_07430_, _06020_, _05984_);
  nor (_07431_, _07430_, _07429_);
  nor (_07432_, _07431_, _05724_);
  and (_07433_, _07362_, _05724_);
  not (_07434_, _07433_);
  and (_07435_, _07434_, _07035_);
  not (_07436_, _07435_);
  nor (_07437_, _07436_, _07432_);
  nor (_07438_, _07035_, _06299_);
  nor (_07439_, _07438_, _05736_);
  not (_07440_, _07439_);
  nor (_07441_, _07440_, _07437_);
  and (_07442_, _07362_, _05736_);
  nor (_07443_, _07442_, _07042_);
  not (_07444_, _07443_);
  nor (_07445_, _07444_, _07441_);
  and (_07446_, _07042_, _05983_);
  nor (_07447_, _07446_, _05732_);
  not (_07448_, _07447_);
  nor (_07449_, _07448_, _07445_);
  and (_07450_, _07362_, _05732_);
  nor (_07451_, _07450_, _07051_);
  not (_07452_, _07451_);
  nor (_07453_, _07452_, _07449_);
  and (_07454_, _07353_, _07051_);
  nor (_07455_, _07454_, _07050_);
  not (_07456_, _07455_);
  nor (_07457_, _07456_, _07453_);
  not (_07458_, _07059_);
  and (_07459_, _07050_, _06299_);
  nor (_07460_, _07459_, _07458_);
  not (_07461_, _07460_);
  nor (_07462_, _07461_, _07457_);
  nor (_07463_, _07362_, _07059_);
  nor (_07464_, _07463_, _07058_);
  not (_07465_, _07464_);
  nor (_07466_, _07465_, _07462_);
  and (_07467_, _07058_, _07414_);
  nor (_07468_, _07467_, _07068_);
  not (_07469_, _07468_);
  nor (_07470_, _07469_, _07466_);
  and (_07471_, _07353_, _07068_);
  nor (_07472_, _07471_, _07067_);
  not (_07473_, _07472_);
  nor (_07474_, _07473_, _07470_);
  nor (_07475_, _06048_, _05984_);
  nor (_07476_, _07475_, _07474_);
  not (_07477_, _06403_);
  and (_07478_, _07067_, _07477_);
  and (_07479_, _06360_, _05652_);
  nor (_07480_, _07356_, \oc8051_golden_model_1.SP [2]);
  nor (_07481_, _07480_, _07357_);
  and (_07482_, _07481_, _05732_);
  and (_07483_, _07477_, _06021_);
  nor (_07484_, _07481_, _05686_);
  and (_07485_, _06976_, _07477_);
  nand (_07486_, _06881_, \oc8051_golden_model_1.IRAM[0] [2]);
  nand (_07487_, _06726_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_07488_, _07487_, _06879_);
  nand (_07489_, _07488_, _07486_);
  nand (_07490_, _06726_, \oc8051_golden_model_1.IRAM[3] [2]);
  nand (_07491_, _06881_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_07492_, _07491_, _06887_);
  nand (_07493_, _07492_, _07490_);
  nand (_07494_, _07493_, _07489_);
  nand (_07495_, _07494_, _06504_);
  nand (_07496_, _06726_, \oc8051_golden_model_1.IRAM[7] [2]);
  nand (_07497_, _06881_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_07498_, _07497_, _06887_);
  nand (_07499_, _07498_, _07496_);
  nand (_07500_, _06881_, \oc8051_golden_model_1.IRAM[4] [2]);
  nand (_07501_, _06726_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_07502_, _07501_, _06879_);
  nand (_07503_, _07502_, _07500_);
  nand (_07504_, _07503_, _07499_);
  nand (_07505_, _07504_, _06894_);
  nand (_07506_, _07505_, _07495_);
  nand (_07507_, _07506_, _06328_);
  nand (_07508_, _06726_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_07509_, _06881_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_07510_, _07509_, _06887_);
  nand (_07511_, _07510_, _07508_);
  nand (_07512_, _06881_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_07513_, _06726_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_07514_, _07513_, _06879_);
  nand (_07515_, _07514_, _07512_);
  nand (_07516_, _07515_, _07511_);
  nand (_07517_, _07516_, _06504_);
  nand (_07518_, _06726_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_07519_, _06881_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_07520_, _07519_, _06887_);
  nand (_07521_, _07520_, _07518_);
  nand (_07522_, _06881_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_07523_, _06726_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_07524_, _07523_, _06879_);
  nand (_07525_, _07524_, _07522_);
  nand (_07526_, _07525_, _07521_);
  nand (_07527_, _07526_, _06894_);
  nand (_07528_, _07527_, _07517_);
  nand (_07529_, _07528_, _06908_);
  nand (_07530_, _07529_, _07507_);
  or (_07531_, _07530_, _05670_);
  and (_07532_, _07531_, _07247_);
  and (_07533_, _06940_, _06403_);
  nor (_07534_, _07533_, _07532_);
  not (_07535_, _07481_);
  and (_07536_, _07535_, _06943_);
  and (_07537_, _06095_, _06042_);
  nor (_07538_, _07537_, _07536_);
  and (_07539_, _07538_, _07534_);
  and (_07540_, _07530_, _06948_);
  nor (_07541_, _07540_, _06955_);
  and (_07542_, _07541_, _07539_);
  and (_07543_, _06955_, _07477_);
  nor (_07544_, _07543_, _07542_);
  and (_07545_, _06953_, _06359_);
  nor (_07546_, _07545_, _07544_);
  or (_07547_, _07481_, _05690_);
  nand (_07548_, _07547_, _07546_);
  and (_07549_, _06095_, _06037_);
  and (_07550_, _06963_, _06403_);
  nor (_07551_, _07550_, _07549_);
  not (_07552_, _07551_);
  nor (_07553_, _07552_, _07548_);
  and (_07554_, _07530_, _06970_);
  nor (_07555_, _07554_, _06976_);
  and (_07556_, _07555_, _07553_);
  nor (_07557_, _07556_, _07485_);
  nor (_07558_, _07557_, _06975_);
  nor (_07559_, _07558_, _06371_);
  nor (_07560_, _07559_, _06038_);
  and (_07561_, _07481_, _06038_);
  nor (_07562_, _07561_, _07560_);
  and (_07563_, _06035_, _06359_);
  nor (_07564_, _07563_, _07562_);
  nand (_07565_, _07564_, _06232_);
  nor (_07566_, _07565_, _07484_);
  and (_07567_, _07530_, _06992_);
  not (_07568_, _07567_);
  and (_07569_, _07568_, _07566_);
  and (_07570_, _06991_, _06359_);
  nor (_07571_, _07570_, _06023_);
  and (_07572_, _07571_, _07569_);
  nor (_07573_, _07535_, _05673_);
  nor (_07574_, _07573_, _07572_);
  nor (_07575_, _07015_, _07477_);
  nor (_07576_, _07575_, _07252_);
  not (_07577_, _07576_);
  nor (_07578_, _07577_, _07574_);
  and (_07579_, _07530_, _07023_);
  nor (_07580_, _07579_, _06021_);
  and (_07581_, _07580_, _07578_);
  nor (_07582_, _07581_, _07483_);
  nor (_07583_, _07582_, _05724_);
  and (_07584_, _07481_, _05724_);
  nor (_07585_, _07584_, _07583_);
  nor (_07586_, _07035_, _07477_);
  nor (_07587_, _07586_, _05736_);
  not (_07588_, _07587_);
  nor (_07589_, _07588_, _07585_);
  and (_07590_, _07481_, _05736_);
  nor (_07591_, _07590_, _07589_);
  and (_07592_, _07042_, _06403_);
  nor (_07593_, _07592_, _05732_);
  not (_07594_, _07593_);
  nor (_07595_, _07594_, _07591_);
  nor (_07596_, _07595_, _07482_);
  and (_07597_, _06095_, _05495_);
  nor (_07598_, _07597_, _07596_);
  and (_07599_, _07530_, _07051_);
  nor (_07600_, _07599_, _07050_);
  and (_07601_, _07600_, _07598_);
  and (_07602_, _07050_, _07477_);
  nor (_07603_, _07602_, _07601_);
  nor (_07604_, _07481_, _07059_);
  nor (_07605_, _07604_, _07058_);
  not (_07606_, _07605_);
  nor (_07607_, _07606_, _07603_);
  nor (_07608_, _07607_, _07479_);
  and (_07609_, _06095_, _05750_);
  nor (_07610_, _07609_, _07608_);
  and (_07611_, _07530_, _07068_);
  nor (_07612_, _07611_, _07067_);
  and (_07613_, _07612_, _07610_);
  nor (_07614_, _07613_, _07478_);
  nor (_07615_, _07614_, _07305_);
  not (_07616_, _07615_);
  nor (_07617_, _07616_, _07476_);
  and (_07618_, _07617_, _07307_);
  or (_07619_, _07618_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_07620_, _07359_, _06029_);
  nor (_07621_, _07481_, _07081_);
  nor (_07622_, _07621_, _07620_);
  and (_07623_, _07360_, _06029_);
  nor (_07624_, _07620_, _07362_);
  nor (_07625_, _07624_, _07623_);
  and (_07626_, _07234_, _07235_);
  and (_07627_, _07626_, _07274_);
  nor (_07628_, _07627_, _07230_);
  and (_07629_, _07628_, _07625_);
  and (_07630_, _07629_, _07622_);
  and (_07631_, _07630_, _07080_);
  not (_07632_, _07631_);
  and (_07633_, _07632_, _07619_);
  not (_07634_, _07618_);
  and (_07635_, _06084_, _05952_);
  and (_07636_, _07635_, _06359_);
  and (_07637_, _07636_, _06758_);
  and (_07638_, _07637_, _05983_);
  nor (_07639_, _06799_, _06016_);
  and (_07640_, _07639_, _07477_);
  and (_07641_, _07640_, _07638_);
  and (_07642_, _07641_, \oc8051_golden_model_1.PCON [7]);
  not (_07643_, _07642_);
  and (_07644_, _06799_, _06016_);
  not (_07645_, _07644_);
  nand (_07646_, _06403_, _06299_);
  nor (_07647_, _07646_, _07645_);
  and (_07648_, _07647_, _07637_);
  and (_07649_, _07648_, \oc8051_golden_model_1.TCON [7]);
  and (_07650_, _06799_, _06017_);
  not (_07651_, _07650_);
  nor (_07652_, _07651_, _07646_);
  and (_07653_, _07652_, _07637_);
  and (_07654_, _07653_, \oc8051_golden_model_1.TMOD [7]);
  not (_07655_, _07637_);
  nor (_07656_, _06799_, _06017_);
  not (_07657_, _07656_);
  or (_07658_, _07657_, _07646_);
  nor (_07659_, _07658_, _07655_);
  and (_07660_, _07659_, \oc8051_golden_model_1.TL0 [7]);
  or (_07661_, _06403_, _05983_);
  or (_07662_, _07661_, _07645_);
  nor (_07663_, _07662_, _07655_);
  and (_07664_, _07663_, \oc8051_golden_model_1.TH0 [7]);
  not (_07665_, _07639_);
  or (_07666_, _07665_, _07646_);
  nor (_07667_, _07666_, _07655_);
  and (_07668_, _07667_, \oc8051_golden_model_1.TL1 [7]);
  or (_07669_, _07661_, _07651_);
  nor (_07670_, _07669_, _07655_);
  and (_07671_, _07670_, \oc8051_golden_model_1.TH1 [7]);
  nand (_07672_, _06403_, _05983_);
  nor (_07673_, _07672_, _07645_);
  not (_07674_, _06758_);
  and (_07675_, _07674_, _06359_);
  and (_07676_, _07675_, _07635_);
  and (_07677_, _07676_, _07673_);
  and (_07678_, _07677_, \oc8051_golden_model_1.P1 [7]);
  and (_07679_, _07676_, _07647_);
  and (_07680_, _07679_, \oc8051_golden_model_1.SCON [7]);
  and (_07681_, _07652_, _07676_);
  and (_07682_, _07681_, \oc8051_golden_model_1.SBUF [7]);
  not (_07683_, _06359_);
  and (_07684_, _06758_, _07683_);
  and (_07685_, _07635_, _07684_);
  and (_07686_, _07685_, _07673_);
  and (_07687_, _07686_, \oc8051_golden_model_1.P2 [7]);
  and (_07688_, _07647_, _07685_);
  and (_07689_, _07688_, \oc8051_golden_model_1.IE [7]);
  nor (_07690_, _06758_, _06359_);
  and (_07691_, _07635_, _07690_);
  and (_07692_, _07691_, _07673_);
  and (_07693_, _07692_, \oc8051_golden_model_1.P3 [7]);
  and (_07694_, _07647_, _07691_);
  and (_07695_, _07694_, \oc8051_golden_model_1.IP [7]);
  nor (_07696_, _06084_, _06053_);
  and (_07697_, _07696_, _07690_);
  and (_07698_, _07697_, _07673_);
  and (_07699_, _07698_, \oc8051_golden_model_1.B [7]);
  and (_07700_, _07684_, _07696_);
  and (_07701_, _07700_, _07673_);
  and (_07702_, _07701_, \oc8051_golden_model_1.ACC [7]);
  nor (_07703_, _07702_, _07699_);
  and (_07704_, _07675_, _07696_);
  and (_07705_, _07704_, _07673_);
  and (_07706_, _07705_, \oc8051_golden_model_1.PSW [7]);
  not (_07707_, _07706_);
  nand (_07708_, _07707_, _07703_);
  or (_07709_, _07708_, _07695_);
  or (_07710_, _07709_, _07693_);
  or (_07711_, _07710_, _07689_);
  or (_07712_, _07711_, _07687_);
  or (_07713_, _07712_, _07682_);
  or (_07714_, _07713_, _07680_);
  or (_07715_, _07714_, _07678_);
  or (_07716_, _07715_, _07671_);
  or (_07717_, _07716_, _07668_);
  or (_07718_, _07717_, _07664_);
  or (_07719_, _07718_, _07660_);
  or (_07720_, _07719_, _07654_);
  nor (_07721_, _07720_, _07649_);
  and (_07722_, _07721_, _07643_);
  and (_07723_, _07639_, _06403_);
  and (_07724_, _07723_, _07638_);
  and (_07725_, _07724_, \oc8051_golden_model_1.DPH [7]);
  and (_07726_, _07650_, _06403_);
  and (_07727_, _07726_, _07638_);
  and (_07728_, _07727_, \oc8051_golden_model_1.SP [7]);
  nor (_07729_, _07728_, _07725_);
  and (_07730_, _07637_, _07673_);
  and (_07731_, _07730_, \oc8051_golden_model_1.P0 [7]);
  and (_07732_, _07656_, _06403_);
  and (_07733_, _07732_, _07638_);
  and (_07734_, _07733_, \oc8051_golden_model_1.DPL [7]);
  nor (_07735_, _07734_, _07731_);
  and (_07736_, _07735_, _07729_);
  and (_07737_, _07736_, _07722_);
  not (_07738_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_07739_, _06726_, _07738_);
  not (_07740_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_07741_, _06881_, _07740_);
  and (_07742_, _07741_, _06879_);
  nand (_07743_, _07742_, _07739_);
  nand (_07744_, _06726_, \oc8051_golden_model_1.IRAM[3] [7]);
  nand (_07745_, _06881_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_07746_, _07745_, _06887_);
  nand (_07747_, _07746_, _07744_);
  nand (_07748_, _07747_, _07743_);
  nand (_07749_, _07748_, _06504_);
  nand (_07750_, _06726_, \oc8051_golden_model_1.IRAM[7] [7]);
  not (_07751_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_07752_, _06726_, _07751_);
  and (_07753_, _07752_, _06887_);
  nand (_07754_, _07753_, _07750_);
  nand (_07755_, _06881_, \oc8051_golden_model_1.IRAM[4] [7]);
  nand (_07756_, _06726_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_07757_, _07756_, _06879_);
  nand (_07758_, _07757_, _07755_);
  nand (_07759_, _07758_, _07754_);
  nand (_07760_, _07759_, _06894_);
  nand (_07761_, _07760_, _07749_);
  nand (_07762_, _07761_, _06328_);
  nand (_07763_, _06726_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand (_07764_, _06881_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_07765_, _07764_, _06887_);
  nand (_07766_, _07765_, _07763_);
  nand (_07767_, _06881_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_07768_, _06726_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_07769_, _07768_, _06879_);
  nand (_07770_, _07769_, _07767_);
  nand (_07771_, _07770_, _07766_);
  nand (_07772_, _07771_, _06504_);
  nand (_07773_, _06726_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_07774_, _06881_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_07775_, _07774_, _06887_);
  nand (_07776_, _07775_, _07773_);
  nand (_07777_, _06881_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand (_07778_, _06726_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_07779_, _07778_, _06879_);
  nand (_07780_, _07779_, _07777_);
  nand (_07781_, _07780_, _07776_);
  nand (_07782_, _07781_, _06894_);
  nand (_07783_, _07782_, _07772_);
  nand (_07784_, _07783_, _06908_);
  nand (_07785_, _07784_, _07762_);
  or (_07786_, _07785_, _05952_);
  and (_07787_, _07786_, _07737_);
  not (_07788_, _07787_);
  and (_07789_, _07686_, \oc8051_golden_model_1.P2 [6]);
  not (_07790_, _07789_);
  and (_07791_, _07681_, \oc8051_golden_model_1.SBUF [6]);
  not (_07792_, _07791_);
  and (_07793_, _07688_, \oc8051_golden_model_1.IE [6]);
  and (_07794_, _07692_, \oc8051_golden_model_1.P3 [6]);
  nor (_07795_, _07794_, _07793_);
  and (_07796_, _07795_, _07792_);
  and (_07797_, _07796_, _07790_);
  and (_07798_, _07730_, \oc8051_golden_model_1.P0 [6]);
  not (_07799_, _07798_);
  and (_07800_, _07733_, \oc8051_golden_model_1.DPL [6]);
  nor (_07801_, _07665_, _07672_);
  and (_07802_, _07801_, _07637_);
  and (_07803_, _07802_, \oc8051_golden_model_1.DPH [6]);
  nor (_07804_, _07803_, _07800_);
  and (_07805_, _07804_, _07799_);
  and (_07806_, _07667_, \oc8051_golden_model_1.TL1 [6]);
  and (_07807_, _07670_, \oc8051_golden_model_1.TH1 [6]);
  nor (_07808_, _07807_, _07806_);
  and (_07809_, _07679_, \oc8051_golden_model_1.SCON [6]);
  and (_07810_, _07677_, \oc8051_golden_model_1.P1 [6]);
  nor (_07811_, _07810_, _07809_);
  and (_07812_, _07811_, _07808_);
  and (_07813_, _07812_, _07805_);
  and (_07814_, _07813_, _07797_);
  and (_07815_, _07694_, \oc8051_golden_model_1.IP [6]);
  not (_07816_, _07815_);
  and (_07817_, _07698_, \oc8051_golden_model_1.B [6]);
  and (_07818_, _07701_, \oc8051_golden_model_1.ACC [6]);
  nor (_07819_, _07818_, _07817_);
  and (_07820_, _07819_, _07816_);
  and (_07821_, _07641_, \oc8051_golden_model_1.PCON [6]);
  and (_07822_, _07705_, \oc8051_golden_model_1.PSW [6]);
  nor (_07823_, _07822_, _07821_);
  and (_07824_, _07823_, _07820_);
  and (_07825_, _07653_, \oc8051_golden_model_1.TMOD [6]);
  not (_07826_, _07825_);
  and (_07827_, _07659_, \oc8051_golden_model_1.TL0 [6]);
  and (_07828_, _07663_, \oc8051_golden_model_1.TH0 [6]);
  nor (_07829_, _07828_, _07827_);
  and (_07830_, _07829_, _07826_);
  and (_07831_, _07648_, \oc8051_golden_model_1.TCON [6]);
  or (_07832_, _07651_, _07672_);
  nor (_07833_, _07832_, _07655_);
  and (_07834_, _07833_, \oc8051_golden_model_1.SP [6]);
  nor (_07835_, _07834_, _07831_);
  and (_07836_, _07835_, _07830_);
  and (_07837_, _07836_, _07824_);
  and (_07838_, _07837_, _07814_);
  nand (_07839_, _06881_, \oc8051_golden_model_1.IRAM[0] [6]);
  nand (_07840_, _06726_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_07841_, _07840_, _06879_);
  nand (_07842_, _07841_, _07839_);
  nand (_07843_, _06726_, \oc8051_golden_model_1.IRAM[3] [6]);
  nand (_07844_, _06881_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_07845_, _07844_, _06887_);
  nand (_07846_, _07845_, _07843_);
  nand (_07847_, _07846_, _07842_);
  nand (_07848_, _07847_, _06504_);
  nand (_07849_, _06726_, \oc8051_golden_model_1.IRAM[7] [6]);
  nand (_07850_, _06881_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_07851_, _07850_, _06887_);
  nand (_07852_, _07851_, _07849_);
  nand (_07853_, _06881_, \oc8051_golden_model_1.IRAM[4] [6]);
  nand (_07854_, _06726_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_07855_, _07854_, _06879_);
  nand (_07856_, _07855_, _07853_);
  nand (_07857_, _07856_, _07852_);
  nand (_07858_, _07857_, _06894_);
  nand (_07859_, _07858_, _07848_);
  nand (_07860_, _07859_, _06328_);
  nand (_07861_, _06726_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_07862_, _06881_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_07863_, _07862_, _06887_);
  nand (_07864_, _07863_, _07861_);
  nand (_07865_, _06881_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_07866_, _06726_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_07867_, _07866_, _06879_);
  nand (_07868_, _07867_, _07865_);
  nand (_07869_, _07868_, _07864_);
  nand (_07870_, _07869_, _06504_);
  nand (_07871_, _06726_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_07872_, _06881_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_07873_, _07872_, _06887_);
  nand (_07874_, _07873_, _07871_);
  nand (_07875_, _06881_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_07876_, _06726_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_07877_, _07876_, _06879_);
  nand (_07878_, _07877_, _07875_);
  nand (_07879_, _07878_, _07874_);
  nand (_07880_, _07879_, _06894_);
  nand (_07881_, _07880_, _07870_);
  nand (_07882_, _07881_, _06908_);
  nand (_07883_, _07882_, _07860_);
  or (_07884_, _07883_, _05952_);
  and (_07885_, _07884_, _07838_);
  not (_07886_, _07885_);
  and (_07887_, _07686_, \oc8051_golden_model_1.P2 [5]);
  not (_07888_, _07887_);
  and (_07889_, _07681_, \oc8051_golden_model_1.SBUF [5]);
  not (_07890_, _07889_);
  and (_07891_, _07688_, \oc8051_golden_model_1.IE [5]);
  and (_07892_, _07692_, \oc8051_golden_model_1.P3 [5]);
  nor (_07893_, _07892_, _07891_);
  and (_07894_, _07893_, _07890_);
  and (_07895_, _07894_, _07888_);
  and (_07896_, _07667_, \oc8051_golden_model_1.TL1 [5]);
  and (_07897_, _07670_, \oc8051_golden_model_1.TH1 [5]);
  nor (_07898_, _07897_, _07896_);
  and (_07899_, _07679_, \oc8051_golden_model_1.SCON [5]);
  and (_07900_, _07677_, \oc8051_golden_model_1.P1 [5]);
  nor (_07901_, _07900_, _07899_);
  and (_07902_, _07901_, _07898_);
  and (_07903_, _07902_, _07895_);
  and (_07904_, _07694_, \oc8051_golden_model_1.IP [5]);
  not (_07905_, _07904_);
  and (_07906_, _07698_, \oc8051_golden_model_1.B [5]);
  and (_07907_, _07701_, \oc8051_golden_model_1.ACC [5]);
  nor (_07908_, _07907_, _07906_);
  and (_07909_, _07908_, _07905_);
  and (_07910_, _07641_, \oc8051_golden_model_1.PCON [5]);
  and (_07911_, _07705_, \oc8051_golden_model_1.PSW [5]);
  nor (_07912_, _07911_, _07910_);
  and (_07913_, _07912_, _07909_);
  and (_07914_, _07648_, \oc8051_golden_model_1.TCON [5]);
  not (_07915_, _07914_);
  and (_07916_, _07663_, \oc8051_golden_model_1.TH0 [5]);
  and (_07917_, _07659_, \oc8051_golden_model_1.TL0 [5]);
  nor (_07918_, _07917_, _07916_);
  and (_07919_, _07918_, _07915_);
  and (_07920_, _07653_, \oc8051_golden_model_1.TMOD [5]);
  not (_07921_, _07920_);
  and (_07922_, _07733_, \oc8051_golden_model_1.DPL [5]);
  and (_07923_, _07802_, \oc8051_golden_model_1.DPH [5]);
  nor (_07924_, _07923_, _07922_);
  and (_07925_, _07730_, \oc8051_golden_model_1.P0 [5]);
  and (_07926_, _07833_, \oc8051_golden_model_1.SP [5]);
  nor (_07927_, _07926_, _07925_);
  and (_07928_, _07927_, _07924_);
  and (_07929_, _07928_, _07921_);
  and (_07930_, _07929_, _07919_);
  and (_07931_, _07930_, _07913_);
  and (_07932_, _07931_, _07903_);
  nand (_07933_, _06881_, \oc8051_golden_model_1.IRAM[0] [5]);
  nand (_07934_, _06726_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_07935_, _07934_, _06879_);
  nand (_07936_, _07935_, _07933_);
  nand (_07937_, _06726_, \oc8051_golden_model_1.IRAM[3] [5]);
  nand (_07938_, _06881_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_07939_, _07938_, _06887_);
  nand (_07940_, _07939_, _07937_);
  nand (_07941_, _07940_, _07936_);
  nand (_07942_, _07941_, _06504_);
  nand (_07943_, _06726_, \oc8051_golden_model_1.IRAM[7] [5]);
  nand (_07944_, _06881_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_07945_, _07944_, _06887_);
  nand (_07946_, _07945_, _07943_);
  nand (_07947_, _06881_, \oc8051_golden_model_1.IRAM[4] [5]);
  nand (_07948_, _06726_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_07949_, _07948_, _06879_);
  nand (_07950_, _07949_, _07947_);
  nand (_07951_, _07950_, _07946_);
  nand (_07952_, _07951_, _06894_);
  nand (_07953_, _07952_, _07942_);
  nand (_07954_, _07953_, _06328_);
  nand (_07955_, _06726_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_07956_, _06881_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_07957_, _07956_, _06887_);
  nand (_07958_, _07957_, _07955_);
  nand (_07959_, _06881_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_07960_, _06726_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_07961_, _07960_, _06879_);
  nand (_07962_, _07961_, _07959_);
  nand (_07963_, _07962_, _07958_);
  nand (_07964_, _07963_, _06504_);
  nand (_07965_, _06726_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_07966_, _06881_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_07967_, _07966_, _06887_);
  nand (_07968_, _07967_, _07965_);
  nand (_07969_, _06881_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand (_07970_, _06726_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_07971_, _07970_, _06879_);
  nand (_07972_, _07971_, _07969_);
  nand (_07973_, _07972_, _07968_);
  nand (_07974_, _07973_, _06894_);
  nand (_07975_, _07974_, _07964_);
  nand (_07976_, _07975_, _06908_);
  nand (_07977_, _07976_, _07954_);
  or (_07978_, _07977_, _05952_);
  and (_07979_, _07978_, _07932_);
  not (_07980_, _07979_);
  and (_07981_, _07667_, \oc8051_golden_model_1.TL1 [3]);
  not (_07982_, _07981_);
  and (_07983_, _07677_, \oc8051_golden_model_1.P1 [3]);
  and (_07984_, _07679_, \oc8051_golden_model_1.SCON [3]);
  nor (_07985_, _07984_, _07983_);
  and (_07986_, _07985_, _07982_);
  and (_07987_, _07681_, \oc8051_golden_model_1.SBUF [3]);
  not (_07988_, _07987_);
  and (_07989_, _07692_, \oc8051_golden_model_1.P3 [3]);
  and (_07990_, _07688_, \oc8051_golden_model_1.IE [3]);
  nor (_07991_, _07990_, _07989_);
  and (_07992_, _07991_, _07988_);
  and (_07993_, _07686_, \oc8051_golden_model_1.P2 [3]);
  and (_07994_, _07670_, \oc8051_golden_model_1.TH1 [3]);
  nor (_07995_, _07994_, _07993_);
  and (_07996_, _07995_, _07992_);
  and (_07997_, _07996_, _07986_);
  and (_07998_, _07694_, \oc8051_golden_model_1.IP [3]);
  not (_07999_, _07998_);
  and (_08000_, _07701_, \oc8051_golden_model_1.ACC [3]);
  and (_08001_, _07698_, \oc8051_golden_model_1.B [3]);
  nor (_08002_, _08001_, _08000_);
  and (_08003_, _08002_, _07999_);
  and (_08004_, _07641_, \oc8051_golden_model_1.PCON [3]);
  and (_08005_, _07705_, \oc8051_golden_model_1.PSW [3]);
  nor (_08006_, _08005_, _08004_);
  and (_08007_, _08006_, _08003_);
  and (_08008_, _07653_, \oc8051_golden_model_1.TMOD [3]);
  not (_08009_, _08008_);
  and (_08010_, _07663_, \oc8051_golden_model_1.TH0 [3]);
  and (_08011_, _07659_, \oc8051_golden_model_1.TL0 [3]);
  nor (_08012_, _08011_, _08010_);
  and (_08013_, _08012_, _08009_);
  and (_08014_, _07648_, \oc8051_golden_model_1.TCON [3]);
  not (_08015_, _08014_);
  and (_08016_, _07733_, \oc8051_golden_model_1.DPL [3]);
  and (_08017_, _07802_, \oc8051_golden_model_1.DPH [3]);
  nor (_08018_, _08017_, _08016_);
  and (_08019_, _07730_, \oc8051_golden_model_1.P0 [3]);
  and (_08020_, _07833_, \oc8051_golden_model_1.SP [3]);
  nor (_08021_, _08020_, _08019_);
  and (_08022_, _08021_, _08018_);
  and (_08023_, _08022_, _08015_);
  and (_08024_, _08023_, _08013_);
  and (_08025_, _08024_, _08007_);
  and (_08026_, _08025_, _07997_);
  or (_08027_, _07353_, _05952_);
  and (_08028_, _08027_, _08026_);
  not (_08029_, _08028_);
  and (_08030_, _07670_, \oc8051_golden_model_1.TH1 [1]);
  not (_08031_, _08030_);
  and (_08032_, _07679_, \oc8051_golden_model_1.SCON [1]);
  and (_08033_, _07677_, \oc8051_golden_model_1.P1 [1]);
  nor (_08034_, _08033_, _08032_);
  and (_08035_, _08034_, _08031_);
  and (_08036_, _07681_, \oc8051_golden_model_1.SBUF [1]);
  not (_08037_, _08036_);
  and (_08038_, _07692_, \oc8051_golden_model_1.P3 [1]);
  and (_08039_, _07688_, \oc8051_golden_model_1.IE [1]);
  nor (_08040_, _08039_, _08038_);
  and (_08041_, _08040_, _08037_);
  and (_08042_, _07686_, \oc8051_golden_model_1.P2 [1]);
  and (_08043_, _07667_, \oc8051_golden_model_1.TL1 [1]);
  nor (_08044_, _08043_, _08042_);
  and (_08045_, _08044_, _08041_);
  and (_08046_, _08045_, _08035_);
  and (_08047_, _07694_, \oc8051_golden_model_1.IP [1]);
  not (_08048_, _08047_);
  and (_08049_, _07701_, \oc8051_golden_model_1.ACC [1]);
  and (_08050_, _07698_, \oc8051_golden_model_1.B [1]);
  nor (_08051_, _08050_, _08049_);
  and (_08052_, _08051_, _08048_);
  and (_08053_, _07641_, \oc8051_golden_model_1.PCON [1]);
  and (_08054_, _07705_, \oc8051_golden_model_1.PSW [1]);
  nor (_08055_, _08054_, _08053_);
  and (_08056_, _08055_, _08052_);
  and (_08057_, _07653_, \oc8051_golden_model_1.TMOD [1]);
  not (_08058_, _08057_);
  and (_08059_, _07659_, \oc8051_golden_model_1.TL0 [1]);
  and (_08060_, _07663_, \oc8051_golden_model_1.TH0 [1]);
  nor (_08061_, _08060_, _08059_);
  and (_08062_, _08061_, _08058_);
  and (_08063_, _07648_, \oc8051_golden_model_1.TCON [1]);
  not (_08064_, _08063_);
  and (_08065_, _07730_, \oc8051_golden_model_1.P0 [1]);
  and (_08066_, _07833_, \oc8051_golden_model_1.SP [1]);
  nor (_08067_, _08066_, _08065_);
  and (_08068_, _07733_, \oc8051_golden_model_1.DPL [1]);
  and (_08069_, _07802_, \oc8051_golden_model_1.DPH [1]);
  nor (_08070_, _08069_, _08068_);
  and (_08071_, _08070_, _08067_);
  and (_08072_, _08071_, _08064_);
  and (_08073_, _08072_, _08062_);
  and (_08074_, _08073_, _08056_);
  and (_08075_, _08074_, _08046_);
  or (_08076_, _07132_, _05952_);
  and (_08077_, _08076_, _08075_);
  not (_08078_, _08077_);
  and (_08079_, _07681_, \oc8051_golden_model_1.SBUF [0]);
  not (_08080_, _08079_);
  and (_08081_, _07686_, \oc8051_golden_model_1.P2 [0]);
  not (_08082_, _08081_);
  and (_08083_, _07692_, \oc8051_golden_model_1.P3 [0]);
  and (_08084_, _07688_, \oc8051_golden_model_1.IE [0]);
  nor (_08085_, _08084_, _08083_);
  and (_08086_, _08085_, _08082_);
  and (_08087_, _08086_, _08080_);
  and (_08088_, _07833_, \oc8051_golden_model_1.SP [0]);
  not (_08089_, _08088_);
  and (_08090_, _07733_, \oc8051_golden_model_1.DPL [0]);
  and (_08091_, _07802_, \oc8051_golden_model_1.DPH [0]);
  nor (_08092_, _08091_, _08090_);
  and (_08093_, _08092_, _08089_);
  and (_08094_, _07677_, \oc8051_golden_model_1.P1 [0]);
  and (_08095_, _07679_, \oc8051_golden_model_1.SCON [0]);
  nor (_08096_, _08095_, _08094_);
  and (_08097_, _07670_, \oc8051_golden_model_1.TH1 [0]);
  and (_08098_, _07667_, \oc8051_golden_model_1.TL1 [0]);
  nor (_08099_, _08098_, _08097_);
  and (_08100_, _08099_, _08096_);
  and (_08101_, _08100_, _08093_);
  and (_08102_, _08101_, _08087_);
  and (_08103_, _07705_, \oc8051_golden_model_1.PSW [0]);
  not (_08104_, _08103_);
  and (_08105_, _07698_, \oc8051_golden_model_1.B [0]);
  and (_08106_, _07701_, \oc8051_golden_model_1.ACC [0]);
  nor (_08107_, _08106_, _08105_);
  and (_08108_, _08107_, _08104_);
  and (_08109_, _07641_, \oc8051_golden_model_1.PCON [0]);
  and (_08110_, _07694_, \oc8051_golden_model_1.IP [0]);
  nor (_08111_, _08110_, _08109_);
  and (_08112_, _08111_, _08108_);
  and (_08113_, _07653_, \oc8051_golden_model_1.TMOD [0]);
  not (_08114_, _08113_);
  and (_08115_, _07659_, \oc8051_golden_model_1.TL0 [0]);
  and (_08116_, _07663_, \oc8051_golden_model_1.TH0 [0]);
  nor (_08117_, _08116_, _08115_);
  and (_08118_, _08117_, _08114_);
  and (_08119_, _07730_, \oc8051_golden_model_1.P0 [0]);
  and (_08120_, _07648_, \oc8051_golden_model_1.TCON [0]);
  nor (_08121_, _08120_, _08119_);
  and (_08122_, _08121_, _08118_);
  and (_08123_, _08122_, _08112_);
  and (_08124_, _08123_, _08102_);
  not (_08125_, _08124_);
  and (_08126_, _06931_, _06053_);
  or (_08127_, _08126_, _08125_);
  and (_08128_, _08127_, _08078_);
  and (_08129_, _07681_, \oc8051_golden_model_1.SBUF [2]);
  not (_08130_, _08129_);
  and (_08131_, _07692_, \oc8051_golden_model_1.P3 [2]);
  and (_08132_, _07688_, \oc8051_golden_model_1.IE [2]);
  nor (_08133_, _08132_, _08131_);
  and (_08134_, _08133_, _08130_);
  and (_08135_, _07686_, \oc8051_golden_model_1.P2 [2]);
  and (_08136_, _07667_, \oc8051_golden_model_1.TL1 [2]);
  nor (_08137_, _08136_, _08135_);
  and (_08138_, _08137_, _08134_);
  and (_08139_, _07653_, \oc8051_golden_model_1.TMOD [2]);
  not (_08140_, _08139_);
  and (_08141_, _07659_, \oc8051_golden_model_1.TL0 [2]);
  and (_08142_, _07663_, \oc8051_golden_model_1.TH0 [2]);
  nor (_08143_, _08142_, _08141_);
  and (_08144_, _08143_, _08140_);
  and (_08145_, _07730_, \oc8051_golden_model_1.P0 [2]);
  and (_08146_, _07648_, \oc8051_golden_model_1.TCON [2]);
  nor (_08147_, _08146_, _08145_);
  and (_08148_, _08147_, _08144_);
  and (_08149_, _08148_, _08138_);
  and (_08150_, _07705_, \oc8051_golden_model_1.PSW [2]);
  not (_08151_, _08150_);
  and (_08152_, _07698_, \oc8051_golden_model_1.B [2]);
  and (_08153_, _07701_, \oc8051_golden_model_1.ACC [2]);
  nor (_08154_, _08153_, _08152_);
  and (_08155_, _08154_, _08151_);
  and (_08156_, _07641_, \oc8051_golden_model_1.PCON [2]);
  and (_08157_, _07694_, \oc8051_golden_model_1.IP [2]);
  nor (_08158_, _08157_, _08156_);
  and (_08159_, _08158_, _08155_);
  and (_08160_, _07833_, \oc8051_golden_model_1.SP [2]);
  not (_08161_, _08160_);
  and (_08162_, _07733_, \oc8051_golden_model_1.DPL [2]);
  and (_08163_, _07802_, \oc8051_golden_model_1.DPH [2]);
  nor (_08164_, _08163_, _08162_);
  and (_08165_, _08164_, _08161_);
  and (_08166_, _07670_, \oc8051_golden_model_1.TH1 [2]);
  not (_08167_, _08166_);
  and (_08168_, _07677_, \oc8051_golden_model_1.P1 [2]);
  and (_08169_, _07679_, \oc8051_golden_model_1.SCON [2]);
  nor (_08170_, _08169_, _08168_);
  and (_08171_, _08170_, _08167_);
  and (_08172_, _08171_, _08165_);
  and (_08173_, _08172_, _08159_);
  and (_08174_, _08173_, _08149_);
  or (_08175_, _07530_, _05952_);
  and (_08176_, _08175_, _08174_);
  not (_08177_, _08176_);
  and (_08178_, _08177_, _08128_);
  and (_08179_, _08178_, _08029_);
  and (_08180_, _07670_, \oc8051_golden_model_1.TH1 [4]);
  not (_08181_, _08180_);
  and (_08182_, _07679_, \oc8051_golden_model_1.SCON [4]);
  and (_08183_, _07677_, \oc8051_golden_model_1.P1 [4]);
  nor (_08184_, _08183_, _08182_);
  and (_08185_, _08184_, _08181_);
  and (_08186_, _07681_, \oc8051_golden_model_1.SBUF [4]);
  not (_08187_, _08186_);
  and (_08188_, _07688_, \oc8051_golden_model_1.IE [4]);
  and (_08189_, _07692_, \oc8051_golden_model_1.P3 [4]);
  nor (_08190_, _08189_, _08188_);
  and (_08191_, _08190_, _08187_);
  and (_08192_, _07686_, \oc8051_golden_model_1.P2 [4]);
  and (_08193_, _07667_, \oc8051_golden_model_1.TL1 [4]);
  nor (_08194_, _08193_, _08192_);
  and (_08195_, _08194_, _08191_);
  and (_08196_, _08195_, _08185_);
  and (_08197_, _07694_, \oc8051_golden_model_1.IP [4]);
  not (_08198_, _08197_);
  and (_08199_, _07698_, \oc8051_golden_model_1.B [4]);
  and (_08200_, _07701_, \oc8051_golden_model_1.ACC [4]);
  nor (_08201_, _08200_, _08199_);
  and (_08202_, _08201_, _08198_);
  and (_08203_, _07641_, \oc8051_golden_model_1.PCON [4]);
  and (_08204_, _07705_, \oc8051_golden_model_1.PSW [4]);
  nor (_08205_, _08204_, _08203_);
  and (_08206_, _08205_, _08202_);
  and (_08207_, _07648_, \oc8051_golden_model_1.TCON [4]);
  not (_08208_, _08207_);
  and (_08209_, _07659_, \oc8051_golden_model_1.TL0 [4]);
  and (_08210_, _07663_, \oc8051_golden_model_1.TH0 [4]);
  nor (_08211_, _08210_, _08209_);
  and (_08212_, _08211_, _08208_);
  and (_08213_, _07653_, \oc8051_golden_model_1.TMOD [4]);
  not (_08214_, _08213_);
  and (_08215_, _07730_, \oc8051_golden_model_1.P0 [4]);
  and (_08216_, _07833_, \oc8051_golden_model_1.SP [4]);
  nor (_08217_, _08216_, _08215_);
  and (_08218_, _07733_, \oc8051_golden_model_1.DPL [4]);
  and (_08219_, _07802_, \oc8051_golden_model_1.DPH [4]);
  nor (_08220_, _08219_, _08218_);
  and (_08221_, _08220_, _08217_);
  and (_08222_, _08221_, _08214_);
  and (_08223_, _08222_, _08212_);
  and (_08224_, _08223_, _08206_);
  and (_08225_, _08224_, _08196_);
  nand (_08226_, _06881_, \oc8051_golden_model_1.IRAM[0] [4]);
  nand (_08227_, _06726_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_08228_, _08227_, _06879_);
  nand (_08229_, _08228_, _08226_);
  nand (_08230_, _06726_, \oc8051_golden_model_1.IRAM[3] [4]);
  nand (_08231_, _06881_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_08232_, _08231_, _06887_);
  nand (_08233_, _08232_, _08230_);
  nand (_08234_, _08233_, _08229_);
  nand (_08235_, _08234_, _06504_);
  nand (_08236_, _06726_, \oc8051_golden_model_1.IRAM[7] [4]);
  nand (_08237_, _06881_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_08238_, _08237_, _06887_);
  nand (_08239_, _08238_, _08236_);
  nand (_08240_, _06881_, \oc8051_golden_model_1.IRAM[4] [4]);
  nand (_08241_, _06726_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_08242_, _08241_, _06879_);
  nand (_08243_, _08242_, _08240_);
  nand (_08244_, _08243_, _08239_);
  nand (_08245_, _08244_, _06894_);
  nand (_08246_, _08245_, _08235_);
  nand (_08247_, _08246_, _06328_);
  nand (_08248_, _06726_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_08249_, _06881_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_08250_, _08249_, _06887_);
  nand (_08251_, _08250_, _08248_);
  nand (_08252_, _06881_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_08253_, _06726_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_08254_, _08253_, _06879_);
  nand (_08255_, _08254_, _08252_);
  nand (_08256_, _08255_, _08251_);
  nand (_08257_, _08256_, _06504_);
  nand (_08258_, _06726_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_08259_, _06881_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_08260_, _08259_, _06887_);
  nand (_08261_, _08260_, _08258_);
  nand (_08262_, _06881_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand (_08263_, _06726_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_08264_, _08263_, _06879_);
  nand (_08265_, _08264_, _08262_);
  nand (_08266_, _08265_, _08261_);
  nand (_08267_, _08266_, _06894_);
  nand (_08268_, _08267_, _08257_);
  nand (_08269_, _08268_, _06908_);
  nand (_08270_, _08269_, _08247_);
  or (_08271_, _08270_, _05952_);
  and (_08272_, _08271_, _08225_);
  not (_08273_, _08272_);
  and (_08274_, _08273_, _08179_);
  and (_08275_, _08274_, _07980_);
  and (_08276_, _08275_, _07886_);
  nor (_08277_, _08276_, _07788_);
  and (_08278_, _08276_, _07788_);
  nor (_08279_, _08278_, _08277_);
  and (_08280_, _08279_, _07067_);
  nor (_08281_, _06137_, _06723_);
  or (_08282_, _07278_, _06458_);
  not (_08283_, _08282_);
  not (_08284_, _06457_);
  and (_08285_, _06866_, _08284_);
  and (_08286_, _08285_, _08283_);
  and (_08287_, _08286_, _07211_);
  not (_08288_, _07785_);
  and (_08289_, _08270_, _07977_);
  and (_08290_, _07530_, _07353_);
  and (_08291_, _07132_, _07022_);
  and (_08292_, _08291_, _08290_);
  and (_08293_, _08292_, _08289_);
  and (_08294_, _08293_, _07883_);
  or (_08295_, _08294_, _08288_);
  nand (_08296_, _08294_, _08288_);
  and (_08297_, _08296_, _08295_);
  and (_08298_, _08297_, _07211_);
  or (_08299_, _08298_, _08287_);
  not (_08300_, _07031_);
  nor (_08301_, _07032_, _05952_);
  and (_08302_, _06166_, _04200_);
  and (_08303_, _06205_, _04168_);
  nor (_08304_, _08303_, _08302_);
  and (_08305_, _06210_, _04205_);
  and (_08306_, _06197_, _04208_);
  nor (_08307_, _08306_, _08305_);
  and (_08308_, _08307_, _08304_);
  and (_08309_, _06161_, _04155_);
  and (_08310_, _06203_, _04197_);
  nor (_08311_, _08310_, _08309_);
  and (_08312_, _06199_, _04180_);
  and (_08313_, _06187_, _04159_);
  nor (_08314_, _08313_, _08312_);
  and (_08315_, _08314_, _08311_);
  and (_08316_, _08315_, _08308_);
  and (_08317_, _06170_, _04193_);
  and (_08318_, _06185_, _04176_);
  nor (_08319_, _08318_, _08317_);
  and (_08320_, _06208_, _04172_);
  and (_08321_, _06182_, _04122_);
  nor (_08322_, _08321_, _08320_);
  and (_08323_, _08322_, _08319_);
  and (_08324_, _06179_, _04149_);
  and (_08325_, _06194_, _04165_);
  nor (_08326_, _08325_, _08324_);
  and (_08327_, _06175_, _04185_);
  and (_08328_, _06192_, _04190_);
  nor (_08329_, _08328_, _08327_);
  and (_08330_, _08329_, _08326_);
  and (_08331_, _08330_, _08323_);
  and (_08332_, _08331_, _08316_);
  nor (_08333_, _08332_, _07787_);
  and (_08334_, _08333_, _08301_);
  nand (_08335_, _08332_, _06021_);
  and (_08336_, _07638_, \oc8051_golden_model_1.P0 [7]);
  not (_08337_, _05984_);
  nor (_08338_, _06759_, _08337_);
  and (_08339_, _08338_, _06361_);
  and (_08340_, _08339_, _06087_);
  and (_08341_, _08340_, _07637_);
  and (_08342_, _08341_, \oc8051_golden_model_1.TCON [7]);
  not (_08343_, _06087_);
  and (_08344_, _08339_, _08343_);
  and (_08345_, _08344_, _07676_);
  and (_08346_, _08345_, \oc8051_golden_model_1.P1 [7]);
  and (_08347_, _08340_, _07676_);
  and (_08348_, _08347_, \oc8051_golden_model_1.SCON [7]);
  and (_08349_, _08344_, _07685_);
  and (_08350_, _08349_, \oc8051_golden_model_1.P2 [7]);
  and (_08351_, _08340_, _07685_);
  and (_08352_, _08351_, \oc8051_golden_model_1.IE [7]);
  and (_08353_, _08344_, _07691_);
  and (_08354_, _08353_, \oc8051_golden_model_1.P3 [7]);
  and (_08355_, _07704_, _08344_);
  and (_08356_, _08355_, \oc8051_golden_model_1.PSW [7]);
  and (_08357_, _08340_, _07691_);
  and (_08358_, _08357_, \oc8051_golden_model_1.IP [7]);
  and (_08359_, _08344_, _07700_);
  and (_08360_, _08359_, \oc8051_golden_model_1.ACC [7]);
  and (_08361_, _08344_, _07697_);
  and (_08362_, _08361_, \oc8051_golden_model_1.B [7]);
  or (_08363_, _08362_, _08360_);
  or (_08364_, _08363_, _08358_);
  or (_08365_, _08364_, _08356_);
  or (_08366_, _08365_, _08354_);
  or (_08367_, _08366_, _08352_);
  or (_08368_, _08367_, _08350_);
  or (_08369_, _08368_, _08348_);
  or (_08370_, _08369_, _08346_);
  or (_08371_, _08370_, _08342_);
  nor (_08372_, _08371_, _08336_);
  and (_08373_, _08372_, _07786_);
  nor (_08374_, _08373_, _07640_);
  and (_08375_, _07640_, \oc8051_golden_model_1.PSW [7]);
  or (_08376_, _08375_, _08374_);
  and (_08377_, _08376_, _06991_);
  not (_08378_, _06975_);
  or (_08379_, _08374_, _08378_);
  not (_08380_, _06953_);
  not (_08381_, _06955_);
  not (_08382_, _05567_);
  or (_08383_, _05689_, _08382_);
  not (_08384_, _08383_);
  and (_08385_, _08384_, _08297_);
  and (_08386_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_08387_, _08386_, \oc8051_golden_model_1.PC [6]);
  and (_08388_, _08387_, _05850_);
  and (_08389_, _08388_, \oc8051_golden_model_1.PC [7]);
  nor (_08390_, _08388_, \oc8051_golden_model_1.PC [7]);
  nor (_08391_, _08390_, _08389_);
  and (_08392_, _08391_, _06943_);
  not (_08393_, \oc8051_golden_model_1.ACC [7]);
  nor (_08394_, _06943_, _08393_);
  or (_08395_, _08394_, _08392_);
  and (_08396_, _08395_, _08383_);
  or (_08397_, _08396_, _08385_);
  and (_08398_, _08397_, _06949_);
  nor (_08399_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_08400_, _08399_, _06447_);
  nor (_08401_, _08400_, _06238_);
  nor (_08402_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_08403_, _08402_, _06238_);
  and (_08404_, _08403_, _06029_);
  nor (_08405_, _08404_, _08401_);
  nor (_08406_, _08405_, _06448_);
  not (_08407_, _08406_);
  nand (_08408_, _07353_, _06993_);
  not (_08409_, _06448_);
  and (_08410_, _06992_, _05983_);
  nor (_08411_, _08410_, _08409_);
  nand (_08412_, _08411_, _08408_);
  and (_08413_, _08412_, _08407_);
  nor (_08414_, _08399_, _06447_);
  nor (_08415_, _08414_, _08400_);
  nor (_08416_, _08415_, _06448_);
  not (_08417_, _08416_);
  nand (_08418_, _07530_, _06993_);
  and (_08419_, _06992_, _06403_);
  nor (_08420_, _08419_, _08409_);
  nand (_08421_, _08420_, _08418_);
  and (_08422_, _08421_, _08417_);
  nor (_08423_, _07132_, _06992_);
  nor (_08424_, _06993_, _06799_);
  or (_08425_, _08424_, _08423_);
  nand (_08426_, _08425_, _06448_);
  nor (_08427_, _07083_, _06448_);
  not (_08428_, _08427_);
  and (_08429_, _08428_, _08426_);
  or (_08430_, _06992_, _06931_);
  and (_08431_, _06992_, _06016_);
  nor (_08432_, _08431_, _08409_);
  nand (_08433_, _08432_, _08430_);
  nor (_08434_, _06448_, \oc8051_golden_model_1.SP [0]);
  not (_08435_, _08434_);
  and (_08436_, _08435_, _08433_);
  or (_08437_, _08436_, _07740_);
  nand (_08438_, _08435_, _08433_);
  or (_08439_, _08438_, _07738_);
  nand (_08440_, _08439_, _08437_);
  and (_08441_, _08440_, _08429_);
  or (_08442_, _08438_, \oc8051_golden_model_1.IRAM[2] [7]);
  nand (_08443_, _08428_, _08426_);
  or (_08444_, _08436_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_08445_, _08444_, _08443_);
  and (_08446_, _08445_, _08442_);
  nor (_08447_, _08446_, _08441_);
  nand (_08448_, _08447_, _08422_);
  not (_08449_, _08422_);
  or (_08450_, _08436_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_08451_, _08438_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_08452_, _08451_, _08429_);
  and (_08453_, _08452_, _08450_);
  or (_08454_, _08438_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_08455_, _08436_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_08456_, _08455_, _08443_);
  and (_08457_, _08456_, _08454_);
  nor (_08458_, _08457_, _08453_);
  nand (_08459_, _08458_, _08449_);
  nand (_08460_, _08459_, _08448_);
  nand (_08461_, _08460_, _08413_);
  not (_08462_, _08413_);
  or (_08463_, _08438_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_08464_, _08436_, \oc8051_golden_model_1.IRAM[9] [7]);
  nand (_08465_, _08464_, _08463_);
  nand (_08466_, _08465_, _08429_);
  or (_08467_, _08438_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_08468_, _08436_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand (_08469_, _08468_, _08467_);
  nand (_08470_, _08469_, _08443_);
  nand (_08471_, _08470_, _08466_);
  nand (_08472_, _08471_, _08422_);
  or (_08473_, _08438_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_08474_, _08436_, \oc8051_golden_model_1.IRAM[13] [7]);
  nand (_08475_, _08474_, _08473_);
  nand (_08476_, _08475_, _08429_);
  or (_08477_, _08438_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_08478_, _08436_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_08479_, _08478_, _08477_);
  nand (_08480_, _08479_, _08443_);
  nand (_08481_, _08480_, _08476_);
  nand (_08482_, _08481_, _08449_);
  nand (_08483_, _08482_, _08472_);
  nand (_08484_, _08483_, _08462_);
  and (_08485_, _08484_, _08461_);
  and (_08486_, _08485_, _06948_);
  or (_08487_, _08486_, _08398_);
  and (_08488_, _08487_, _08381_);
  and (_08489_, _08272_, _07979_);
  not (_08490_, _08127_);
  and (_08491_, _08490_, _08077_);
  and (_08492_, _08176_, _08028_);
  and (_08493_, _08492_, _08491_);
  and (_08494_, _08493_, _08489_);
  and (_08495_, _08494_, _07885_);
  or (_08496_, _08495_, _07788_);
  nand (_08497_, _08495_, _07788_);
  and (_08498_, _08497_, _08496_);
  and (_08499_, _08498_, _06955_);
  or (_08500_, _08499_, _08488_);
  and (_08501_, _08500_, _08380_);
  not (_08502_, _07640_);
  nand (_08503_, _08373_, _08502_);
  and (_08504_, _08503_, _06953_);
  or (_08505_, _08504_, _07272_);
  or (_08506_, _08505_, _08501_);
  nor (_08507_, _08391_, _05690_);
  nor (_08508_, _08507_, _06963_);
  and (_08509_, _08508_, _08506_);
  and (_08510_, _08288_, _06963_);
  or (_08511_, _08510_, _06975_);
  or (_08512_, _08511_, _08509_);
  and (_08513_, _08512_, _08379_);
  or (_08514_, _08513_, _06038_);
  nand (_08515_, _07787_, _06038_);
  and (_08516_, _08515_, _06036_);
  and (_08517_, _08516_, _08514_);
  nor (_08518_, _08373_, _08502_);
  not (_08519_, _08518_);
  and (_08520_, _08519_, _08503_);
  and (_08521_, _08520_, _06035_);
  or (_08522_, _08521_, _08517_);
  and (_08523_, _08522_, _05686_);
  not (_08524_, _08391_);
  or (_08525_, _08524_, _05686_);
  nand (_08526_, _08525_, _06233_);
  or (_08527_, _08526_, _08523_);
  nand (_08528_, _07787_, _06573_);
  and (_08529_, _08528_, _08527_);
  or (_08530_, _08529_, _06992_);
  and (_08531_, _08485_, _06053_);
  nand (_08532_, _07737_, _06992_);
  or (_08533_, _08532_, _08531_);
  and (_08534_, _08533_, _07308_);
  and (_08535_, _08534_, _08530_);
  or (_08536_, _08535_, _08377_);
  and (_08537_, _08536_, _05673_);
  or (_08538_, _08524_, _05673_);
  nand (_08539_, _08538_, _07009_);
  or (_08540_, _08539_, _08537_);
  not (_08541_, _07009_);
  nand (_08542_, _07785_, _08541_);
  and (_08543_, _08542_, _08540_);
  or (_08544_, _08543_, _07013_);
  not (_08545_, _07010_);
  or (_08546_, _08485_, _07231_);
  and (_08547_, _08546_, _08545_);
  and (_08548_, _08547_, _08544_);
  not (_08549_, _08332_);
  nor (_08550_, _08549_, _07785_);
  and (_08551_, _06170_, _04508_);
  and (_08552_, _06166_, _04532_);
  nor (_08553_, _08552_, _08551_);
  and (_08554_, _06161_, _04492_);
  and (_08555_, _06187_, _04503_);
  nor (_08556_, _08555_, _08554_);
  and (_08557_, _08556_, _08553_);
  and (_08558_, _06182_, _04510_);
  and (_08559_, _06205_, _04525_);
  nor (_08560_, _08559_, _08558_);
  and (_08561_, _06197_, _04515_);
  and (_08562_, _06192_, _04505_);
  nor (_08563_, _08562_, _08561_);
  and (_08564_, _08563_, _08560_);
  and (_08565_, _08564_, _08557_);
  and (_08566_, _06199_, _04494_);
  and (_08567_, _06194_, _04521_);
  nor (_08568_, _08567_, _08566_);
  and (_08569_, _06185_, _04513_);
  and (_08570_, _06179_, _04523_);
  nor (_08571_, _08570_, _08569_);
  and (_08572_, _08571_, _08568_);
  and (_08573_, _06210_, _04497_);
  and (_08574_, _06203_, _04530_);
  nor (_08575_, _08574_, _08573_);
  and (_08576_, _06208_, _04499_);
  and (_08577_, _06175_, _04519_);
  nor (_08578_, _08577_, _08576_);
  and (_08579_, _08578_, _08575_);
  and (_08580_, _08579_, _08572_);
  and (_08581_, _08580_, _08565_);
  and (_08582_, _06185_, _04579_);
  and (_08583_, _06208_, _04538_);
  nor (_08584_, _08583_, _08582_);
  and (_08585_, _06197_, _04560_);
  and (_08586_, _06187_, _04552_);
  nor (_08587_, _08586_, _08585_);
  and (_08588_, _08587_, _08584_);
  and (_08589_, _06205_, _04568_);
  and (_08590_, _06194_, _04572_);
  nor (_08591_, _08590_, _08589_);
  and (_08592_, _06175_, _04566_);
  and (_08593_, _06192_, _04550_);
  nor (_08594_, _08593_, _08592_);
  and (_08595_, _08594_, _08591_);
  and (_08596_, _08595_, _08588_);
  and (_08597_, _06179_, _04570_);
  and (_08598_, _06203_, _04557_);
  nor (_08599_, _08598_, _08597_);
  and (_08600_, _06170_, _04577_);
  and (_08601_, _06210_, _04544_);
  nor (_08602_, _08601_, _08600_);
  and (_08603_, _08602_, _08599_);
  and (_08604_, _06199_, _04546_);
  and (_08605_, _06166_, _04562_);
  nor (_08606_, _08605_, _08604_);
  and (_08607_, _06161_, _04540_);
  and (_08608_, _06182_, _04555_);
  nor (_08609_, _08608_, _08607_);
  and (_08610_, _08609_, _08606_);
  and (_08611_, _08610_, _08603_);
  and (_08612_, _08611_, _08596_);
  nor (_08613_, _08612_, _08581_);
  and (_08614_, _06832_, _06633_);
  and (_08615_, _06445_, _06215_);
  and (_08616_, _08615_, _08614_);
  and (_08617_, _06170_, _04623_);
  and (_08618_, _06203_, _04603_);
  nor (_08619_, _08618_, _08617_);
  and (_08620_, _06161_, _04585_);
  and (_08621_, _06166_, _04608_);
  nor (_08622_, _08621_, _08620_);
  and (_08623_, _08622_, _08619_);
  and (_08624_, _06197_, _04606_);
  and (_08625_, _06199_, _04592_);
  nor (_08626_, _08625_, _08624_);
  and (_08627_, _06185_, _04625_);
  and (_08628_, _06210_, _04587_);
  nor (_08629_, _08628_, _08627_);
  and (_08630_, _08629_, _08626_);
  and (_08631_, _08630_, _08623_);
  and (_08632_, _06192_, _04596_);
  and (_08633_, _06205_, _04614_);
  nor (_08634_, _08633_, _08632_);
  and (_08635_, _06187_, _04598_);
  and (_08636_, _06194_, _04618_);
  nor (_08637_, _08636_, _08635_);
  and (_08638_, _08637_, _08634_);
  and (_08639_, _06182_, _04601_);
  and (_08640_, _06179_, _04616_);
  nor (_08641_, _08640_, _08639_);
  and (_08642_, _06208_, _04590_);
  and (_08643_, _06175_, _04612_);
  nor (_08644_, _08643_, _08642_);
  and (_08645_, _08644_, _08641_);
  and (_08646_, _08645_, _08638_);
  and (_08647_, _08646_, _08631_);
  nor (_08648_, _08647_, _08332_);
  and (_08649_, _08648_, _08616_);
  and (_08650_, _08649_, _08613_);
  and (_08651_, _08650_, \oc8051_golden_model_1.B [7]);
  not (_08652_, _08612_);
  and (_08653_, _08652_, _08581_);
  and (_08654_, _08653_, _08649_);
  and (_08655_, _08654_, \oc8051_golden_model_1.ACC [7]);
  or (_08656_, _08655_, _08651_);
  and (_08657_, _08647_, _08549_);
  and (_08658_, _08612_, _08581_);
  and (_08659_, _08658_, _08657_);
  and (_08660_, _08659_, _08616_);
  and (_08661_, _08660_, \oc8051_golden_model_1.P0 [7]);
  not (_08662_, _06215_);
  and (_08663_, _06445_, _08662_);
  and (_08664_, _08663_, _08614_);
  not (_08665_, _08581_);
  and (_08666_, _08612_, _08665_);
  and (_08667_, _08666_, _08657_);
  and (_08668_, _08667_, _08664_);
  and (_08669_, _08668_, \oc8051_golden_model_1.SCON [7]);
  or (_08670_, _08669_, _08661_);
  or (_08671_, _08670_, _08656_);
  not (_08672_, _06633_);
  and (_08673_, _06832_, _08672_);
  and (_08674_, _08673_, _08663_);
  and (_08675_, _08674_, _08659_);
  and (_08676_, _08675_, \oc8051_golden_model_1.TMOD [7]);
  and (_08677_, _08674_, _08667_);
  and (_08678_, _08677_, \oc8051_golden_model_1.SBUF [7]);
  or (_08679_, _08678_, _08676_);
  and (_08680_, _08664_, _08659_);
  and (_08681_, _08680_, \oc8051_golden_model_1.TCON [7]);
  and (_08682_, _08667_, _08616_);
  and (_08683_, _08682_, \oc8051_golden_model_1.P1 [7]);
  or (_08684_, _08683_, _08681_);
  or (_08685_, _08684_, _08679_);
  and (_08686_, _08657_, _08653_);
  and (_08687_, _08686_, _08616_);
  and (_08688_, _08687_, \oc8051_golden_model_1.P2 [7]);
  and (_08689_, _08657_, _08613_);
  and (_08690_, _08689_, _08664_);
  and (_08691_, _08690_, \oc8051_golden_model_1.IP [7]);
  or (_08692_, _08691_, _08688_);
  and (_08693_, _08686_, _08664_);
  and (_08694_, _08693_, \oc8051_golden_model_1.IE [7]);
  and (_08695_, _08689_, _08616_);
  and (_08696_, _08695_, \oc8051_golden_model_1.P3 [7]);
  or (_08697_, _08696_, _08694_);
  or (_08698_, _08697_, _08692_);
  not (_08699_, _06832_);
  and (_08700_, _08699_, _06633_);
  and (_08701_, _08700_, _08663_);
  and (_08702_, _08701_, _08659_);
  and (_08703_, _08702_, \oc8051_golden_model_1.TL0 [7]);
  and (_08704_, _08666_, _08649_);
  and (_08705_, _08704_, \oc8051_golden_model_1.PSW [7]);
  or (_08706_, _08705_, _08703_);
  or (_08707_, _08706_, _08698_);
  or (_08708_, _08707_, _08685_);
  or (_08709_, _08708_, _08671_);
  nor (_08710_, _06445_, _06215_);
  and (_08711_, _08710_, _08659_);
  and (_08712_, _08711_, _08614_);
  and (_08713_, _08712_, \oc8051_golden_model_1.TH0 [7]);
  nor (_08714_, _06832_, _06633_);
  and (_08715_, _08714_, _08659_);
  and (_08716_, _08715_, _08663_);
  and (_08717_, _08716_, \oc8051_golden_model_1.TL1 [7]);
  and (_08718_, _08659_, _08615_);
  and (_08719_, _08673_, _08718_);
  and (_08720_, _08719_, \oc8051_golden_model_1.SP [7]);
  or (_08721_, _08720_, _08717_);
  or (_08722_, _08721_, _08713_);
  and (_08723_, _08715_, _08615_);
  and (_08724_, _08723_, \oc8051_golden_model_1.DPH [7]);
  and (_08725_, _08711_, _08673_);
  and (_08726_, _08725_, \oc8051_golden_model_1.TH1 [7]);
  or (_08727_, _08726_, _08724_);
  and (_08728_, _08700_, _08718_);
  and (_08729_, _08728_, \oc8051_golden_model_1.DPL [7]);
  not (_08730_, _06445_);
  and (_08731_, _08730_, _06215_);
  and (_08732_, _08731_, _08715_);
  and (_08733_, _08732_, \oc8051_golden_model_1.PCON [7]);
  or (_08734_, _08733_, _08729_);
  or (_08735_, _08734_, _08727_);
  or (_08736_, _08735_, _08722_);
  or (_08737_, _08736_, _08709_);
  or (_08738_, _08737_, _08550_);
  and (_08739_, _08738_, _07010_);
  nor (_08740_, _07267_, _07254_);
  nor (_08741_, _07023_, _07252_);
  and (_08742_, _08741_, _08740_);
  not (_08743_, _08742_);
  or (_08744_, _08743_, _08739_);
  or (_08745_, _08744_, _08548_);
  or (_08746_, _08742_, _05952_);
  and (_08747_, _08746_, _08745_);
  or (_08748_, _08747_, _06021_);
  and (_08749_, _08748_, _08335_);
  or (_08750_, _08749_, _05724_);
  not (_08751_, _06112_);
  nor (_08752_, _08751_, _05952_);
  and (_08753_, _08524_, _05724_);
  nor (_08754_, _08753_, _08752_);
  and (_08755_, _08754_, _08750_);
  not (_08756_, _06284_);
  nor (_08757_, _08756_, _05952_);
  not (_08758_, _08333_);
  nand (_08759_, _08332_, _07787_);
  and (_08760_, _08759_, _08758_);
  and (_08761_, _08760_, _08752_);
  or (_08762_, _08761_, _08757_);
  or (_08763_, _08762_, _08755_);
  not (_08764_, _08301_);
  not (_08765_, _08757_);
  nor (_08766_, _07787_, _08393_);
  and (_08767_, _07787_, _08393_);
  nor (_08768_, _08767_, _08766_);
  or (_08769_, _08768_, _08765_);
  and (_08770_, _08769_, _08764_);
  and (_08771_, _08770_, _08763_);
  or (_08772_, _08771_, _08334_);
  and (_08773_, _08772_, _08300_);
  and (_08774_, _08766_, _07031_);
  or (_08775_, _08774_, _05736_);
  or (_08776_, _08775_, _08773_);
  not (_08777_, _06130_);
  nor (_08778_, _08777_, _05952_);
  and (_08779_, _08524_, _05736_);
  nor (_08780_, _08779_, _08778_);
  and (_08781_, _08780_, _08776_);
  not (_08782_, _06292_);
  nor (_08783_, _08782_, _05952_);
  and (_08784_, _08759_, _08778_);
  or (_08785_, _08784_, _08783_);
  or (_08786_, _08785_, _08781_);
  nand (_08787_, _08767_, _08783_);
  and (_08788_, _08787_, _05734_);
  and (_08789_, _08788_, _08786_);
  nand (_08790_, _08391_, _05732_);
  nand (_08791_, _08790_, _08286_);
  or (_08792_, _08791_, _08789_);
  and (_08793_, _08792_, _08299_);
  and (_08794_, _08297_, _07210_);
  or (_08795_, _08794_, _07051_);
  or (_08796_, _08795_, _08793_);
  not (_08797_, _07050_);
  nand (_08798_, _08484_, _08461_);
  or (_08799_, _08436_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_08800_, _08438_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_08801_, _08800_, _08429_);
  and (_08802_, _08801_, _08799_);
  or (_08803_, _08438_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_08804_, _08436_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_08805_, _08804_, _08443_);
  and (_08806_, _08805_, _08803_);
  nor (_08807_, _08806_, _08802_);
  nand (_08808_, _08807_, _08422_);
  or (_08809_, _08436_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_08810_, _08438_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_08811_, _08810_, _08429_);
  and (_08812_, _08811_, _08809_);
  or (_08813_, _08438_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_08814_, _08436_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_08815_, _08814_, _08443_);
  and (_08816_, _08815_, _08813_);
  nor (_08817_, _08816_, _08812_);
  nand (_08818_, _08817_, _08449_);
  nand (_08819_, _08818_, _08808_);
  nand (_08820_, _08819_, _08413_);
  or (_08821_, _08438_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_08822_, _08436_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_08823_, _08822_, _08821_);
  nand (_08824_, _08823_, _08429_);
  or (_08825_, _08438_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_08826_, _08436_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_08827_, _08826_, _08825_);
  nand (_08828_, _08827_, _08443_);
  nand (_08829_, _08828_, _08824_);
  nand (_08830_, _08829_, _08422_);
  or (_08831_, _08438_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_08832_, _08436_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand (_08833_, _08832_, _08831_);
  nand (_08834_, _08833_, _08429_);
  or (_08835_, _08438_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_08836_, _08436_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_08837_, _08836_, _08835_);
  nand (_08838_, _08837_, _08443_);
  nand (_08839_, _08838_, _08834_);
  nand (_08840_, _08839_, _08449_);
  nand (_08841_, _08840_, _08830_);
  nand (_08842_, _08841_, _08462_);
  nand (_08843_, _08842_, _08820_);
  or (_08844_, _08436_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_08845_, _08438_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_08846_, _08845_, _08429_);
  and (_08847_, _08846_, _08844_);
  or (_08848_, _08438_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_08849_, _08436_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_08850_, _08849_, _08443_);
  and (_08851_, _08850_, _08848_);
  nor (_08852_, _08851_, _08847_);
  nand (_08853_, _08852_, _08422_);
  or (_08854_, _08436_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_08855_, _08438_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_08856_, _08855_, _08429_);
  and (_08857_, _08856_, _08854_);
  or (_08858_, _08438_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_08859_, _08436_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_08860_, _08859_, _08443_);
  and (_08861_, _08860_, _08858_);
  nor (_08862_, _08861_, _08857_);
  nand (_08863_, _08862_, _08449_);
  nand (_08864_, _08863_, _08853_);
  nand (_08865_, _08864_, _08413_);
  or (_08866_, _08438_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_08867_, _08436_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_08868_, _08867_, _08866_);
  nand (_08869_, _08868_, _08429_);
  or (_08870_, _08438_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_08871_, _08436_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_08872_, _08871_, _08870_);
  nand (_08873_, _08872_, _08443_);
  nand (_08874_, _08873_, _08869_);
  nand (_08875_, _08874_, _08422_);
  or (_08876_, _08438_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_08877_, _08436_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand (_08878_, _08877_, _08876_);
  nand (_08879_, _08878_, _08429_);
  or (_08880_, _08438_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_08881_, _08436_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_08882_, _08881_, _08880_);
  nand (_08883_, _08882_, _08443_);
  nand (_08884_, _08883_, _08879_);
  nand (_08885_, _08884_, _08449_);
  nand (_08886_, _08885_, _08875_);
  nand (_08887_, _08886_, _08462_);
  nand (_08888_, _08887_, _08865_);
  or (_08889_, _08436_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_08890_, _08438_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_08891_, _08890_, _08429_);
  and (_08892_, _08891_, _08889_);
  or (_08893_, _08438_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_08894_, _08436_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_08895_, _08894_, _08443_);
  and (_08896_, _08895_, _08893_);
  nor (_08897_, _08896_, _08892_);
  nand (_08898_, _08897_, _08422_);
  or (_08899_, _08436_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_08900_, _08438_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_08901_, _08900_, _08429_);
  and (_08902_, _08901_, _08899_);
  or (_08904_, _08438_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_08905_, _08436_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_08906_, _08905_, _08443_);
  and (_08907_, _08906_, _08904_);
  nor (_08908_, _08907_, _08902_);
  nand (_08909_, _08908_, _08449_);
  nand (_08910_, _08909_, _08898_);
  nand (_08911_, _08910_, _08413_);
  or (_08912_, _08438_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_08913_, _08436_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_08915_, _08913_, _08912_);
  nand (_08916_, _08915_, _08429_);
  or (_08917_, _08438_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_08918_, _08436_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_08919_, _08918_, _08917_);
  nand (_08920_, _08919_, _08443_);
  nand (_08921_, _08920_, _08916_);
  nand (_08922_, _08921_, _08422_);
  or (_08923_, _08438_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_08924_, _08436_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand (_08926_, _08924_, _08923_);
  nand (_08927_, _08926_, _08429_);
  or (_08928_, _08438_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_08929_, _08436_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_08930_, _08929_, _08928_);
  nand (_08931_, _08930_, _08443_);
  nand (_08932_, _08931_, _08927_);
  nand (_08933_, _08932_, _08449_);
  nand (_08934_, _08933_, _08922_);
  nand (_08935_, _08934_, _08462_);
  nand (_08937_, _08935_, _08911_);
  or (_08938_, _08436_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_08939_, _08438_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_08940_, _08939_, _08429_);
  and (_08941_, _08940_, _08938_);
  or (_08942_, _08438_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_08943_, _08436_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_08944_, _08943_, _08443_);
  and (_08945_, _08944_, _08942_);
  nor (_08946_, _08945_, _08941_);
  nand (_08948_, _08946_, _08422_);
  or (_08949_, _08436_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_08950_, _08438_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_08951_, _08950_, _08429_);
  and (_08952_, _08951_, _08949_);
  or (_08953_, _08438_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_08954_, _08436_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_08955_, _08954_, _08443_);
  and (_08956_, _08955_, _08953_);
  nor (_08957_, _08956_, _08952_);
  nand (_08959_, _08957_, _08449_);
  nand (_08960_, _08959_, _08948_);
  nand (_08961_, _08960_, _08413_);
  or (_08962_, _08438_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_08963_, _08436_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_08964_, _08963_, _08962_);
  nand (_08965_, _08964_, _08429_);
  or (_08966_, _08438_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_08967_, _08436_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_08968_, _08967_, _08966_);
  nand (_08970_, _08968_, _08443_);
  nand (_08971_, _08970_, _08965_);
  nand (_08972_, _08971_, _08422_);
  or (_08973_, _08438_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_08974_, _08436_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_08975_, _08974_, _08973_);
  nand (_08976_, _08975_, _08429_);
  or (_08977_, _08438_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_08978_, _08436_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_08979_, _08978_, _08977_);
  nand (_08980_, _08979_, _08443_);
  nand (_08981_, _08980_, _08976_);
  nand (_08982_, _08981_, _08449_);
  nand (_08983_, _08982_, _08972_);
  nand (_08984_, _08983_, _08462_);
  nand (_08985_, _08984_, _08961_);
  or (_08986_, _08436_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_08987_, _08438_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_08988_, _08987_, _08429_);
  and (_08989_, _08988_, _08986_);
  or (_08990_, _08438_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_08991_, _08436_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_08992_, _08991_, _08443_);
  and (_08993_, _08992_, _08990_);
  nor (_08994_, _08993_, _08989_);
  nand (_08995_, _08994_, _08422_);
  or (_08996_, _08436_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_08997_, _08438_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_08998_, _08997_, _08429_);
  and (_08999_, _08998_, _08996_);
  or (_09000_, _08438_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_09001_, _08436_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_09002_, _09001_, _08443_);
  and (_09003_, _09002_, _09000_);
  nor (_09004_, _09003_, _08999_);
  nand (_09005_, _09004_, _08449_);
  nand (_09006_, _09005_, _08995_);
  nand (_09007_, _09006_, _08413_);
  or (_09008_, _08438_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_09009_, _08436_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_09010_, _09009_, _09008_);
  nand (_09011_, _09010_, _08429_);
  or (_09012_, _08438_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_09013_, _08436_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_09014_, _09013_, _09012_);
  nand (_09015_, _09014_, _08443_);
  nand (_09016_, _09015_, _09011_);
  nand (_09017_, _09016_, _08422_);
  or (_09018_, _08438_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_09019_, _08436_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_09020_, _09019_, _09018_);
  nand (_09021_, _09020_, _08429_);
  or (_09022_, _08438_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_09023_, _08436_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_09024_, _09023_, _09022_);
  nand (_09025_, _09024_, _08443_);
  nand (_09026_, _09025_, _09021_);
  nand (_09027_, _09026_, _08449_);
  nand (_09028_, _09027_, _09017_);
  nand (_09029_, _09028_, _08462_);
  nand (_09030_, _09029_, _09007_);
  or (_09031_, _08436_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_09032_, _08438_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_09033_, _09032_, _08429_);
  and (_09034_, _09033_, _09031_);
  or (_09035_, _08438_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_09036_, _08436_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_09037_, _09036_, _08443_);
  and (_09038_, _09037_, _09035_);
  nor (_09039_, _09038_, _09034_);
  nand (_09040_, _09039_, _08422_);
  or (_09041_, _08436_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_09042_, _08438_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_09043_, _09042_, _08429_);
  and (_09044_, _09043_, _09041_);
  or (_09045_, _08438_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_09046_, _08436_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_09047_, _09046_, _08443_);
  and (_09048_, _09047_, _09045_);
  nor (_09049_, _09048_, _09044_);
  nand (_09050_, _09049_, _08449_);
  nand (_09051_, _09050_, _09040_);
  nand (_09052_, _09051_, _08413_);
  or (_09053_, _08438_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_09054_, _08436_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_09055_, _09054_, _09053_);
  nand (_09056_, _09055_, _08429_);
  or (_09057_, _08438_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_09058_, _08436_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_09059_, _09058_, _09057_);
  nand (_09060_, _09059_, _08443_);
  nand (_09061_, _09060_, _09056_);
  nand (_09062_, _09061_, _08422_);
  or (_09063_, _08438_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_09064_, _08436_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_09065_, _09064_, _09063_);
  nand (_09066_, _09065_, _08429_);
  or (_09067_, _08438_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_09068_, _08436_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_09069_, _09068_, _09067_);
  nand (_09070_, _09069_, _08443_);
  nand (_09071_, _09070_, _09066_);
  nand (_09072_, _09071_, _08449_);
  nand (_09073_, _09072_, _09062_);
  nand (_09074_, _09073_, _08462_);
  and (_09075_, _09074_, _09052_);
  or (_09076_, _08436_, \oc8051_golden_model_1.IRAM[1] [0]);
  or (_09077_, _08438_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_09078_, _09077_, _08429_);
  and (_09079_, _09078_, _09076_);
  or (_09080_, _08438_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_09081_, _08436_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_09082_, _09081_, _08443_);
  and (_09083_, _09082_, _09080_);
  nor (_09084_, _09083_, _09079_);
  nand (_09085_, _09084_, _08422_);
  or (_09086_, _08436_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_09087_, _08438_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_09088_, _09087_, _08429_);
  and (_09089_, _09088_, _09086_);
  or (_09090_, _08438_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_09091_, _08436_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_09092_, _09091_, _08443_);
  and (_09093_, _09092_, _09090_);
  nor (_09094_, _09093_, _09089_);
  nand (_09095_, _09094_, _08449_);
  nand (_09096_, _09095_, _09085_);
  nand (_09097_, _09096_, _08413_);
  or (_09098_, _08438_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_09099_, _08436_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_09100_, _09099_, _09098_);
  nand (_09101_, _09100_, _08429_);
  or (_09102_, _08438_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_09103_, _08436_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_09104_, _09103_, _09102_);
  nand (_09105_, _09104_, _08443_);
  nand (_09106_, _09105_, _09101_);
  nand (_09107_, _09106_, _08422_);
  or (_09108_, _08438_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_09109_, _08436_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand (_09110_, _09109_, _09108_);
  nand (_09111_, _09110_, _08429_);
  or (_09112_, _08438_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_09113_, _08436_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_09114_, _09113_, _09112_);
  nand (_09115_, _09114_, _08443_);
  nand (_09116_, _09115_, _09111_);
  nand (_09117_, _09116_, _08449_);
  nand (_09118_, _09117_, _09107_);
  nand (_09119_, _09118_, _08462_);
  and (_09120_, _09119_, _09097_);
  nor (_09121_, _09120_, _09075_);
  and (_09122_, _09121_, _09030_);
  and (_09123_, _09122_, _08985_);
  and (_09124_, _09123_, _08937_);
  and (_09125_, _09124_, _08888_);
  and (_09126_, _09125_, _08843_);
  nor (_09127_, _09126_, _08798_);
  and (_09128_, _09126_, _08798_);
  or (_09129_, _09128_, _09127_);
  or (_09130_, _09129_, _07052_);
  and (_09131_, _09130_, _08797_);
  and (_09132_, _09131_, _08796_);
  and (_09133_, _08498_, _07050_);
  or (_09134_, _09133_, _06127_);
  or (_09135_, _09134_, _09132_);
  and (_09136_, _05350_, \oc8051_golden_model_1.PC [2]);
  and (_09137_, _09136_, \oc8051_golden_model_1.PC [3]);
  and (_09138_, _09137_, _08387_);
  and (_09139_, _09138_, \oc8051_golden_model_1.PC [7]);
  nor (_09140_, _09138_, \oc8051_golden_model_1.PC [7]);
  nor (_09141_, _09140_, _09139_);
  not (_09142_, _09141_);
  nand (_09143_, _09142_, _06127_);
  and (_09144_, _09143_, _09135_);
  or (_09145_, _09144_, _05752_);
  and (_09146_, _08524_, _05752_);
  nor (_09147_, _09146_, _07058_);
  and (_09148_, _09147_, _09145_);
  and (_09149_, _08374_, _07058_);
  and (_09150_, _07005_, _05750_);
  or (_09151_, _09150_, _09149_);
  or (_09152_, _09151_, _09148_);
  nor (_09153_, _09152_, _08281_);
  nor (_09154_, _07609_, _06464_);
  not (_09155_, _07223_);
  not (_09156_, _07883_);
  not (_09157_, _07977_);
  not (_09158_, _08270_);
  not (_09159_, _07353_);
  not (_09160_, _07530_);
  not (_09161_, _07132_);
  and (_09162_, _09161_, _06931_);
  and (_09163_, _09162_, _09160_);
  and (_09164_, _09163_, _09159_);
  and (_09165_, _09164_, _09158_);
  and (_09166_, _09165_, _09157_);
  and (_09167_, _09166_, _09156_);
  nor (_09168_, _09167_, _08288_);
  and (_09169_, _09167_, _08288_);
  nor (_09170_, _09169_, _09168_);
  and (_09171_, _09170_, _09155_);
  nor (_09172_, _09171_, _09154_);
  nor (_09173_, _09172_, _09153_);
  and (_09174_, _09170_, _07223_);
  nor (_09175_, _09174_, _07068_);
  not (_09176_, _09175_);
  nor (_09177_, _09176_, _09173_);
  and (_09178_, _08842_, _08820_);
  and (_09179_, _08887_, _08865_);
  and (_09180_, _08935_, _08911_);
  and (_09181_, _08984_, _08961_);
  and (_09182_, _09029_, _09007_);
  and (_09183_, _09120_, _09075_);
  and (_09184_, _09183_, _09182_);
  and (_09185_, _09184_, _09181_);
  and (_09186_, _09185_, _09180_);
  and (_09187_, _09186_, _09179_);
  and (_09188_, _09187_, _09178_);
  nor (_09189_, _09188_, _08798_);
  and (_09190_, _09188_, _08798_);
  or (_09191_, _09190_, _09189_);
  nor (_09192_, _09191_, _07069_);
  nor (_09193_, _09192_, _07067_);
  not (_09194_, _09193_);
  nor (_09195_, _09194_, _09177_);
  nor (_09196_, _09195_, _08280_);
  nor (_09197_, _09196_, _07305_);
  or (_09198_, _09197_, _07634_);
  and (_09199_, _09198_, _07633_);
  not (_09200_, _06127_);
  and (_09201_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_09202_, _09201_, \oc8051_golden_model_1.PC [10]);
  and (_09203_, _09202_, _08389_);
  and (_09204_, _09203_, \oc8051_golden_model_1.PC [11]);
  and (_09205_, _09204_, \oc8051_golden_model_1.PC [12]);
  and (_09206_, _09205_, \oc8051_golden_model_1.PC [13]);
  and (_09207_, _09206_, \oc8051_golden_model_1.PC [14]);
  nor (_09208_, _09207_, \oc8051_golden_model_1.PC [15]);
  and (_09209_, _09201_, _08389_);
  and (_09210_, _09209_, \oc8051_golden_model_1.PC [10]);
  and (_09211_, _09210_, \oc8051_golden_model_1.PC [11]);
  and (_09212_, _09211_, \oc8051_golden_model_1.PC [12]);
  and (_09213_, _09212_, \oc8051_golden_model_1.PC [13]);
  and (_09214_, _09213_, \oc8051_golden_model_1.PC [14]);
  and (_09215_, _09214_, \oc8051_golden_model_1.PC [15]);
  nor (_09216_, _09215_, _09208_);
  and (_09217_, _09216_, _09200_);
  not (_09218_, \oc8051_golden_model_1.PC [15]);
  and (_09219_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and (_09220_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_09221_, _09220_, _09201_);
  and (_09222_, _09221_, _09139_);
  and (_09223_, _09222_, _09219_);
  and (_09224_, _09223_, \oc8051_golden_model_1.PC [14]);
  and (_09225_, _09224_, _09218_);
  nor (_09226_, _09224_, _09218_);
  or (_09227_, _09226_, _09225_);
  and (_09228_, _09227_, _06127_);
  or (_09229_, _09228_, _09217_);
  and (_09230_, _09229_, _07628_);
  and (_09231_, _09230_, _07631_);
  or (_40751_, _09231_, _09199_);
  not (_09232_, \oc8051_golden_model_1.B [7]);
  nor (_09233_, _01336_, _09232_);
  nor (_09234_, _07698_, _09232_);
  and (_09235_, _08768_, _07698_);
  or (_09236_, _09235_, _09234_);
  and (_09237_, _09236_, _06284_);
  nor (_09238_, _08361_, _09232_);
  and (_09239_, _08374_, _08361_);
  or (_09240_, _09239_, _09238_);
  and (_09241_, _09240_, _06039_);
  and (_09242_, _08498_, _07698_);
  or (_09243_, _09242_, _09234_);
  or (_09244_, _09243_, _06954_);
  and (_09245_, _07698_, \oc8051_golden_model_1.ACC [7]);
  or (_09246_, _09245_, _09234_);
  and (_09247_, _09246_, _06938_);
  nor (_09248_, _06938_, _09232_);
  or (_09249_, _09248_, _06102_);
  or (_09250_, _09249_, _09247_);
  and (_09251_, _09250_, _06044_);
  and (_09252_, _09251_, _09244_);
  and (_09253_, _08503_, _08361_);
  or (_09254_, _09253_, _09238_);
  and (_09255_, _09254_, _06043_);
  or (_09256_, _09255_, _06239_);
  or (_09257_, _09256_, _09252_);
  not (_09258_, _07698_);
  nor (_09259_, _07785_, _09258_);
  or (_09260_, _09259_, _09234_);
  or (_09261_, _09260_, _06848_);
  and (_09262_, _09261_, _09257_);
  or (_09263_, _09262_, _06219_);
  or (_09264_, _09246_, _06220_);
  and (_09265_, _09264_, _06040_);
  and (_09266_, _09265_, _09263_);
  or (_09267_, _09266_, _09241_);
  and (_09268_, _09267_, _06033_);
  and (_09269_, _06114_, _06221_);
  or (_09270_, _09238_, _08519_);
  and (_09271_, _09254_, _06032_);
  and (_09272_, _09271_, _09270_);
  or (_09273_, _09272_, _09269_);
  or (_09274_, _09273_, _09268_);
  and (_09275_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_09276_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_09277_, _09276_, _09275_);
  and (_09278_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [2]);
  and (_09279_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and (_09280_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor (_09281_, _09280_, _09279_);
  nor (_09282_, _09281_, _09277_);
  and (_09283_, _09282_, _09278_);
  nor (_09284_, _09283_, _09277_);
  and (_09285_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_09286_, _09285_, _09280_);
  and (_09287_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_09288_, _09287_, _09275_);
  nor (_09289_, _09288_, _09286_);
  not (_09290_, _09289_);
  nor (_09291_, _09290_, _09284_);
  and (_09292_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_09293_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [3]);
  and (_09294_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [4]);
  and (_09295_, _09294_, _09293_);
  nor (_09296_, _09294_, _09293_);
  nor (_09297_, _09296_, _09295_);
  and (_09298_, _09297_, _09292_);
  nor (_09299_, _09297_, _09292_);
  nor (_09300_, _09299_, _09298_);
  and (_09301_, _09290_, _09284_);
  nor (_09302_, _09301_, _09291_);
  and (_09303_, _09302_, _09300_);
  nor (_09304_, _09303_, _09291_);
  not (_09305_, _09280_);
  and (_09306_, _09285_, _09305_);
  and (_09307_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [5]);
  and (_09308_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_09309_, _09308_, _09293_);
  and (_09310_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [4]);
  and (_09311_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_09312_, _09311_, _09310_);
  nor (_09313_, _09312_, _09309_);
  and (_09314_, _09313_, _09307_);
  nor (_09315_, _09313_, _09307_);
  nor (_09316_, _09315_, _09314_);
  and (_09317_, _09316_, _09306_);
  nor (_09318_, _09316_, _09306_);
  nor (_09319_, _09318_, _09317_);
  not (_09320_, _09319_);
  nor (_09321_, _09320_, _09304_);
  and (_09322_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_09323_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [7]);
  and (_09324_, _09323_, _09322_);
  nor (_09325_, _09298_, _09295_);
  and (_09326_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.B [7]);
  and (_09327_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_09328_, _09327_, _09326_);
  nor (_09329_, _09327_, _09326_);
  nor (_09330_, _09329_, _09328_);
  not (_09331_, _09330_);
  nor (_09332_, _09331_, _09325_);
  and (_09333_, _09331_, _09325_);
  nor (_09334_, _09333_, _09332_);
  and (_09335_, _09334_, _09324_);
  nor (_09336_, _09334_, _09324_);
  nor (_09337_, _09336_, _09335_);
  and (_09338_, _09320_, _09304_);
  nor (_09339_, _09338_, _09321_);
  and (_09340_, _09339_, _09337_);
  nor (_09341_, _09340_, _09321_);
  nor (_09342_, _09314_, _09309_);
  and (_09343_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.B [7]);
  and (_09344_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [6]);
  and (_09345_, _09344_, _09343_);
  nor (_09346_, _09344_, _09343_);
  nor (_09347_, _09346_, _09345_);
  not (_09348_, _09347_);
  nor (_09349_, _09348_, _09342_);
  and (_09350_, _09348_, _09342_);
  nor (_09351_, _09350_, _09349_);
  and (_09352_, _09351_, _09328_);
  nor (_09353_, _09351_, _09328_);
  nor (_09354_, _09353_, _09352_);
  nor (_09355_, _09317_, _09286_);
  and (_09356_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [5]);
  and (_09357_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_09358_, _09357_, _09308_);
  nor (_09359_, _09357_, _09308_);
  nor (_09360_, _09359_, _09358_);
  and (_09361_, _09360_, _09356_);
  nor (_09362_, _09360_, _09356_);
  nor (_09363_, _09362_, _09361_);
  not (_09364_, _09363_);
  nor (_09365_, _09364_, _09355_);
  and (_09366_, _09364_, _09355_);
  nor (_09367_, _09366_, _09365_);
  and (_09368_, _09367_, _09354_);
  nor (_09369_, _09367_, _09354_);
  nor (_09370_, _09369_, _09368_);
  not (_09371_, _09370_);
  nor (_09372_, _09371_, _09341_);
  nor (_09373_, _09335_, _09332_);
  not (_09374_, _09373_);
  and (_09375_, _09371_, _09341_);
  nor (_09376_, _09375_, _09372_);
  and (_09377_, _09376_, _09374_);
  nor (_09378_, _09377_, _09372_);
  nor (_09379_, _09352_, _09349_);
  not (_09380_, _09379_);
  nor (_09381_, _09368_, _09365_);
  not (_09382_, _09381_);
  and (_09383_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_09384_, _09383_, _09308_);
  and (_09385_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_09386_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_09387_, _09386_, _09385_);
  nor (_09388_, _09387_, _09384_);
  nor (_09389_, _09361_, _09358_);
  and (_09390_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [7]);
  and (_09391_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [6]);
  and (_09392_, _09391_, _09390_);
  nor (_09393_, _09391_, _09390_);
  nor (_09394_, _09393_, _09392_);
  not (_09395_, _09394_);
  nor (_09396_, _09395_, _09389_);
  and (_09397_, _09395_, _09389_);
  nor (_09398_, _09397_, _09396_);
  and (_09399_, _09398_, _09345_);
  nor (_09400_, _09398_, _09345_);
  nor (_09401_, _09400_, _09399_);
  and (_09402_, _09401_, _09388_);
  nor (_09403_, _09401_, _09388_);
  nor (_09404_, _09403_, _09402_);
  and (_09405_, _09404_, _09382_);
  nor (_09406_, _09404_, _09382_);
  nor (_09407_, _09406_, _09405_);
  and (_09408_, _09407_, _09380_);
  nor (_09409_, _09407_, _09380_);
  nor (_09410_, _09409_, _09408_);
  not (_09411_, _09410_);
  nor (_09412_, _09411_, _09378_);
  nor (_09413_, _09408_, _09405_);
  nor (_09414_, _09399_, _09396_);
  not (_09415_, _09414_);
  and (_09416_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [7]);
  and (_09417_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_09418_, _09417_, _09416_);
  nor (_09419_, _09417_, _09416_);
  nor (_09420_, _09419_, _09418_);
  and (_09421_, _09420_, _09384_);
  nor (_09422_, _09420_, _09384_);
  nor (_09423_, _09422_, _09421_);
  and (_09424_, _09423_, _09392_);
  nor (_09425_, _09423_, _09392_);
  nor (_09426_, _09425_, _09424_);
  and (_09427_, _09426_, _09383_);
  nor (_09428_, _09426_, _09383_);
  nor (_09429_, _09428_, _09427_);
  and (_09430_, _09429_, _09402_);
  nor (_09431_, _09429_, _09402_);
  nor (_09432_, _09431_, _09430_);
  and (_09433_, _09432_, _09415_);
  nor (_09434_, _09432_, _09415_);
  nor (_09435_, _09434_, _09433_);
  not (_09436_, _09435_);
  nor (_09437_, _09436_, _09413_);
  and (_09438_, _09436_, _09413_);
  nor (_09439_, _09438_, _09437_);
  and (_09440_, _09439_, _09412_);
  nor (_09441_, _09433_, _09430_);
  nor (_09442_, _09424_, _09421_);
  not (_09443_, _09442_);
  and (_09444_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.B [7]);
  and (_09445_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_09446_, _09445_, _09444_);
  nor (_09447_, _09445_, _09444_);
  nor (_09448_, _09447_, _09446_);
  and (_09449_, _09448_, _09418_);
  nor (_09450_, _09448_, _09418_);
  nor (_09451_, _09450_, _09449_);
  and (_09452_, _09451_, _09427_);
  nor (_09453_, _09451_, _09427_);
  nor (_09454_, _09453_, _09452_);
  and (_09455_, _09454_, _09443_);
  nor (_09456_, _09454_, _09443_);
  nor (_09457_, _09456_, _09455_);
  not (_09458_, _09457_);
  nor (_09459_, _09458_, _09441_);
  and (_09460_, _09458_, _09441_);
  nor (_09461_, _09460_, _09459_);
  and (_09462_, _09461_, _09437_);
  nor (_09463_, _09461_, _09437_);
  nor (_09464_, _09463_, _09462_);
  and (_09465_, _09464_, _09440_);
  nor (_09466_, _09464_, _09440_);
  and (_09467_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  and (_09468_, _09467_, _09280_);
  and (_09469_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [2]);
  and (_09470_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [1]);
  nor (_09471_, _09470_, _09276_);
  nor (_09472_, _09471_, _09468_);
  and (_09473_, _09472_, _09469_);
  nor (_09474_, _09473_, _09468_);
  not (_09475_, _09474_);
  nor (_09476_, _09282_, _09278_);
  nor (_09477_, _09476_, _09283_);
  and (_09478_, _09477_, _09475_);
  and (_09479_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_09480_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [3]);
  and (_09481_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_09482_, _09481_, _09480_);
  nor (_09483_, _09481_, _09480_);
  nor (_09484_, _09483_, _09482_);
  and (_09485_, _09484_, _09479_);
  nor (_09486_, _09484_, _09479_);
  nor (_09487_, _09486_, _09485_);
  nor (_09488_, _09477_, _09475_);
  nor (_09489_, _09488_, _09478_);
  and (_09490_, _09489_, _09487_);
  nor (_09491_, _09490_, _09478_);
  nor (_09492_, _09302_, _09300_);
  nor (_09493_, _09492_, _09303_);
  not (_09494_, _09493_);
  nor (_09495_, _09494_, _09491_);
  and (_09496_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_09497_, _09496_, _09323_);
  nor (_09498_, _09485_, _09482_);
  nor (_09499_, _09323_, _09322_);
  nor (_09500_, _09499_, _09324_);
  not (_09501_, _09500_);
  nor (_09502_, _09501_, _09498_);
  and (_09503_, _09501_, _09498_);
  nor (_09504_, _09503_, _09502_);
  and (_09505_, _09504_, _09497_);
  nor (_09506_, _09504_, _09497_);
  nor (_09507_, _09506_, _09505_);
  and (_09508_, _09494_, _09491_);
  nor (_09509_, _09508_, _09495_);
  and (_09510_, _09509_, _09507_);
  nor (_09511_, _09510_, _09495_);
  nor (_09512_, _09339_, _09337_);
  nor (_09513_, _09512_, _09340_);
  not (_09514_, _09513_);
  nor (_09515_, _09514_, _09511_);
  nor (_09516_, _09505_, _09502_);
  not (_09517_, _09516_);
  and (_09518_, _09514_, _09511_);
  nor (_09520_, _09518_, _09515_);
  and (_09521_, _09520_, _09517_);
  nor (_09522_, _09521_, _09515_);
  nor (_09523_, _09376_, _09374_);
  nor (_09524_, _09523_, _09377_);
  not (_09525_, _09524_);
  nor (_09526_, _09525_, _09522_);
  and (_09527_, _09411_, _09378_);
  nor (_09528_, _09527_, _09412_);
  and (_09529_, _09528_, _09526_);
  nor (_09530_, _09439_, _09412_);
  nor (_09531_, _09530_, _09440_);
  nand (_09532_, _09531_, _09529_);
  and (_09533_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [1]);
  and (_09534_, _09533_, _09467_);
  and (_09535_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_09536_, _09533_, _09467_);
  nor (_09537_, _09536_, _09534_);
  and (_09538_, _09537_, _09535_);
  nor (_09539_, _09538_, _09534_);
  not (_09541_, _09539_);
  nor (_09542_, _09472_, _09469_);
  nor (_09543_, _09542_, _09473_);
  and (_09544_, _09543_, _09541_);
  and (_09545_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [5]);
  and (_09546_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_09547_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_09548_, _09547_, _09546_);
  nor (_09549_, _09547_, _09546_);
  nor (_09550_, _09549_, _09548_);
  and (_09551_, _09550_, _09545_);
  nor (_09552_, _09550_, _09545_);
  nor (_09553_, _09552_, _09551_);
  nor (_09554_, _09543_, _09541_);
  nor (_09555_, _09554_, _09544_);
  and (_09556_, _09555_, _09553_);
  nor (_09557_, _09556_, _09544_);
  not (_09558_, _09557_);
  nor (_09559_, _09489_, _09487_);
  nor (_09560_, _09559_, _09490_);
  and (_09561_, _09560_, _09558_);
  nor (_09562_, _09551_, _09548_);
  and (_09563_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [6]);
  and (_09564_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.B [7]);
  nor (_09565_, _09564_, _09563_);
  nor (_09566_, _09565_, _09497_);
  not (_09567_, _09566_);
  nor (_09568_, _09567_, _09562_);
  and (_09569_, _09567_, _09562_);
  nor (_09570_, _09569_, _09568_);
  nor (_09571_, _09560_, _09558_);
  nor (_09572_, _09571_, _09561_);
  and (_09573_, _09572_, _09570_);
  nor (_09574_, _09573_, _09561_);
  nor (_09575_, _09509_, _09507_);
  nor (_09576_, _09575_, _09510_);
  not (_09577_, _09576_);
  nor (_09578_, _09577_, _09574_);
  and (_09579_, _09577_, _09574_);
  nor (_09580_, _09579_, _09578_);
  and (_09581_, _09580_, _09568_);
  nor (_09582_, _09581_, _09578_);
  nor (_09583_, _09520_, _09517_);
  nor (_09584_, _09583_, _09521_);
  not (_09585_, _09584_);
  nor (_09586_, _09585_, _09582_);
  and (_09587_, _09525_, _09522_);
  nor (_09588_, _09587_, _09526_);
  and (_09589_, _09588_, _09586_);
  nor (_09590_, _09528_, _09526_);
  nor (_09591_, _09590_, _09529_);
  and (_09592_, _09591_, _09589_);
  nor (_09593_, _09591_, _09589_);
  nor (_09594_, _09593_, _09592_);
  and (_09595_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [0]);
  and (_09596_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_09597_, _09596_, _09595_);
  and (_09598_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_09599_, _09596_, _09595_);
  nor (_09600_, _09599_, _09597_);
  and (_09601_, _09600_, _09598_);
  nor (_09602_, _09601_, _09597_);
  not (_09603_, _09602_);
  nor (_09604_, _09537_, _09535_);
  nor (_09605_, _09604_, _09538_);
  and (_09606_, _09605_, _09603_);
  and (_09607_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_09608_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_09609_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [4]);
  and (_09610_, _09609_, _09608_);
  nor (_09611_, _09609_, _09608_);
  nor (_09612_, _09611_, _09610_);
  and (_09613_, _09612_, _09607_);
  nor (_09614_, _09612_, _09607_);
  nor (_09615_, _09614_, _09613_);
  nor (_09616_, _09605_, _09603_);
  nor (_09617_, _09616_, _09606_);
  and (_09618_, _09617_, _09615_);
  nor (_09619_, _09618_, _09606_);
  not (_09620_, _09619_);
  nor (_09621_, _09555_, _09553_);
  nor (_09622_, _09621_, _09556_);
  and (_09623_, _09622_, _09620_);
  not (_09624_, _09496_);
  nor (_09625_, _09613_, _09610_);
  nor (_09626_, _09625_, _09624_);
  and (_09627_, _09625_, _09624_);
  nor (_09628_, _09627_, _09626_);
  nor (_09629_, _09622_, _09620_);
  nor (_09630_, _09629_, _09623_);
  and (_09631_, _09630_, _09628_);
  nor (_09632_, _09631_, _09623_);
  not (_09633_, _09632_);
  nor (_09634_, _09572_, _09570_);
  nor (_09635_, _09634_, _09573_);
  and (_09636_, _09635_, _09633_);
  nor (_09637_, _09635_, _09633_);
  nor (_09638_, _09637_, _09636_);
  and (_09639_, _09638_, _09626_);
  nor (_09640_, _09639_, _09636_);
  nor (_09641_, _09580_, _09568_);
  nor (_09642_, _09641_, _09581_);
  not (_09643_, _09642_);
  nor (_09644_, _09643_, _09640_);
  and (_09645_, _09585_, _09582_);
  nor (_09646_, _09645_, _09586_);
  and (_09647_, _09646_, _09644_);
  nor (_09648_, _09588_, _09586_);
  nor (_09649_, _09648_, _09589_);
  nand (_09650_, _09649_, _09647_);
  or (_09651_, _09649_, _09647_);
  and (_09652_, _09651_, _09650_);
  and (_09653_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_09654_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_09655_, _09654_, _09653_);
  and (_09656_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [2]);
  nor (_09657_, _09654_, _09653_);
  nor (_09658_, _09657_, _09655_);
  and (_09659_, _09658_, _09656_);
  nor (_09660_, _09659_, _09655_);
  not (_09661_, _09660_);
  nor (_09662_, _09600_, _09598_);
  nor (_09663_, _09662_, _09601_);
  and (_09664_, _09663_, _09661_);
  and (_09665_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_09666_, _09665_, _09609_);
  and (_09667_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [3]);
  and (_09668_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_09669_, _09668_, _09667_);
  nor (_09670_, _09669_, _09666_);
  nor (_09671_, _09663_, _09661_);
  nor (_09672_, _09671_, _09664_);
  and (_09673_, _09672_, _09670_);
  nor (_09674_, _09673_, _09664_);
  not (_09675_, _09674_);
  nor (_09676_, _09617_, _09615_);
  nor (_09677_, _09676_, _09618_);
  and (_09678_, _09677_, _09675_);
  nor (_09679_, _09677_, _09675_);
  nor (_09680_, _09679_, _09678_);
  and (_09681_, _09680_, _09666_);
  nor (_09682_, _09681_, _09678_);
  not (_09683_, _09682_);
  nor (_09684_, _09630_, _09628_);
  nor (_09685_, _09684_, _09631_);
  and (_09686_, _09685_, _09683_);
  nor (_09687_, _09638_, _09626_);
  nor (_09688_, _09687_, _09639_);
  and (_09689_, _09688_, _09686_);
  and (_09690_, _09643_, _09640_);
  nor (_09691_, _09690_, _09644_);
  and (_09692_, _09691_, _09689_);
  nor (_09693_, _09646_, _09644_);
  nor (_09694_, _09693_, _09647_);
  and (_09696_, _09694_, _09692_);
  nor (_09697_, _09694_, _09692_);
  nor (_09699_, _09697_, _09696_);
  and (_09700_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_09702_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [1]);
  and (_09703_, _09702_, _09700_);
  and (_09705_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_09706_, _09702_, _09700_);
  nor (_09708_, _09706_, _09703_);
  and (_09709_, _09708_, _09705_);
  nor (_09711_, _09709_, _09703_);
  not (_09712_, _09711_);
  nor (_09714_, _09658_, _09656_);
  nor (_09715_, _09714_, _09659_);
  and (_09717_, _09715_, _09712_);
  nor (_09718_, _09715_, _09712_);
  nor (_09720_, _09718_, _09717_);
  and (_09721_, _09720_, _09665_);
  nor (_09723_, _09721_, _09717_);
  not (_09724_, _09723_);
  nor (_09726_, _09672_, _09670_);
  nor (_09727_, _09726_, _09673_);
  and (_09729_, _09727_, _09724_);
  nor (_09730_, _09680_, _09666_);
  nor (_09732_, _09730_, _09681_);
  and (_09733_, _09732_, _09729_);
  nor (_09734_, _09685_, _09683_);
  nor (_09735_, _09734_, _09686_);
  and (_09736_, _09735_, _09733_);
  nor (_09737_, _09688_, _09686_);
  nor (_09738_, _09737_, _09689_);
  and (_09739_, _09738_, _09736_);
  nor (_09740_, _09691_, _09689_);
  nor (_09741_, _09740_, _09692_);
  and (_09742_, _09741_, _09739_);
  and (_09743_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  and (_09744_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  and (_09745_, _09744_, _09743_);
  nor (_09746_, _09708_, _09705_);
  nor (_09747_, _09746_, _09709_);
  and (_09748_, _09747_, _09745_);
  nor (_09749_, _09720_, _09665_);
  nor (_09750_, _09749_, _09721_);
  and (_09751_, _09750_, _09748_);
  nor (_09752_, _09727_, _09724_);
  nor (_09753_, _09752_, _09729_);
  and (_09754_, _09753_, _09751_);
  nor (_09755_, _09732_, _09729_);
  nor (_09756_, _09755_, _09733_);
  and (_09757_, _09756_, _09754_);
  nor (_09758_, _09735_, _09733_);
  nor (_09759_, _09758_, _09736_);
  and (_09760_, _09759_, _09757_);
  nor (_09761_, _09738_, _09736_);
  nor (_09762_, _09761_, _09739_);
  and (_09763_, _09762_, _09760_);
  nor (_09764_, _09741_, _09739_);
  nor (_09765_, _09764_, _09742_);
  and (_09766_, _09765_, _09763_);
  nor (_09767_, _09766_, _09742_);
  not (_09768_, _09767_);
  and (_09769_, _09768_, _09699_);
  or (_09770_, _09769_, _09696_);
  nand (_09771_, _09770_, _09652_);
  and (_09772_, _09771_, _09650_);
  not (_09773_, _09772_);
  and (_09774_, _09773_, _09594_);
  or (_09775_, _09774_, _09592_);
  or (_09776_, _09531_, _09529_);
  and (_09777_, _09776_, _09532_);
  nand (_09778_, _09777_, _09775_);
  and (_09779_, _09778_, _09532_);
  nor (_09780_, _09779_, _09466_);
  or (_09781_, _09780_, _09465_);
  and (_09782_, \oc8051_golden_model_1.ACC [7], \oc8051_golden_model_1.B [7]);
  not (_09783_, _09782_);
  nor (_09784_, _09783_, _09417_);
  nor (_09785_, _09784_, _09449_);
  nor (_09786_, _09455_, _09452_);
  nor (_09787_, _09786_, _09785_);
  and (_09788_, _09786_, _09785_);
  nor (_09789_, _09788_, _09787_);
  not (_09791_, _09789_);
  nor (_09793_, _09462_, _09459_);
  and (_09794_, _09793_, _09791_);
  nor (_09796_, _09793_, _09791_);
  nor (_09797_, _09796_, _09794_);
  and (_09799_, _09797_, _09781_);
  not (_09800_, _09269_);
  or (_09802_, _09787_, _09446_);
  or (_09803_, _09802_, _09796_);
  or (_09805_, _09803_, _09800_);
  or (_09806_, _09805_, _09799_);
  and (_09808_, _09806_, _06027_);
  and (_09809_, _09808_, _09274_);
  and (_09811_, _08376_, _08361_);
  or (_09812_, _09811_, _09238_);
  and (_09814_, _09812_, _06026_);
  and (_09815_, _05659_, _05567_);
  nor (_09817_, _09815_, _07011_);
  not (_09818_, _09817_);
  or (_09820_, _09818_, _09814_);
  or (_09821_, _09820_, _09809_);
  and (_09823_, _08485_, _07698_);
  or (_09824_, _09234_, _07012_);
  or (_09826_, _09824_, _09823_);
  not (_09827_, _09815_);
  or (_09828_, _09827_, _09260_);
  and (_09829_, _09828_, _05669_);
  and (_09830_, _09829_, _09826_);
  and (_09831_, _09830_, _09821_);
  and (_09832_, _06114_, _05659_);
  not (_09833_, _05669_);
  and (_09834_, _08738_, _07698_);
  or (_09835_, _09834_, _09234_);
  and (_09836_, _09835_, _09833_);
  or (_09837_, _09836_, _09832_);
  or (_09838_, _09837_, _09831_);
  not (_09839_, _09832_);
  nor (_09840_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_09841_, _09840_, _09279_);
  not (_09842_, \oc8051_golden_model_1.B [1]);
  nor (_09843_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor (_09844_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and (_09845_, _09844_, _09843_);
  and (_09846_, _09845_, _09842_);
  nor (_09847_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not (_09848_, _09847_);
  and (_09849_, \oc8051_golden_model_1.B [0], _08393_);
  nor (_09850_, _09849_, _09848_);
  and (_09851_, _09850_, _09846_);
  and (_09852_, _09851_, _09841_);
  or (_09853_, _09851_, _08393_);
  not (_09854_, \oc8051_golden_model_1.B [4]);
  not (_09855_, \oc8051_golden_model_1.B [5]);
  nor (_09856_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_09857_, _09856_, _09855_);
  and (_09858_, _09857_, _09854_);
  nor (_09859_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.B [2]);
  and (_09860_, _09859_, _09858_);
  not (_09861_, \oc8051_golden_model_1.ACC [6]);
  and (_09862_, \oc8051_golden_model_1.B [0], _09861_);
  nor (_09863_, _09862_, _08393_);
  nor (_09864_, _09863_, _09842_);
  not (_09865_, _09864_);
  and (_09866_, _09865_, _09860_);
  nor (_09867_, _09866_, _09853_);
  nor (_09868_, _09867_, _09852_);
  and (_09869_, _09866_, \oc8051_golden_model_1.B [0]);
  nor (_09870_, _09869_, _09861_);
  and (_09871_, _09870_, _09842_);
  nor (_09872_, _09870_, _09842_);
  nor (_09873_, _09872_, _09871_);
  nor (_09874_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  nor (_09875_, _09874_, _09467_);
  nor (_09876_, _09875_, \oc8051_golden_model_1.ACC [4]);
  not (_09877_, \oc8051_golden_model_1.B [0]);
  and (_09878_, \oc8051_golden_model_1.ACC [4], _09877_);
  nor (_09879_, _09878_, \oc8051_golden_model_1.ACC [5]);
  not (_09880_, \oc8051_golden_model_1.ACC [4]);
  and (_09881_, _09880_, \oc8051_golden_model_1.B [0]);
  nor (_09882_, _09881_, _09879_);
  nor (_09883_, _09882_, _09876_);
  not (_09884_, _09883_);
  and (_09885_, _09884_, _09873_);
  nor (_09886_, _09868_, \oc8051_golden_model_1.B [2]);
  nor (_09887_, _09886_, _09871_);
  not (_09888_, _09887_);
  nor (_09889_, _09888_, _09885_);
  not (_09890_, _09889_);
  and (_09891_, \oc8051_golden_model_1.B [2], _08393_);
  nor (_09892_, _09891_, \oc8051_golden_model_1.B [7]);
  and (_09893_, _09892_, _09845_);
  and (_09894_, _09893_, _09890_);
  nor (_09895_, _09894_, _09868_);
  nor (_09896_, _09895_, _09852_);
  nor (_09897_, _09884_, _09873_);
  nor (_09898_, _09897_, _09885_);
  and (_09899_, _09898_, _09894_);
  not (_09900_, _09870_);
  nor (_09901_, _09894_, _09900_);
  nor (_09902_, _09901_, _09899_);
  nor (_09903_, _09902_, \oc8051_golden_model_1.B [2]);
  and (_09904_, _09902_, \oc8051_golden_model_1.B [2]);
  nor (_09905_, _09904_, _09903_);
  not (_09906_, \oc8051_golden_model_1.ACC [5]);
  nor (_09907_, _09894_, _09906_);
  and (_09908_, _09894_, _09875_);
  or (_09909_, _09908_, _09907_);
  and (_09910_, _09909_, _09842_);
  nor (_09911_, _09909_, _09842_);
  nor (_09912_, _09911_, _09881_);
  nor (_09913_, _09912_, _09910_);
  not (_09914_, _09913_);
  and (_09915_, _09914_, _09905_);
  nor (_09916_, _09896_, \oc8051_golden_model_1.B [3]);
  nor (_09917_, _09916_, _09903_);
  not (_09918_, _09917_);
  nor (_09919_, _09918_, _09915_);
  not (_09920_, _09919_);
  and (_09921_, \oc8051_golden_model_1.B [3], _08393_);
  not (_09922_, _09921_);
  and (_09923_, _09922_, _09858_);
  and (_09924_, _09923_, _09920_);
  nor (_09925_, _09924_, _09896_);
  nor (_09926_, _09925_, _09852_);
  not (_09927_, \oc8051_golden_model_1.B [3]);
  nor (_09928_, _09924_, _09902_);
  nor (_09929_, _09914_, _09905_);
  nor (_09930_, _09929_, _09915_);
  and (_09931_, _09930_, _09924_);
  or (_09932_, _09931_, _09928_);
  and (_09933_, _09932_, _09927_);
  nor (_09934_, _09932_, _09927_);
  nor (_09935_, _09934_, _09933_);
  not (_09936_, _09935_);
  nor (_09937_, _09924_, _09909_);
  nor (_09938_, _09911_, _09910_);
  and (_09939_, _09938_, _09881_);
  nor (_09940_, _09938_, _09881_);
  nor (_09941_, _09940_, _09939_);
  and (_09942_, _09941_, _09924_);
  or (_09943_, _09942_, _09937_);
  nor (_09944_, _09943_, \oc8051_golden_model_1.B [2]);
  and (_09945_, _09943_, \oc8051_golden_model_1.B [2]);
  nor (_09946_, _09881_, _09878_);
  and (_09947_, _09924_, _09946_);
  nor (_09948_, _09924_, \oc8051_golden_model_1.ACC [4]);
  nor (_09949_, _09948_, _09947_);
  and (_09950_, _09949_, _09842_);
  nor (_09951_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_09952_, _09951_, _09653_);
  nor (_09953_, _09952_, \oc8051_golden_model_1.ACC [2]);
  and (_09954_, _09877_, \oc8051_golden_model_1.ACC [2]);
  nor (_09955_, _09954_, \oc8051_golden_model_1.ACC [3]);
  not (_09956_, \oc8051_golden_model_1.ACC [2]);
  and (_09957_, \oc8051_golden_model_1.B [0], _09956_);
  nor (_09958_, _09957_, _09955_);
  nor (_09959_, _09958_, _09953_);
  not (_09960_, _09959_);
  nor (_09961_, _09949_, _09842_);
  nor (_09962_, _09961_, _09950_);
  and (_09963_, _09962_, _09960_);
  nor (_09964_, _09963_, _09950_);
  nor (_09965_, _09964_, _09945_);
  nor (_09966_, _09965_, _09944_);
  nor (_09967_, _09966_, _09936_);
  nor (_09968_, _09926_, \oc8051_golden_model_1.B [4]);
  nor (_09969_, _09968_, _09933_);
  not (_09970_, _09969_);
  nor (_09971_, _09970_, _09967_);
  not (_09972_, _09857_);
  and (_09973_, \oc8051_golden_model_1.B [4], _08393_);
  nor (_09974_, _09973_, _09972_);
  not (_09975_, _09974_);
  nor (_09976_, _09975_, _09971_);
  nor (_09977_, _09976_, _09926_);
  nor (_09978_, _09977_, _09852_);
  and (_09979_, _09856_, \oc8051_golden_model_1.ACC [7]);
  nor (_09980_, _09979_, _09857_);
  nor (_09981_, _09978_, \oc8051_golden_model_1.B [5]);
  and (_09982_, _09966_, _09936_);
  nor (_09983_, _09982_, _09967_);
  not (_09984_, _09983_);
  and (_09985_, _09984_, _09976_);
  nor (_09986_, _09976_, _09932_);
  nor (_09987_, _09986_, _09985_);
  and (_09988_, _09987_, _09854_);
  nor (_09989_, _09987_, _09854_);
  nor (_09990_, _09989_, _09988_);
  not (_09991_, _09990_);
  nor (_09992_, _09976_, _09943_);
  nor (_09993_, _09945_, _09944_);
  and (_09994_, _09993_, _09964_);
  nor (_09995_, _09993_, _09964_);
  nor (_09996_, _09995_, _09994_);
  not (_09997_, _09996_);
  and (_09998_, _09997_, _09976_);
  nor (_09999_, _09998_, _09992_);
  nor (_10000_, _09999_, \oc8051_golden_model_1.B [3]);
  and (_10001_, _09999_, \oc8051_golden_model_1.B [3]);
  not (_10002_, \oc8051_golden_model_1.B [2]);
  nor (_10003_, _09962_, _09960_);
  nor (_10004_, _10003_, _09963_);
  not (_10005_, _10004_);
  and (_10006_, _10005_, _09976_);
  nor (_10007_, _09976_, _09949_);
  nor (_10008_, _10007_, _10006_);
  and (_10009_, _10008_, _10002_);
  not (_10010_, \oc8051_golden_model_1.ACC [3]);
  nor (_10011_, _09976_, _10010_);
  and (_10012_, _09976_, _09952_);
  or (_10013_, _10012_, _10011_);
  and (_10014_, _10013_, _09842_);
  nor (_10015_, _10013_, _09842_);
  nor (_10016_, _10015_, _09957_);
  nor (_10017_, _10016_, _10014_);
  nor (_10018_, _10008_, _10002_);
  nor (_10019_, _10018_, _10009_);
  not (_10020_, _10019_);
  nor (_10021_, _10020_, _10017_);
  nor (_10022_, _10021_, _10009_);
  nor (_10023_, _10022_, _10001_);
  nor (_10024_, _10023_, _10000_);
  nor (_10025_, _10024_, _09991_);
  or (_10026_, _10025_, _09988_);
  nor (_10027_, _10026_, _09981_);
  nor (_10028_, _10027_, _09980_);
  nor (_10029_, _10028_, _09978_);
  nor (_10030_, _10029_, _09852_);
  not (_10031_, _10028_);
  and (_10032_, _10024_, _09991_);
  nor (_10033_, _10032_, _10025_);
  nor (_10034_, _10033_, _10031_);
  nor (_10035_, _10028_, _09987_);
  nor (_10036_, _10035_, _10034_);
  and (_10037_, _10036_, _09855_);
  nor (_10038_, _10036_, _09855_);
  nor (_10039_, _10038_, _10037_);
  nor (_10040_, _10028_, _09999_);
  nor (_10041_, _10001_, _10000_);
  nor (_10042_, _10041_, _10022_);
  and (_10043_, _10041_, _10022_);
  or (_10044_, _10043_, _10042_);
  and (_10045_, _10044_, _10028_);
  or (_10046_, _10045_, _10040_);
  and (_10047_, _10046_, _09854_);
  nor (_10048_, _10046_, _09854_);
  and (_10049_, _10020_, _10017_);
  nor (_10050_, _10049_, _10021_);
  nor (_10051_, _10050_, _10031_);
  nor (_10052_, _10028_, _10008_);
  nor (_10053_, _10052_, _10051_);
  and (_10054_, _10053_, _09927_);
  nor (_10055_, _10015_, _10014_);
  nor (_10056_, _10055_, _09957_);
  and (_10057_, _10055_, _09957_);
  or (_10058_, _10057_, _10056_);
  nor (_10059_, _10058_, _10031_);
  nor (_10060_, _10028_, _10013_);
  nor (_10061_, _10060_, _10059_);
  and (_10062_, _10061_, _10002_);
  nor (_10063_, _10061_, _10002_);
  nor (_10064_, _10028_, \oc8051_golden_model_1.ACC [2]);
  nor (_10065_, _09957_, _09954_);
  and (_10066_, _10028_, _10065_);
  nor (_10067_, _10066_, _10064_);
  and (_10068_, _10067_, _09842_);
  and (_10069_, _05784_, \oc8051_golden_model_1.B [0]);
  not (_10070_, _10069_);
  nor (_10071_, _10067_, _09842_);
  nor (_10072_, _10071_, _10068_);
  and (_10073_, _10072_, _10070_);
  nor (_10074_, _10073_, _10068_);
  nor (_10075_, _10074_, _10063_);
  nor (_10076_, _10075_, _10062_);
  not (_10077_, _10076_);
  nor (_10078_, _10053_, _09927_);
  nor (_10079_, _10078_, _10054_);
  and (_10080_, _10079_, _10077_);
  nor (_10081_, _10080_, _10054_);
  nor (_10082_, _10081_, _10048_);
  nor (_10083_, _10082_, _10047_);
  not (_10084_, _10083_);
  and (_10085_, _10084_, _10039_);
  nor (_10086_, _10030_, \oc8051_golden_model_1.B [6]);
  or (_10087_, _10086_, _10037_);
  or (_10088_, _10087_, _10085_);
  not (_10089_, \oc8051_golden_model_1.B [6]);
  or (_10090_, _10089_, \oc8051_golden_model_1.ACC [7]);
  and (_10091_, _10090_, _09232_);
  and (_10092_, _10091_, _10088_);
  nor (_10093_, _10092_, _10030_);
  or (_10094_, _10093_, _09852_);
  nor (_10095_, _10094_, \oc8051_golden_model_1.B [7]);
  nor (_10096_, _10095_, _09782_);
  nor (_10097_, _10084_, _10039_);
  nor (_10098_, _10097_, _10085_);
  and (_10099_, _10098_, _10092_);
  not (_10100_, _10036_);
  nor (_10101_, _10092_, _10100_);
  nor (_10102_, _10101_, _10099_);
  and (_10103_, _10102_, \oc8051_golden_model_1.B [6]);
  not (_10104_, _10103_);
  nor (_10105_, _10104_, _10096_);
  nor (_10106_, _10063_, _10062_);
  or (_10107_, _10106_, _10074_);
  nand (_10108_, _10106_, _10074_);
  and (_10109_, _10108_, _10107_);
  and (_10110_, _10109_, _10092_);
  nor (_10111_, _10092_, _10061_);
  nor (_10112_, _10111_, _10110_);
  and (_10113_, _10112_, _09927_);
  nor (_10114_, _10112_, _09927_);
  nor (_10115_, _10114_, _10113_);
  nor (_10116_, _10072_, _10070_);
  nor (_10117_, _10116_, _10073_);
  and (_10118_, _10117_, _10092_);
  not (_10119_, _10067_);
  nor (_10120_, _10092_, _10119_);
  nor (_10121_, _10120_, _10118_);
  and (_10122_, _10121_, \oc8051_golden_model_1.B [2]);
  nor (_10123_, _10121_, \oc8051_golden_model_1.B [2]);
  nor (_10124_, _10123_, _10122_);
  and (_10125_, _10124_, _10115_);
  or (_10126_, _10092_, \oc8051_golden_model_1.ACC [1]);
  nor (_10127_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  or (_10128_, _10127_, _09743_);
  nand (_10129_, _10092_, _10128_);
  and (_10130_, _10129_, _10126_);
  and (_10131_, _10130_, _09842_);
  nor (_10132_, _10130_, _09842_);
  and (_10133_, _09877_, \oc8051_golden_model_1.ACC [0]);
  not (_10134_, _10133_);
  nor (_10135_, _10134_, _10132_);
  nor (_10136_, _10135_, _10131_);
  and (_10137_, _10136_, _10125_);
  not (_10138_, _10137_);
  and (_10139_, _10122_, _10115_);
  nor (_10140_, _10139_, _10114_);
  and (_10141_, _10140_, _10138_);
  nor (_10142_, _10079_, _10077_);
  nor (_10143_, _10142_, _10080_);
  and (_10144_, _10143_, _10092_);
  not (_10145_, _10053_);
  nor (_10146_, _10092_, _10145_);
  nor (_10147_, _10146_, _10144_);
  and (_10148_, _10147_, \oc8051_golden_model_1.B [4]);
  nor (_10149_, _10147_, \oc8051_golden_model_1.B [4]);
  nor (_10150_, _10149_, _10148_);
  nor (_10151_, _10048_, _10047_);
  or (_10152_, _10151_, _10081_);
  nand (_10153_, _10151_, _10081_);
  and (_10154_, _10153_, _10152_);
  and (_10155_, _10154_, _10092_);
  nor (_10156_, _10092_, _10046_);
  nor (_10157_, _10156_, _10155_);
  nor (_10158_, _10157_, _09855_);
  and (_10159_, _10157_, _09855_);
  nor (_10160_, _10159_, _10158_);
  and (_10161_, _10160_, _10150_);
  nor (_10162_, _10102_, \oc8051_golden_model_1.B [6]);
  nor (_10163_, _10162_, _10103_);
  not (_10164_, _10163_);
  nor (_10165_, _10164_, _10096_);
  and (_10166_, _10165_, _10161_);
  not (_10167_, _10166_);
  nor (_10168_, _10167_, _10141_);
  and (_10169_, _10030_, \oc8051_golden_model_1.B [7]);
  and (_10170_, _10160_, _10148_);
  nor (_10171_, _10170_, _10158_);
  not (_10172_, _10171_);
  and (_10173_, _10172_, _10165_);
  or (_10174_, _10173_, _10169_);
  or (_10175_, _10174_, _10168_);
  nor (_10176_, _10175_, _10105_);
  nor (_10177_, _10132_, _10131_);
  and (_10178_, \oc8051_golden_model_1.B [0], _05758_);
  not (_10179_, _10178_);
  and (_10180_, _10179_, _10177_);
  and (_10181_, _10180_, _10134_);
  and (_10182_, _10181_, _10125_);
  and (_10183_, _10182_, _10166_);
  nor (_10184_, _10183_, _10176_);
  and (_10185_, _10184_, _10094_);
  or (_10186_, _10185_, _09852_);
  or (_10187_, _10186_, _09839_);
  and (_10188_, _10187_, _06020_);
  and (_10189_, _10188_, _09838_);
  and (_10190_, _08549_, _07698_);
  or (_10191_, _10190_, _09234_);
  and (_10192_, _10191_, _06019_);
  or (_10193_, _10192_, _06112_);
  or (_10194_, _10193_, _10189_);
  and (_10195_, _08760_, _07698_);
  or (_10196_, _10195_, _09234_);
  or (_10197_, _10196_, _08751_);
  and (_10198_, _10197_, _08756_);
  and (_10199_, _10198_, _10194_);
  or (_10200_, _10199_, _09237_);
  and (_10201_, _10200_, _07032_);
  or (_10202_, _09234_, _07788_);
  and (_10203_, _10191_, _06108_);
  and (_10204_, _10203_, _10202_);
  or (_10205_, _10204_, _10201_);
  and (_10206_, _10205_, _06278_);
  and (_10207_, _09246_, _06277_);
  and (_10208_, _10207_, _10202_);
  or (_10209_, _10208_, _06130_);
  or (_10210_, _10209_, _10206_);
  and (_10211_, _08759_, _07698_);
  or (_10212_, _09234_, _08777_);
  or (_10213_, _10212_, _10211_);
  and (_10214_, _10213_, _08782_);
  and (_10215_, _10214_, _10210_);
  nor (_10216_, _08767_, _09258_);
  or (_10217_, _10216_, _09234_);
  and (_10218_, _10217_, _06292_);
  or (_10219_, _10218_, _06316_);
  or (_10220_, _10219_, _10215_);
  or (_10221_, _09243_, _06718_);
  and (_10222_, _10221_, _05653_);
  and (_10223_, _10222_, _10220_);
  and (_10224_, _09240_, _05652_);
  or (_10225_, _10224_, _06047_);
  or (_10226_, _10225_, _10223_);
  and (_10227_, _08279_, _07698_);
  or (_10228_, _09234_, _06048_);
  or (_10229_, _10228_, _10227_);
  and (_10230_, _10229_, _01336_);
  and (_10231_, _10230_, _10226_);
  or (_10232_, _10231_, _09233_);
  and (_40752_, _10232_, _42882_);
  nor (_10233_, _01336_, _08393_);
  and (_10234_, _06931_, \oc8051_golden_model_1.PSW [7]);
  and (_10235_, _10234_, _09161_);
  and (_10236_, _10235_, _09160_);
  and (_10237_, _10236_, _09159_);
  and (_10238_, _10237_, _09158_);
  and (_10239_, _10238_, _09157_);
  and (_10240_, _10239_, _09156_);
  and (_10241_, _10240_, _08288_);
  nor (_10242_, _10240_, _08288_);
  or (_10243_, _10242_, _10241_);
  and (_10244_, _10243_, \oc8051_golden_model_1.ACC [7]);
  nor (_10245_, _10243_, \oc8051_golden_model_1.ACC [7]);
  nor (_10246_, _10245_, _10244_);
  nor (_10247_, _10239_, _09156_);
  nor (_10248_, _10247_, _10240_);
  and (_10249_, _10248_, \oc8051_golden_model_1.ACC [6]);
  nor (_10250_, _10248_, _09861_);
  and (_10251_, _10248_, _09861_);
  nor (_10252_, _10251_, _10250_);
  not (_10253_, _10252_);
  nor (_10254_, _10238_, _09157_);
  nor (_10255_, _10254_, _10239_);
  and (_10256_, _10255_, \oc8051_golden_model_1.ACC [5]);
  nor (_10257_, _10255_, _09906_);
  and (_10258_, _10255_, _09906_);
  nor (_10259_, _10258_, _10257_);
  nor (_10260_, _10237_, _09158_);
  nor (_10261_, _10260_, _10238_);
  nand (_10262_, _10261_, \oc8051_golden_model_1.ACC [4]);
  nor (_10263_, _10261_, _09880_);
  and (_10264_, _10261_, _09880_);
  or (_10265_, _10264_, _10263_);
  nor (_10266_, _10236_, _09159_);
  nor (_10267_, _10266_, _10237_);
  and (_10268_, _10267_, \oc8051_golden_model_1.ACC [3]);
  nor (_10269_, _10267_, _10010_);
  and (_10270_, _10267_, _10010_);
  nor (_10271_, _10270_, _10269_);
  nor (_10272_, _10235_, _09160_);
  nor (_10273_, _10272_, _10236_);
  and (_10274_, _10273_, \oc8051_golden_model_1.ACC [2]);
  nor (_10275_, _10273_, _09956_);
  and (_10276_, _10273_, _09956_);
  nor (_10277_, _10276_, _10275_);
  nor (_10278_, _10234_, _09161_);
  nor (_10279_, _10278_, _10235_);
  and (_10280_, _10279_, \oc8051_golden_model_1.ACC [1]);
  and (_10281_, _10279_, _05784_);
  nor (_10282_, _10279_, _05784_);
  nor (_10283_, _10282_, _10281_);
  nor (_10284_, _06931_, \oc8051_golden_model_1.PSW [7]);
  nor (_10285_, _10284_, _10234_);
  and (_10286_, _10285_, \oc8051_golden_model_1.ACC [0]);
  not (_10287_, _10286_);
  nor (_10288_, _10287_, _10283_);
  nor (_10289_, _10288_, _10280_);
  nor (_10290_, _10289_, _10277_);
  nor (_10291_, _10290_, _10274_);
  nor (_10292_, _10291_, _10271_);
  or (_10293_, _10292_, _10268_);
  nand (_10294_, _10293_, _10265_);
  and (_10295_, _10294_, _10262_);
  nor (_10296_, _10295_, _10259_);
  or (_10297_, _10296_, _10256_);
  and (_10298_, _10297_, _10253_);
  nor (_10299_, _10298_, _10249_);
  nor (_10300_, _10299_, _10246_);
  and (_10301_, _10299_, _10246_);
  nor (_10302_, _10301_, _10300_);
  and (_10303_, _05731_, _05567_);
  not (_10304_, _10303_);
  or (_10305_, _10304_, _10302_);
  and (_10306_, _06114_, _05671_);
  not (_10307_, _10306_);
  and (_10308_, _08127_, \oc8051_golden_model_1.PSW [7]);
  and (_10309_, _10308_, _08078_);
  and (_10310_, _10309_, _08177_);
  and (_10311_, _10310_, _08029_);
  and (_10312_, _10311_, _08273_);
  and (_10313_, _10312_, _07980_);
  and (_10314_, _10313_, _07886_);
  nor (_10315_, _10314_, _07787_);
  and (_10316_, _10314_, _07787_);
  nor (_10317_, _10316_, _10315_);
  and (_10318_, _10317_, \oc8051_golden_model_1.ACC [7]);
  nor (_10319_, _10317_, \oc8051_golden_model_1.ACC [7]);
  nor (_10320_, _10319_, _10318_);
  not (_10321_, _10320_);
  nor (_10322_, _10313_, _07886_);
  nor (_10323_, _10322_, _10314_);
  nor (_10324_, _10323_, _09861_);
  nor (_10325_, _10312_, _07980_);
  nor (_10326_, _10325_, _10313_);
  and (_10327_, _10326_, _09906_);
  nor (_10328_, _10326_, _09906_);
  nor (_10329_, _10328_, _10327_);
  not (_10330_, _10329_);
  nor (_10331_, _10311_, _08273_);
  nor (_10332_, _10331_, _10312_);
  nor (_10333_, _10332_, _09880_);
  and (_10334_, _10332_, _09880_);
  or (_10335_, _10334_, _10333_);
  or (_10336_, _10335_, _10330_);
  nor (_10337_, _10310_, _08029_);
  nor (_10338_, _10337_, _10311_);
  nor (_10339_, _10338_, _10010_);
  and (_10340_, _10338_, _10010_);
  nor (_10341_, _10340_, _10339_);
  nor (_10342_, _10309_, _08177_);
  nor (_10343_, _10342_, _10310_);
  nor (_10344_, _10343_, _09956_);
  and (_10345_, _10343_, _09956_);
  nor (_10346_, _10345_, _10344_);
  and (_10347_, _10346_, _10341_);
  nor (_10348_, _10308_, _08078_);
  nor (_10349_, _10348_, _10309_);
  nor (_10350_, _10349_, _05784_);
  and (_10351_, _10349_, _05784_);
  nor (_10352_, _08127_, \oc8051_golden_model_1.PSW [7]);
  nor (_10353_, _10352_, _10308_);
  and (_10354_, _10353_, _05758_);
  nor (_10355_, _10354_, _10351_);
  or (_10356_, _10355_, _10350_);
  nand (_10357_, _10356_, _10347_);
  and (_10358_, _10344_, _10341_);
  nor (_10359_, _10358_, _10339_);
  and (_10360_, _10359_, _10357_);
  nor (_10361_, _10360_, _10336_);
  and (_10362_, _10333_, _10329_);
  nor (_10363_, _10362_, _10328_);
  not (_10364_, _10363_);
  nor (_10365_, _10364_, _10361_);
  and (_10366_, _10323_, _09861_);
  nor (_10367_, _10324_, _10366_);
  not (_10368_, _10367_);
  nor (_10369_, _10368_, _10365_);
  or (_10370_, _10369_, _10324_);
  and (_10371_, _10370_, _10321_);
  nor (_10372_, _10370_, _10321_);
  or (_10373_, _10372_, _10371_);
  or (_10374_, _10373_, _06267_);
  and (_10375_, _10374_, _10307_);
  and (_10376_, _06114_, _06037_);
  nand (_10377_, _10376_, _10010_);
  nor (_10378_, _05693_, _08382_);
  nand (_10379_, _10378_, _07785_);
  nor (_10380_, _08359_, _08393_);
  and (_10381_, _08503_, _08359_);
  or (_10382_, _10381_, _10380_);
  or (_10383_, _10382_, _06044_);
  and (_10384_, _10383_, _06848_);
  nor (_10385_, _07701_, _08393_);
  and (_10386_, _08498_, _07701_);
  or (_10387_, _10386_, _10385_);
  and (_10388_, _10387_, _06102_);
  and (_10389_, _06114_, _06523_);
  not (_10390_, _10389_);
  or (_10391_, _10390_, _08485_);
  nor (_10392_, _06137_, _05697_);
  not (_10393_, _10392_);
  nor (_10394_, _05667_, _05661_);
  and (_10395_, _10394_, _06523_);
  nor (_10396_, _10395_, _06528_);
  and (_10397_, _06133_, _06523_);
  nor (_10398_, _10397_, _06525_);
  and (_10399_, _10398_, _10396_);
  and (_10400_, _10399_, _10393_);
  nor (_10401_, _10400_, _07785_);
  or (_10402_, _06530_, \oc8051_golden_model_1.ACC [7]);
  nand (_10403_, _06530_, \oc8051_golden_model_1.ACC [7]);
  and (_10404_, _10403_, _10402_);
  and (_10405_, _10404_, _10400_);
  or (_10406_, _10405_, _10389_);
  or (_10407_, _10406_, _10401_);
  and (_10408_, _06954_, _05698_);
  and (_10409_, _10408_, _10407_);
  and (_10410_, _10409_, _10391_);
  or (_10411_, _10410_, _10388_);
  and (_10412_, _06114_, _06042_);
  not (_10413_, _10412_);
  and (_10414_, _10413_, _10411_);
  nor (_10415_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [2]);
  nor (_10416_, _10415_, _10010_);
  and (_10417_, _10416_, \oc8051_golden_model_1.ACC [4]);
  and (_10418_, _10417_, \oc8051_golden_model_1.ACC [5]);
  and (_10419_, _10418_, \oc8051_golden_model_1.ACC [6]);
  and (_10420_, _10419_, \oc8051_golden_model_1.ACC [7]);
  nor (_10421_, _10419_, \oc8051_golden_model_1.ACC [7]);
  nor (_10422_, _10421_, _10420_);
  nor (_10423_, _10417_, \oc8051_golden_model_1.ACC [5]);
  nor (_10424_, _10423_, _10418_);
  nor (_10425_, _10418_, \oc8051_golden_model_1.ACC [6]);
  nor (_10426_, _10425_, _10419_);
  nor (_10427_, _10426_, _10424_);
  not (_10428_, _10427_);
  nand (_10429_, _10428_, _10422_);
  nor (_10430_, _10420_, \oc8051_golden_model_1.PSW [7]);
  and (_10431_, _10430_, _10429_);
  nor (_10432_, _10431_, _10427_);
  or (_10433_, _10432_, _10422_);
  and (_10434_, _10429_, _10412_);
  and (_10435_, _10434_, _10433_);
  or (_10436_, _10435_, _06043_);
  or (_10437_, _10436_, _10414_);
  and (_10438_, _10437_, _10384_);
  not (_10439_, _07701_);
  nor (_10440_, _07785_, _10439_);
  or (_10441_, _10440_, _10385_);
  and (_10442_, _10441_, _06239_);
  or (_10443_, _10442_, _10378_);
  or (_10444_, _10443_, _10438_);
  and (_10445_, _10444_, _10379_);
  or (_10446_, _10445_, _06970_);
  or (_10447_, _08485_, _06971_);
  and (_10448_, _10447_, _06220_);
  and (_10449_, _10448_, _10446_);
  nor (_10450_, _07787_, _06220_);
  or (_10451_, _10450_, _10376_);
  or (_10452_, _10451_, _10449_);
  and (_10453_, _10452_, _10377_);
  or (_10454_, _10453_, _06039_);
  and (_10455_, _08374_, _08359_);
  or (_10456_, _10455_, _10380_);
  or (_10457_, _10456_, _06040_);
  and (_10458_, _10457_, _06033_);
  and (_10459_, _10458_, _10454_);
  or (_10460_, _10380_, _08519_);
  and (_10461_, _10382_, _06032_);
  and (_10462_, _10461_, _10460_);
  or (_10463_, _10462_, _09269_);
  or (_10464_, _10463_, _10459_);
  nor (_10465_, _09762_, _09760_);
  nor (_10466_, _10465_, _09763_);
  or (_10467_, _10466_, _09800_);
  and (_10468_, _05671_, _05567_);
  not (_10469_, _10468_);
  and (_10470_, _10469_, _10467_);
  and (_10471_, _10470_, _10464_);
  nor (_10472_, _10263_, _10257_);
  nor (_10473_, _10472_, _10258_);
  not (_10474_, _10259_);
  or (_10475_, _10265_, _10474_);
  and (_10476_, _10277_, _10271_);
  and (_10477_, _10285_, _05758_);
  nor (_10478_, _10477_, _10281_);
  or (_10479_, _10478_, _10282_);
  nand (_10480_, _10479_, _10476_);
  and (_10481_, _10275_, _10271_);
  nor (_10482_, _10481_, _10269_);
  and (_10483_, _10482_, _10480_);
  nor (_10484_, _10483_, _10475_);
  nor (_10485_, _10484_, _10473_);
  nor (_10486_, _10485_, _10253_);
  or (_10487_, _10486_, _10250_);
  nor (_10488_, _10487_, _10246_);
  and (_10489_, _10487_, _10246_);
  or (_10490_, _10489_, _10488_);
  nor (_10491_, _10490_, _10469_);
  nor (_10492_, _10491_, _10471_);
  and (_10493_, _10394_, _05671_);
  nor (_10494_, _10493_, _10492_);
  and (_10495_, _09188_, \oc8051_golden_model_1.PSW [7]);
  nor (_10496_, _10495_, _08798_);
  and (_10497_, _10495_, _08798_);
  nor (_10498_, _10497_, _10496_);
  and (_10499_, _10498_, \oc8051_golden_model_1.ACC [7]);
  nor (_10500_, _10498_, \oc8051_golden_model_1.ACC [7]);
  nor (_10501_, _10500_, _10499_);
  not (_10502_, _10501_);
  and (_10503_, _09187_, \oc8051_golden_model_1.PSW [7]);
  nor (_10504_, _10503_, _09178_);
  nor (_10505_, _10504_, _10495_);
  nor (_10506_, _10505_, _09861_);
  and (_10507_, _09186_, \oc8051_golden_model_1.PSW [7]);
  nor (_10508_, _10507_, _09179_);
  nor (_10509_, _10508_, _10503_);
  and (_10510_, _10509_, _09906_);
  nor (_10511_, _10509_, _09906_);
  and (_10512_, _09185_, \oc8051_golden_model_1.PSW [7]);
  nor (_10513_, _10512_, _09180_);
  nor (_10514_, _10513_, _10507_);
  nor (_10515_, _10514_, _09880_);
  nor (_10516_, _10515_, _10511_);
  nor (_10517_, _10516_, _10510_);
  nor (_10518_, _10511_, _10510_);
  not (_10519_, _10518_);
  and (_10520_, _10514_, _09880_);
  or (_10521_, _10520_, _10515_);
  or (_10522_, _10521_, _10519_);
  and (_10523_, _09184_, \oc8051_golden_model_1.PSW [7]);
  nor (_10524_, _10523_, _09181_);
  nor (_10525_, _10524_, _10512_);
  nor (_10526_, _10525_, _10010_);
  and (_10527_, _10525_, _10010_);
  nor (_10528_, _10527_, _10526_);
  and (_10529_, _09183_, \oc8051_golden_model_1.PSW [7]);
  nor (_10530_, _10529_, _09182_);
  nor (_10531_, _10530_, _10523_);
  nor (_10532_, _10531_, _09956_);
  and (_10533_, _10531_, _09956_);
  nor (_10534_, _10533_, _10532_);
  and (_10535_, _10534_, _10528_);
  and (_10536_, _09120_, \oc8051_golden_model_1.PSW [7]);
  nor (_10537_, _10536_, _09075_);
  nor (_10538_, _10537_, _10529_);
  nor (_10539_, _10538_, _05784_);
  and (_10540_, _10538_, _05784_);
  nor (_10541_, _09120_, \oc8051_golden_model_1.PSW [7]);
  nor (_10542_, _10541_, _10536_);
  and (_10543_, _10542_, _05758_);
  nor (_10544_, _10543_, _10540_);
  or (_10545_, _10544_, _10539_);
  nand (_10546_, _10545_, _10535_);
  and (_10547_, _10532_, _10528_);
  nor (_10548_, _10547_, _10526_);
  and (_10549_, _10548_, _10546_);
  nor (_10550_, _10549_, _10522_);
  nor (_10551_, _10550_, _10517_);
  and (_10552_, _10505_, _09861_);
  nor (_10553_, _10506_, _10552_);
  not (_10554_, _10553_);
  nor (_10555_, _10554_, _10551_);
  or (_10556_, _10555_, _10506_);
  and (_10557_, _10556_, _10502_);
  nor (_10558_, _10556_, _10502_);
  or (_10559_, _10558_, _10557_);
  and (_10560_, _10559_, _10493_);
  nor (_10561_, _10560_, _10494_);
  nor (_10562_, _10561_, _06591_);
  and (_10563_, _10559_, _06591_);
  or (_10564_, _10563_, _10562_);
  or (_10565_, _10564_, _06261_);
  and (_10566_, _10565_, _10375_);
  and (_10567_, _08375_, _06299_);
  and (_10568_, _10567_, _07697_);
  and (_10569_, _10567_, _07690_);
  and (_10570_, _10569_, _07414_);
  nor (_10571_, _10570_, _05952_);
  nor (_10572_, _10571_, _10568_);
  nor (_10573_, _10572_, _08393_);
  and (_10574_, _10572_, _08393_);
  nor (_10575_, _10574_, _10573_);
  nor (_10576_, _10569_, _07414_);
  nor (_10577_, _10576_, _10570_);
  nor (_10578_, _10577_, _09861_);
  and (_10579_, _10567_, _07674_);
  nor (_10580_, _10579_, _07683_);
  nor (_10581_, _10580_, _10569_);
  and (_10582_, _10581_, _09906_);
  nor (_10583_, _10581_, _09906_);
  nor (_10584_, _10567_, _07674_);
  nor (_10585_, _10584_, _10579_);
  nor (_10586_, _10585_, _09880_);
  nor (_10587_, _10586_, _10583_);
  nor (_10588_, _10587_, _10582_);
  nor (_10589_, _10583_, _10582_);
  not (_10590_, _10589_);
  and (_10591_, _10585_, _09880_);
  or (_10592_, _10591_, _10586_);
  or (_10593_, _10592_, _10590_);
  nor (_10594_, _08375_, _06299_);
  nor (_10595_, _10594_, _10567_);
  nor (_10596_, _10595_, _10010_);
  and (_10597_, _10595_, _10010_);
  nor (_10598_, _10597_, _10596_);
  and (_10599_, _07639_, \oc8051_golden_model_1.PSW [7]);
  nor (_10600_, _10599_, _07477_);
  or (_10601_, _10600_, _08375_);
  and (_10602_, _10601_, \oc8051_golden_model_1.ACC [2]);
  nor (_10603_, _10601_, \oc8051_golden_model_1.ACC [2]);
  nor (_10604_, _10603_, _10602_);
  and (_10605_, _10604_, _10598_);
  not (_10606_, \oc8051_golden_model_1.PSW [7]);
  nor (_10607_, _06016_, _10606_);
  nor (_10608_, _10607_, _07076_);
  nor (_10609_, _10608_, _10599_);
  nor (_10610_, _10609_, _05784_);
  and (_10611_, _10609_, _05784_);
  nor (_10612_, _06016_, \oc8051_golden_model_1.PSW [7]);
  and (_10613_, _06016_, \oc8051_golden_model_1.PSW [7]);
  nor (_10614_, _10613_, _10612_);
  nor (_10615_, _10614_, \oc8051_golden_model_1.ACC [0]);
  nor (_10616_, _10615_, _10611_);
  or (_10617_, _10616_, _10610_);
  nand (_10618_, _10617_, _10605_);
  and (_10619_, _10602_, _10598_);
  nor (_10620_, _10619_, _10596_);
  and (_10621_, _10620_, _10618_);
  nor (_10622_, _10621_, _10593_);
  nor (_10623_, _10622_, _10588_);
  and (_10624_, _10577_, _09861_);
  nor (_10625_, _10578_, _10624_);
  not (_10626_, _10625_);
  nor (_10627_, _10626_, _10623_);
  or (_10628_, _10627_, _10578_);
  nor (_10629_, _10628_, _10575_);
  and (_10630_, _10628_, _10575_);
  or (_10631_, _10630_, _10629_);
  nor (_10632_, _10631_, _10307_);
  or (_10633_, _10632_, _05676_);
  or (_10634_, _10633_, _10566_);
  or (_10635_, _05952_, _05675_);
  and (_10636_, _10635_, _06027_);
  and (_10637_, _10636_, _10634_);
  and (_10638_, _08376_, _08359_);
  or (_10639_, _10638_, _10380_);
  and (_10640_, _10639_, _06026_);
  or (_10641_, _10640_, _09818_);
  or (_10642_, _10641_, _10637_);
  and (_10643_, _08485_, _07701_);
  or (_10644_, _10385_, _07012_);
  or (_10645_, _10644_, _10643_);
  or (_10646_, _10441_, _09827_);
  and (_10647_, _10646_, _05669_);
  and (_10648_, _10647_, _10645_);
  and (_10649_, _10648_, _10642_);
  and (_10650_, _08738_, _07701_);
  or (_10651_, _10650_, _10385_);
  and (_10652_, _10651_, _09833_);
  or (_10653_, _10652_, _09832_);
  or (_10654_, _10653_, _10649_);
  or (_10655_, _09851_, _09839_);
  and (_10656_, _10655_, _05664_);
  and (_10657_, _10656_, _10654_);
  and (_10658_, _05952_, _05663_);
  or (_10659_, _10658_, _06019_);
  or (_10660_, _10659_, _10657_);
  and (_10661_, _06114_, _05723_);
  not (_10662_, _10661_);
  and (_10663_, _08549_, _07701_);
  or (_10664_, _10663_, _10385_);
  or (_10665_, _10664_, _06020_);
  and (_10666_, _10665_, _10662_);
  and (_10667_, _10666_, _10660_);
  and (_10668_, _10661_, _05952_);
  and (_10669_, _07005_, _05726_);
  or (_10670_, _10669_, _10668_);
  or (_10671_, _10670_, _10667_);
  and (_10672_, _07785_, _08393_);
  nor (_10673_, _07785_, _08393_);
  nor (_10674_, _10673_, _10672_);
  not (_10675_, _10669_);
  or (_10676_, _10675_, _10674_);
  nor (_10677_, _06137_, _06644_);
  not (_10678_, _10677_);
  and (_10679_, _10678_, _10676_);
  and (_10680_, _10679_, _10671_);
  and (_10681_, _07002_, _05726_);
  and (_10682_, _10677_, _10674_);
  or (_10683_, _10682_, _10681_);
  or (_10684_, _10683_, _10680_);
  and (_10685_, _06103_, _05726_);
  not (_10686_, _10685_);
  not (_10687_, _10681_);
  or (_10688_, _10687_, _10674_);
  and (_10689_, _10688_, _10686_);
  and (_10690_, _10689_, _10684_);
  and (_10691_, _08798_, _08393_);
  and (_10692_, _08485_, \oc8051_golden_model_1.ACC [7]);
  nor (_10693_, _10692_, _10691_);
  and (_10694_, _10685_, _10693_);
  or (_10695_, _10694_, _06282_);
  or (_10697_, _10695_, _10690_);
  and (_10698_, _06114_, _05726_);
  not (_10699_, _10698_);
  or (_10700_, _08768_, _06283_);
  and (_10701_, _10700_, _10699_);
  and (_10702_, _10701_, _10697_);
  nor (_10703_, _05952_, \oc8051_golden_model_1.ACC [7]);
  and (_10704_, _05952_, \oc8051_golden_model_1.ACC [7]);
  nor (_10705_, _10704_, _10703_);
  and (_10706_, _10698_, _10705_);
  or (_10708_, _10706_, _06112_);
  or (_10709_, _10708_, _10702_);
  and (_10710_, _08760_, _07701_);
  or (_10711_, _10710_, _10385_);
  or (_10712_, _10711_, _08751_);
  and (_10713_, _10712_, _08756_);
  and (_10714_, _10713_, _10709_);
  and (_10715_, _10385_, _06284_);
  or (_10716_, _10715_, _06482_);
  or (_10717_, _10716_, _10714_);
  not (_10719_, _10673_);
  nand (_10720_, _10719_, _06482_);
  and (_10721_, _06096_, _05735_);
  not (_10722_, _10721_);
  not (_10723_, _06490_);
  and (_10724_, _06133_, _05735_);
  nor (_10725_, _10724_, _06835_);
  and (_10726_, _10725_, _10723_);
  and (_10727_, _10726_, _10722_);
  and (_10728_, _10727_, _10720_);
  and (_10730_, _10728_, _10717_);
  and (_10731_, _06103_, _05735_);
  nor (_10732_, _10727_, _10719_);
  or (_10733_, _10732_, _10731_);
  or (_10734_, _10733_, _10730_);
  not (_10735_, _06279_);
  not (_10736_, _10731_);
  or (_10737_, _10736_, _10692_);
  and (_10738_, _10737_, _10735_);
  and (_10739_, _10738_, _10734_);
  and (_10741_, _06114_, _05735_);
  nor (_10742_, _10741_, _06279_);
  not (_10743_, _10742_);
  or (_10744_, _10741_, _08766_);
  and (_10745_, _10744_, _10743_);
  or (_10746_, _10745_, _10739_);
  not (_10747_, _10741_);
  or (_10748_, _10747_, _10704_);
  and (_10749_, _10748_, _07032_);
  and (_10750_, _10749_, _10746_);
  and (_10752_, _06450_, _05739_);
  nand (_10753_, _10664_, _06108_);
  nor (_10754_, _10753_, _08767_);
  or (_10755_, _10754_, _10752_);
  or (_10756_, _10755_, _10750_);
  not (_10757_, _05739_);
  nor (_10758_, _06460_, _06229_);
  nor (_10759_, _10758_, _10757_);
  not (_10760_, _10759_);
  nand (_10761_, _10672_, _10752_);
  and (_10763_, _10761_, _10760_);
  and (_10764_, _10763_, _10756_);
  and (_10765_, _06133_, _05739_);
  nor (_10766_, _10765_, _06665_);
  not (_10767_, _10766_);
  nor (_10768_, _10760_, _10672_);
  or (_10769_, _10768_, _10767_);
  or (_10770_, _10769_, _10764_);
  nand (_10771_, _10767_, _10672_);
  and (_10772_, _10771_, _06668_);
  and (_10773_, _10772_, _10770_);
  nor (_10774_, _10672_, _06668_);
  and (_10775_, _06103_, _05739_);
  or (_10776_, _10775_, _10774_);
  or (_10777_, _10776_, _10773_);
  nand (_10778_, _10775_, _10691_);
  and (_10779_, _10778_, _06291_);
  and (_10780_, _10779_, _10777_);
  and (_10781_, _06114_, _05739_);
  nor (_10782_, _08767_, _06291_);
  or (_10783_, _10782_, _10781_);
  or (_10784_, _10783_, _10780_);
  nand (_10785_, _10781_, _10703_);
  and (_10786_, _10785_, _08777_);
  and (_10787_, _10786_, _10784_);
  and (_10788_, _08759_, _07701_);
  or (_10789_, _10788_, _10385_);
  and (_10790_, _10789_, _06130_);
  or (_10791_, _10790_, _10303_);
  or (_10792_, _10791_, _10787_);
  and (_10793_, _10792_, _10305_);
  and (_10794_, _06103_, _05731_);
  or (_10795_, _10794_, _10793_);
  not (_10796_, _10794_);
  nand (_10797_, _10505_, \oc8051_golden_model_1.ACC [6]);
  and (_10798_, _10509_, \oc8051_golden_model_1.ACC [5]);
  nand (_10799_, _10514_, \oc8051_golden_model_1.ACC [4]);
  and (_10800_, _10525_, \oc8051_golden_model_1.ACC [3]);
  and (_10801_, _10531_, \oc8051_golden_model_1.ACC [2]);
  and (_10802_, _10538_, \oc8051_golden_model_1.ACC [1]);
  nor (_10803_, _10540_, _10539_);
  and (_10804_, _10542_, \oc8051_golden_model_1.ACC [0]);
  not (_10805_, _10804_);
  nor (_10806_, _10805_, _10803_);
  nor (_10807_, _10806_, _10802_);
  nor (_10808_, _10807_, _10534_);
  nor (_10809_, _10808_, _10801_);
  nor (_10810_, _10809_, _10528_);
  or (_10811_, _10810_, _10800_);
  nand (_10812_, _10811_, _10521_);
  and (_10813_, _10812_, _10799_);
  nor (_10814_, _10813_, _10518_);
  or (_10815_, _10814_, _10798_);
  nand (_10816_, _10815_, _10554_);
  and (_10817_, _10816_, _10797_);
  nor (_10818_, _10817_, _10501_);
  and (_10819_, _10817_, _10501_);
  nor (_10820_, _10819_, _10818_);
  or (_10821_, _10820_, _10796_);
  and (_10822_, _10821_, _06289_);
  and (_10823_, _10822_, _10795_);
  and (_10824_, _06114_, _05731_);
  nor (_10825_, _10824_, _06288_);
  not (_10826_, _10825_);
  and (_10827_, _10323_, \oc8051_golden_model_1.ACC [6]);
  and (_10828_, _10326_, \oc8051_golden_model_1.ACC [5]);
  nand (_10829_, _10332_, \oc8051_golden_model_1.ACC [4]);
  and (_10830_, _10338_, \oc8051_golden_model_1.ACC [3]);
  and (_10831_, _10343_, \oc8051_golden_model_1.ACC [2]);
  and (_10832_, _10349_, \oc8051_golden_model_1.ACC [1]);
  nor (_10833_, _10351_, _10350_);
  not (_10834_, _10833_);
  and (_10835_, _10353_, \oc8051_golden_model_1.ACC [0]);
  and (_10836_, _10835_, _10834_);
  nor (_10837_, _10836_, _10832_);
  nor (_10838_, _10837_, _10346_);
  nor (_10839_, _10838_, _10831_);
  nor (_10840_, _10839_, _10341_);
  or (_10841_, _10840_, _10830_);
  nand (_10842_, _10841_, _10335_);
  and (_10843_, _10842_, _10829_);
  nor (_10844_, _10843_, _10329_);
  or (_10845_, _10844_, _10828_);
  and (_10846_, _10845_, _10368_);
  nor (_10847_, _10846_, _10827_);
  nor (_10848_, _10847_, _10320_);
  and (_10849_, _10847_, _10320_);
  nor (_10850_, _10849_, _10848_);
  or (_10851_, _10850_, _10824_);
  and (_10852_, _10851_, _10826_);
  or (_10853_, _10852_, _10823_);
  and (_10854_, _05731_, _06107_);
  not (_10855_, _10854_);
  not (_10856_, _10824_);
  nand (_10857_, _10577_, \oc8051_golden_model_1.ACC [6]);
  and (_10858_, _10581_, \oc8051_golden_model_1.ACC [5]);
  nand (_10859_, _10585_, \oc8051_golden_model_1.ACC [4]);
  and (_10860_, _10595_, \oc8051_golden_model_1.ACC [3]);
  nor (_10861_, _10601_, _09956_);
  and (_10862_, _10609_, \oc8051_golden_model_1.ACC [1]);
  nor (_10863_, _10611_, _10610_);
  not (_10864_, _10863_);
  nor (_10865_, _10614_, _05758_);
  and (_10866_, _10865_, _10864_);
  nor (_10867_, _10866_, _10862_);
  nor (_10868_, _10867_, _10604_);
  nor (_10869_, _10868_, _10861_);
  nor (_10870_, _10869_, _10598_);
  or (_10871_, _10870_, _10860_);
  nand (_10872_, _10871_, _10592_);
  and (_10873_, _10872_, _10859_);
  nor (_10874_, _10873_, _10589_);
  or (_10875_, _10874_, _10858_);
  nand (_10876_, _10875_, _10626_);
  and (_10877_, _10876_, _10857_);
  nor (_10878_, _10877_, _10575_);
  and (_10879_, _10877_, _10575_);
  nor (_10880_, _10879_, _10878_);
  or (_10881_, _10880_, _10856_);
  and (_10882_, _10881_, _10855_);
  and (_10883_, _10882_, _10853_);
  nand (_10884_, _10854_, \oc8051_golden_model_1.ACC [6]);
  and (_10885_, _07002_, _05746_);
  not (_10886_, _10885_);
  and (_10887_, _07005_, _05746_);
  nor (_10888_, _06137_, _06841_);
  nor (_10889_, _10888_, _10887_);
  and (_10890_, _10889_, _10886_);
  nand (_10891_, _10890_, _10884_);
  or (_10892_, _10891_, _10883_);
  nor (_10893_, _07883_, _09861_);
  not (_10894_, _10893_);
  nand (_10895_, _07883_, _09861_);
  and (_10896_, _10894_, _10895_);
  nor (_10897_, _07977_, _09906_);
  and (_10898_, _07977_, _09906_);
  nor (_10899_, _10898_, _10897_);
  not (_10900_, _10899_);
  nor (_10901_, _08270_, _09880_);
  nand (_10902_, _08270_, _09880_);
  not (_10903_, _10901_);
  and (_10904_, _10903_, _10902_);
  nor (_10905_, _07353_, _10010_);
  and (_10906_, _07353_, _10010_);
  nor (_10907_, _07530_, _09956_);
  and (_10908_, _07530_, _09956_);
  nor (_10909_, _10907_, _10908_);
  nor (_10910_, _07132_, _05784_);
  and (_10911_, _07132_, _05784_);
  nor (_10912_, _10910_, _10911_);
  and (_10913_, _06931_, \oc8051_golden_model_1.ACC [0]);
  and (_10914_, _10913_, _10912_);
  nor (_10915_, _10914_, _10910_);
  not (_10916_, _10915_);
  and (_10917_, _10916_, _10909_);
  nor (_10918_, _10917_, _10907_);
  nor (_10919_, _10918_, _10906_);
  or (_10920_, _10919_, _10905_);
  and (_10921_, _10920_, _10904_);
  nor (_10922_, _10921_, _10901_);
  nor (_10923_, _10922_, _10900_);
  or (_10924_, _10923_, _10897_);
  nand (_10925_, _10924_, _10896_);
  and (_10926_, _10925_, _10894_);
  nor (_10927_, _10926_, _10674_);
  and (_10928_, _10926_, _10674_);
  or (_10929_, _10928_, _10927_);
  or (_10930_, _10929_, _10890_);
  and (_10931_, _10930_, _10892_);
  and (_10932_, _06103_, _05746_);
  or (_10933_, _10932_, _10931_);
  not (_10934_, _10932_);
  and (_10935_, _09178_, \oc8051_golden_model_1.ACC [6]);
  or (_10936_, _09178_, \oc8051_golden_model_1.ACC [6]);
  not (_10937_, _10935_);
  and (_10938_, _10937_, _10936_);
  and (_10939_, _09179_, \oc8051_golden_model_1.ACC [5]);
  and (_10940_, _08888_, _09906_);
  or (_10941_, _10940_, _10939_);
  or (_10942_, _08937_, _09880_);
  or (_10943_, _09180_, \oc8051_golden_model_1.ACC [4]);
  and (_10944_, _10942_, _10943_);
  and (_10945_, _09181_, \oc8051_golden_model_1.ACC [3]);
  and (_10946_, _08985_, _10010_);
  and (_10947_, _09182_, \oc8051_golden_model_1.ACC [2]);
  and (_10948_, _09030_, _09956_);
  nor (_10949_, _10947_, _10948_);
  not (_10950_, _10949_);
  and (_10951_, _09075_, \oc8051_golden_model_1.ACC [1]);
  or (_10952_, _09075_, \oc8051_golden_model_1.ACC [1]);
  not (_10953_, _10951_);
  and (_10954_, _10953_, _10952_);
  and (_10955_, _09120_, \oc8051_golden_model_1.ACC [0]);
  and (_10956_, _10955_, _10954_);
  nor (_10957_, _10956_, _10951_);
  nor (_10958_, _10957_, _10950_);
  nor (_10959_, _10958_, _10947_);
  nor (_10960_, _10959_, _10946_);
  or (_10961_, _10960_, _10945_);
  nand (_10962_, _10961_, _10944_);
  and (_10963_, _10962_, _10942_);
  nor (_10964_, _10963_, _10941_);
  or (_10965_, _10964_, _10939_);
  and (_10966_, _10965_, _10938_);
  nor (_10967_, _10966_, _10935_);
  and (_10968_, _10967_, _10693_);
  nor (_10969_, _10967_, _10693_);
  or (_10970_, _10969_, _10968_);
  or (_10971_, _10970_, _10934_);
  and (_10972_, _10971_, _06052_);
  and (_10973_, _10972_, _10933_);
  and (_10974_, _06114_, _05746_);
  nor (_10975_, _10974_, _06051_);
  not (_10976_, _10975_);
  nor (_10977_, _07885_, _09861_);
  not (_10978_, _10977_);
  and (_10979_, _07885_, _09861_);
  nor (_10980_, _10979_, _10977_);
  nor (_10981_, _07979_, _09906_);
  and (_10982_, _07979_, _09906_);
  nor (_10983_, _08272_, _09880_);
  not (_10984_, _10983_);
  and (_10985_, _08272_, _09880_);
  nor (_10986_, _10985_, _10983_);
  nor (_10987_, _08028_, _10010_);
  and (_10988_, _08028_, _10010_);
  nor (_10989_, _08176_, _09956_);
  and (_10990_, _08176_, _09956_);
  nor (_10991_, _10990_, _10989_);
  nor (_10992_, _08077_, _05784_);
  and (_10993_, _08077_, _05784_);
  nor (_10994_, _10993_, _10992_);
  and (_10995_, _08127_, \oc8051_golden_model_1.ACC [0]);
  and (_10996_, _10995_, _10994_);
  nor (_10997_, _10996_, _10992_);
  not (_10998_, _10997_);
  and (_10999_, _10998_, _10991_);
  nor (_11000_, _10999_, _10989_);
  nor (_11001_, _11000_, _10988_);
  or (_11002_, _11001_, _10987_);
  nand (_11003_, _11002_, _10986_);
  and (_11004_, _11003_, _10984_);
  nor (_11005_, _11004_, _10982_);
  or (_11006_, _11005_, _10981_);
  nand (_11007_, _11006_, _10980_);
  and (_11008_, _11007_, _10978_);
  and (_11009_, _11008_, _08768_);
  nor (_11010_, _11008_, _08768_);
  or (_11011_, _11010_, _10974_);
  or (_11012_, _11011_, _11009_);
  and (_11013_, _11012_, _10976_);
  or (_11014_, _11013_, _10973_);
  and (_11015_, _05746_, _06107_);
  not (_11016_, _11015_);
  nor (_11017_, _06084_, _09861_);
  not (_11018_, _11017_);
  and (_11019_, _06084_, _09861_);
  nor (_11020_, _11017_, _11019_);
  nor (_11021_, _06359_, _09906_);
  and (_11022_, _06359_, _09906_);
  nor (_11023_, _06758_, _09880_);
  not (_11024_, _11023_);
  and (_11025_, _06758_, _09880_);
  or (_11026_, _11025_, _11023_);
  not (_11027_, _11026_);
  nor (_11028_, _05983_, _10010_);
  and (_11029_, _05983_, _10010_);
  nor (_11030_, _06403_, _09956_);
  and (_11031_, _06403_, _09956_);
  or (_11032_, _11031_, _11030_);
  nor (_11033_, _06799_, _05784_);
  and (_11034_, _06799_, _05784_);
  nor (_11035_, _11033_, _11034_);
  nor (_11036_, _06016_, _05758_);
  and (_11037_, _11036_, _11035_);
  nor (_11038_, _11037_, _11033_);
  nor (_11039_, _11038_, _11032_);
  nor (_11040_, _11039_, _11030_);
  nor (_11041_, _11040_, _11029_);
  or (_11042_, _11041_, _11028_);
  nand (_11043_, _11042_, _11027_);
  and (_11044_, _11043_, _11024_);
  nor (_11045_, _11044_, _11022_);
  or (_11046_, _11045_, _11021_);
  nand (_11047_, _11046_, _11020_);
  and (_11048_, _11047_, _11018_);
  and (_11049_, _11048_, _10705_);
  not (_11050_, _10974_);
  nor (_11051_, _11048_, _10705_);
  or (_11052_, _11051_, _11050_);
  or (_11053_, _11052_, _11049_);
  and (_11054_, _11053_, _11016_);
  and (_11055_, _11054_, _11014_);
  and (_11056_, _11015_, \oc8051_golden_model_1.ACC [6]);
  or (_11057_, _11056_, _06316_);
  or (_11058_, _11057_, _11055_);
  and (_11059_, _06114_, _05495_);
  not (_11060_, _11059_);
  or (_11061_, _10387_, _06718_);
  and (_11062_, _11061_, _11060_);
  and (_11063_, _11062_, _11058_);
  and (_11064_, _06107_, _05495_);
  and (_11065_, _10415_, _05758_);
  and (_11066_, _11065_, _10010_);
  and (_11067_, _11066_, _09880_);
  and (_11068_, _11067_, _09906_);
  and (_11069_, _11068_, _09861_);
  nor (_11070_, _11069_, _08393_);
  and (_11071_, _11069_, _08393_);
  or (_11072_, _11071_, _11070_);
  and (_11073_, _11072_, _11059_);
  or (_11074_, _11073_, _11064_);
  or (_11075_, _11074_, _11063_);
  nand (_11076_, _11064_, _10606_);
  and (_11077_, _11076_, _05653_);
  and (_11078_, _11077_, _11075_);
  and (_11079_, _10456_, _05652_);
  or (_11080_, _11079_, _06047_);
  or (_11081_, _11080_, _11078_);
  and (_11082_, _06114_, _05750_);
  not (_11083_, _11082_);
  and (_11084_, _08279_, _07701_);
  or (_11085_, _10385_, _06048_);
  or (_11086_, _11085_, _11084_);
  and (_11087_, _11086_, _11083_);
  and (_11088_, _11087_, _11081_);
  and (_11089_, _05750_, _06107_);
  and (_11090_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  and (_11091_, _11090_, \oc8051_golden_model_1.ACC [2]);
  and (_11092_, _11091_, \oc8051_golden_model_1.ACC [3]);
  and (_11093_, _11092_, \oc8051_golden_model_1.ACC [4]);
  and (_11094_, _11093_, \oc8051_golden_model_1.ACC [5]);
  and (_11095_, _11094_, \oc8051_golden_model_1.ACC [6]);
  or (_11096_, _11095_, \oc8051_golden_model_1.ACC [7]);
  nand (_11097_, _11095_, \oc8051_golden_model_1.ACC [7]);
  and (_11098_, _11097_, _11096_);
  and (_11099_, _11098_, _11082_);
  or (_11100_, _11099_, _11089_);
  or (_11101_, _11100_, _11088_);
  nand (_11102_, _11089_, _05758_);
  and (_11103_, _11102_, _01336_);
  and (_11104_, _11103_, _11101_);
  or (_11105_, _11104_, _10233_);
  and (_40753_, _11105_, _42882_);
  not (_11106_, \oc8051_golden_model_1.PCON [7]);
  nor (_11107_, _01336_, _11106_);
  nor (_11108_, _07641_, _11106_);
  not (_11109_, _07641_);
  nor (_11110_, _08767_, _11109_);
  or (_11111_, _11110_, _11108_);
  and (_11112_, _11111_, _06292_);
  or (_11113_, _11108_, _07788_);
  and (_11114_, _08549_, _07641_);
  or (_11115_, _11114_, _11108_);
  and (_11116_, _11115_, _06108_);
  and (_11117_, _11116_, _11113_);
  and (_11118_, _08768_, _07641_);
  or (_11119_, _11118_, _11108_);
  and (_11120_, _11119_, _06284_);
  or (_11121_, _11115_, _06020_);
  and (_11122_, _08498_, _07641_);
  or (_11123_, _11122_, _11108_);
  or (_11124_, _11123_, _06954_);
  and (_11125_, _07641_, \oc8051_golden_model_1.ACC [7]);
  or (_11126_, _11125_, _11108_);
  and (_11127_, _11126_, _06938_);
  nor (_11128_, _06938_, _11106_);
  or (_11129_, _11128_, _06102_);
  or (_11130_, _11129_, _11127_);
  and (_11131_, _11130_, _06848_);
  and (_11132_, _11131_, _11124_);
  nor (_11133_, _07785_, _11109_);
  or (_11134_, _11133_, _11108_);
  and (_11135_, _11134_, _06239_);
  or (_11136_, _11135_, _11132_);
  and (_11137_, _11136_, _06220_);
  and (_11138_, _11126_, _06219_);
  or (_11139_, _11138_, _09818_);
  or (_11140_, _11139_, _11137_);
  and (_11141_, _08485_, _07641_);
  or (_11142_, _11108_, _07012_);
  or (_11143_, _11142_, _11141_);
  or (_11144_, _11134_, _09827_);
  and (_11145_, _11144_, _05669_);
  and (_11146_, _11145_, _11143_);
  and (_11147_, _11146_, _11140_);
  and (_11148_, _08738_, _07641_);
  or (_11149_, _11148_, _11108_);
  and (_11150_, _11149_, _09833_);
  or (_11151_, _11150_, _06019_);
  or (_11152_, _11151_, _11147_);
  and (_11153_, _11152_, _11121_);
  or (_11154_, _11153_, _06112_);
  and (_11155_, _08760_, _07641_);
  or (_11156_, _11155_, _11108_);
  or (_11157_, _11156_, _08751_);
  and (_11158_, _11157_, _08756_);
  and (_11159_, _11158_, _11154_);
  or (_11160_, _11159_, _11120_);
  and (_11161_, _11160_, _07032_);
  or (_11162_, _11161_, _11117_);
  and (_11163_, _11162_, _06278_);
  and (_11164_, _11126_, _06277_);
  and (_11165_, _11164_, _11113_);
  or (_11166_, _11165_, _06130_);
  or (_11167_, _11166_, _11163_);
  and (_11168_, _08759_, _07641_);
  or (_11169_, _11108_, _08777_);
  or (_11170_, _11169_, _11168_);
  and (_11171_, _11170_, _08782_);
  and (_11172_, _11171_, _11167_);
  or (_11173_, _11172_, _11112_);
  and (_11174_, _11173_, _06718_);
  and (_11175_, _11123_, _06316_);
  or (_11176_, _11175_, _06047_);
  or (_11177_, _11176_, _11174_);
  and (_11178_, _08279_, _07641_);
  or (_11179_, _11108_, _06048_);
  or (_11180_, _11179_, _11178_);
  and (_11181_, _11180_, _01336_);
  and (_11182_, _11181_, _11177_);
  or (_11183_, _11182_, _11107_);
  and (_40756_, _11183_, _42882_);
  and (_11184_, _01340_, \oc8051_golden_model_1.TMOD [7]);
  not (_11185_, _07653_);
  and (_11186_, _11185_, \oc8051_golden_model_1.TMOD [7]);
  nor (_11187_, _08767_, _11185_);
  or (_11188_, _11187_, _11186_);
  and (_11189_, _11188_, _06292_);
  and (_11190_, _08768_, _07653_);
  or (_11191_, _11190_, _11186_);
  and (_11192_, _11191_, _06284_);
  and (_11193_, _08549_, _07653_);
  or (_11194_, _11193_, _11186_);
  or (_11195_, _11194_, _06020_);
  and (_11196_, _08498_, _07653_);
  or (_11197_, _11196_, _11186_);
  or (_11198_, _11197_, _06954_);
  and (_11199_, _07653_, \oc8051_golden_model_1.ACC [7]);
  or (_11200_, _11199_, _11186_);
  and (_11201_, _11200_, _06938_);
  and (_11202_, _06939_, \oc8051_golden_model_1.TMOD [7]);
  or (_11203_, _11202_, _06102_);
  or (_11204_, _11203_, _11201_);
  and (_11205_, _11204_, _06848_);
  and (_11206_, _11205_, _11198_);
  nor (_11207_, _07785_, _11185_);
  or (_11208_, _11207_, _11186_);
  and (_11209_, _11208_, _06239_);
  or (_11210_, _11209_, _11206_);
  and (_11211_, _11210_, _06220_);
  and (_11212_, _11200_, _06219_);
  or (_11213_, _11212_, _09818_);
  or (_11214_, _11213_, _11211_);
  and (_11215_, _08485_, _07653_);
  or (_11216_, _11186_, _07012_);
  or (_11217_, _11216_, _11215_);
  or (_11218_, _11208_, _09827_);
  and (_11219_, _11218_, _05669_);
  and (_11220_, _11219_, _11217_);
  and (_11221_, _11220_, _11214_);
  and (_11222_, _08738_, _07653_);
  or (_11223_, _11222_, _11186_);
  and (_11224_, _11223_, _09833_);
  or (_11225_, _11224_, _06019_);
  or (_11226_, _11225_, _11221_);
  and (_11227_, _11226_, _11195_);
  or (_11228_, _11227_, _06112_);
  and (_11229_, _08760_, _07653_);
  or (_11230_, _11186_, _08751_);
  or (_11231_, _11230_, _11229_);
  and (_11232_, _11231_, _08756_);
  and (_11233_, _11232_, _11228_);
  or (_11234_, _11233_, _11192_);
  and (_11235_, _11234_, _07032_);
  or (_11236_, _11186_, _07788_);
  and (_11237_, _11194_, _06108_);
  and (_11238_, _11237_, _11236_);
  or (_11239_, _11238_, _11235_);
  and (_11240_, _11239_, _06278_);
  and (_11241_, _11200_, _06277_);
  and (_11242_, _11241_, _11236_);
  or (_11243_, _11242_, _06130_);
  or (_11244_, _11243_, _11240_);
  and (_11245_, _08759_, _07653_);
  or (_11246_, _11186_, _08777_);
  or (_11247_, _11246_, _11245_);
  and (_11248_, _11247_, _08782_);
  and (_11249_, _11248_, _11244_);
  or (_11250_, _11249_, _11189_);
  and (_11251_, _11250_, _06718_);
  and (_11252_, _11197_, _06316_);
  or (_11253_, _11252_, _06047_);
  or (_11254_, _11253_, _11251_);
  and (_11255_, _08279_, _07653_);
  or (_11256_, _11186_, _06048_);
  or (_11257_, _11256_, _11255_);
  and (_11258_, _11257_, _01336_);
  and (_11259_, _11258_, _11254_);
  or (_11260_, _11259_, _11184_);
  and (_40757_, _11260_, _42882_);
  not (_11261_, \oc8051_golden_model_1.DPL [7]);
  nor (_11262_, _01336_, _11261_);
  nor (_11263_, _07733_, _11261_);
  not (_11264_, _07733_);
  nor (_11265_, _08767_, _11264_);
  or (_11266_, _11265_, _11263_);
  and (_11267_, _11266_, _06292_);
  and (_11268_, _08768_, _07733_);
  or (_11269_, _11268_, _11263_);
  and (_11270_, _11269_, _06284_);
  and (_11271_, _08549_, _07733_);
  or (_11272_, _11271_, _11263_);
  or (_11273_, _11272_, _06020_);
  and (_11274_, _08498_, _07733_);
  or (_11275_, _11274_, _11263_);
  or (_11276_, _11275_, _06954_);
  and (_11277_, _07733_, \oc8051_golden_model_1.ACC [7]);
  or (_11278_, _11277_, _11263_);
  and (_11279_, _11278_, _06938_);
  nor (_11280_, _06938_, _11261_);
  or (_11281_, _11280_, _06102_);
  or (_11282_, _11281_, _11279_);
  and (_11283_, _11282_, _06848_);
  and (_11284_, _11283_, _11276_);
  nor (_11285_, _07785_, _11264_);
  or (_11286_, _11285_, _11263_);
  and (_11287_, _11286_, _06239_);
  or (_11288_, _11287_, _06219_);
  or (_11289_, _11288_, _11284_);
  nor (_11290_, _05701_, _05662_);
  not (_11291_, _11290_);
  or (_11292_, _11278_, _06220_);
  and (_11293_, _11292_, _11291_);
  and (_11294_, _11293_, _11289_);
  and (_11295_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_11296_, _11295_, \oc8051_golden_model_1.DPL [2]);
  and (_11297_, _11296_, \oc8051_golden_model_1.DPL [3]);
  and (_11298_, _11297_, \oc8051_golden_model_1.DPL [4]);
  and (_11299_, _11298_, \oc8051_golden_model_1.DPL [5]);
  and (_11300_, _11299_, \oc8051_golden_model_1.DPL [6]);
  nor (_11301_, _11300_, \oc8051_golden_model_1.DPL [7]);
  and (_11302_, _11300_, \oc8051_golden_model_1.DPL [7]);
  nor (_11303_, _11302_, _11301_);
  and (_11304_, _11303_, _11290_);
  or (_11305_, _11304_, _11294_);
  and (_11306_, _11305_, _06111_);
  nor (_11307_, _08332_, _06111_);
  or (_11308_, _11307_, _09818_);
  or (_11309_, _11308_, _11306_);
  and (_11310_, _08485_, _07733_);
  or (_11311_, _11263_, _07012_);
  or (_11312_, _11311_, _11310_);
  or (_11313_, _11286_, _09827_);
  and (_11314_, _11313_, _05669_);
  and (_11315_, _11314_, _11312_);
  and (_11316_, _11315_, _11309_);
  and (_11317_, _08738_, _07733_);
  or (_11318_, _11317_, _11263_);
  and (_11319_, _11318_, _09833_);
  or (_11320_, _11319_, _06019_);
  or (_11321_, _11320_, _11316_);
  and (_11322_, _11321_, _11273_);
  or (_11323_, _11322_, _06112_);
  and (_11324_, _08760_, _07733_);
  or (_11325_, _11263_, _08751_);
  or (_11326_, _11325_, _11324_);
  and (_11327_, _11326_, _08756_);
  and (_11328_, _11327_, _11323_);
  or (_11329_, _11328_, _11270_);
  and (_11330_, _11329_, _07032_);
  or (_11331_, _11263_, _07788_);
  and (_11332_, _11272_, _06108_);
  and (_11333_, _11332_, _11331_);
  or (_11334_, _11333_, _11330_);
  and (_11335_, _11334_, _06278_);
  and (_11336_, _11278_, _06277_);
  and (_11337_, _11336_, _11331_);
  or (_11338_, _11337_, _06130_);
  or (_11339_, _11338_, _11335_);
  and (_11340_, _08759_, _07733_);
  or (_11341_, _11263_, _08777_);
  or (_11342_, _11341_, _11340_);
  and (_11343_, _11342_, _08782_);
  and (_11344_, _11343_, _11339_);
  or (_11345_, _11344_, _11267_);
  and (_11346_, _11345_, _06718_);
  and (_11347_, _11275_, _06316_);
  or (_11348_, _11347_, _06047_);
  or (_11349_, _11348_, _11346_);
  and (_11350_, _08279_, _07733_);
  or (_11351_, _11263_, _06048_);
  or (_11352_, _11351_, _11350_);
  and (_11353_, _11352_, _01336_);
  and (_11354_, _11353_, _11349_);
  or (_11355_, _11354_, _11262_);
  and (_40758_, _11355_, _42882_);
  not (_11356_, \oc8051_golden_model_1.DPH [7]);
  nor (_11357_, _01336_, _11356_);
  nor (_11358_, _07802_, _11356_);
  not (_11359_, _07724_);
  nor (_11360_, _08767_, _11359_);
  or (_11361_, _11360_, _11358_);
  and (_11362_, _11361_, _06292_);
  and (_11363_, _08768_, _07724_);
  or (_11364_, _11363_, _11358_);
  and (_11365_, _11364_, _06284_);
  and (_11366_, _08549_, _07802_);
  or (_11367_, _11366_, _11358_);
  or (_11368_, _11367_, _06020_);
  and (_11369_, _08498_, _07724_);
  or (_11370_, _11369_, _11358_);
  or (_11371_, _11370_, _06954_);
  and (_11372_, _07802_, \oc8051_golden_model_1.ACC [7]);
  or (_11373_, _11372_, _11358_);
  and (_11374_, _11373_, _06938_);
  nor (_11375_, _06938_, _11356_);
  or (_11376_, _11375_, _06102_);
  or (_11377_, _11376_, _11374_);
  and (_11378_, _11377_, _06848_);
  and (_11379_, _11378_, _11371_);
  nor (_11380_, _07785_, _11359_);
  or (_11381_, _11380_, _11358_);
  and (_11382_, _11381_, _06239_);
  or (_11383_, _11382_, _06219_);
  or (_11384_, _11383_, _11379_);
  or (_11385_, _11373_, _06220_);
  and (_11386_, _11385_, _11291_);
  and (_11387_, _11386_, _11384_);
  and (_11388_, _11302_, \oc8051_golden_model_1.DPH [0]);
  and (_11389_, _11388_, \oc8051_golden_model_1.DPH [1]);
  and (_11390_, _11389_, \oc8051_golden_model_1.DPH [2]);
  and (_11391_, _11390_, \oc8051_golden_model_1.DPH [3]);
  and (_11392_, _11391_, \oc8051_golden_model_1.DPH [4]);
  and (_11393_, _11392_, \oc8051_golden_model_1.DPH [5]);
  and (_11394_, _11393_, \oc8051_golden_model_1.DPH [6]);
  nand (_11395_, _11394_, \oc8051_golden_model_1.DPH [7]);
  or (_11396_, _11394_, \oc8051_golden_model_1.DPH [7]);
  and (_11397_, _11396_, _11290_);
  and (_11398_, _11397_, _11395_);
  or (_11399_, _11398_, _11387_);
  and (_11400_, _11399_, _06111_);
  and (_11401_, _06110_, _05952_);
  or (_11402_, _11401_, _09818_);
  or (_11403_, _11402_, _11400_);
  or (_11404_, _11358_, _07012_);
  and (_11405_, _08485_, _07802_);
  or (_11406_, _11405_, _11404_);
  or (_11407_, _11381_, _09827_);
  and (_11408_, _11407_, _05669_);
  and (_11409_, _11408_, _11406_);
  and (_11410_, _11409_, _11403_);
  and (_11411_, _08738_, _07724_);
  or (_11412_, _11411_, _11358_);
  and (_11413_, _11412_, _09833_);
  or (_11414_, _11413_, _06019_);
  or (_11415_, _11414_, _11410_);
  and (_11416_, _11415_, _11368_);
  or (_11417_, _11416_, _06112_);
  and (_11418_, _08760_, _07724_);
  or (_11419_, _11358_, _08751_);
  or (_11420_, _11419_, _11418_);
  and (_11421_, _11420_, _08756_);
  and (_11422_, _11421_, _11417_);
  or (_11423_, _11422_, _11365_);
  and (_11424_, _11423_, _07032_);
  or (_11425_, _11358_, _07788_);
  and (_11426_, _11367_, _06108_);
  and (_11427_, _11426_, _11425_);
  or (_11428_, _11427_, _11424_);
  and (_11429_, _11428_, _06278_);
  and (_11430_, _11373_, _06277_);
  and (_11431_, _11430_, _11425_);
  or (_11432_, _11431_, _06130_);
  or (_11433_, _11432_, _11429_);
  and (_11434_, _08759_, _07724_);
  or (_11435_, _11358_, _08777_);
  or (_11436_, _11435_, _11434_);
  and (_11437_, _11436_, _08782_);
  and (_11438_, _11437_, _11433_);
  or (_11439_, _11438_, _11362_);
  and (_11440_, _11439_, _06718_);
  and (_11441_, _11370_, _06316_);
  or (_11442_, _11441_, _06047_);
  or (_11443_, _11442_, _11440_);
  and (_11444_, _08279_, _07724_);
  or (_11445_, _11358_, _06048_);
  or (_11446_, _11445_, _11444_);
  and (_11447_, _11446_, _01336_);
  and (_11448_, _11447_, _11443_);
  or (_11449_, _11448_, _11357_);
  and (_40759_, _11449_, _42882_);
  and (_11450_, _01340_, \oc8051_golden_model_1.TL1 [7]);
  not (_11451_, _07667_);
  and (_11452_, _11451_, \oc8051_golden_model_1.TL1 [7]);
  nor (_11453_, _08767_, _11451_);
  or (_11454_, _11453_, _11452_);
  and (_11455_, _11454_, _06292_);
  and (_11456_, _08768_, _07667_);
  or (_11457_, _11456_, _11452_);
  and (_11458_, _11457_, _06284_);
  and (_11459_, _08549_, _07667_);
  or (_11460_, _11459_, _11452_);
  or (_11461_, _11460_, _06020_);
  and (_11462_, _08498_, _07667_);
  or (_11463_, _11462_, _11452_);
  or (_11464_, _11463_, _06954_);
  and (_11465_, _07667_, \oc8051_golden_model_1.ACC [7]);
  or (_11466_, _11465_, _11452_);
  and (_11467_, _11466_, _06938_);
  and (_11468_, _06939_, \oc8051_golden_model_1.TL1 [7]);
  or (_11469_, _11468_, _06102_);
  or (_11470_, _11469_, _11467_);
  and (_11471_, _11470_, _06848_);
  and (_11472_, _11471_, _11464_);
  nor (_11473_, _07785_, _11451_);
  or (_11474_, _11473_, _11452_);
  and (_11475_, _11474_, _06239_);
  or (_11476_, _11475_, _11472_);
  and (_11477_, _11476_, _06220_);
  and (_11478_, _11466_, _06219_);
  or (_11479_, _11478_, _09818_);
  or (_11480_, _11479_, _11477_);
  and (_11481_, _08485_, _07667_);
  or (_11482_, _11452_, _07012_);
  or (_11483_, _11482_, _11481_);
  or (_11484_, _11474_, _09827_);
  and (_11485_, _11484_, _05669_);
  and (_11486_, _11485_, _11483_);
  and (_11487_, _11486_, _11480_);
  and (_11488_, _08738_, _07667_);
  or (_11489_, _11488_, _11452_);
  and (_11490_, _11489_, _09833_);
  or (_11491_, _11490_, _06019_);
  or (_11492_, _11491_, _11487_);
  and (_11493_, _11492_, _11461_);
  or (_11494_, _11493_, _06112_);
  and (_11495_, _08760_, _07667_);
  or (_11496_, _11495_, _11452_);
  or (_11497_, _11496_, _08751_);
  and (_11498_, _11497_, _08756_);
  and (_11499_, _11498_, _11494_);
  or (_11500_, _11499_, _11458_);
  and (_11501_, _11500_, _07032_);
  or (_11502_, _11452_, _07788_);
  and (_11503_, _11460_, _06108_);
  and (_11504_, _11503_, _11502_);
  or (_11505_, _11504_, _11501_);
  and (_11506_, _11505_, _06278_);
  and (_11507_, _11466_, _06277_);
  and (_11508_, _11507_, _11502_);
  or (_11509_, _11508_, _06130_);
  or (_11510_, _11509_, _11506_);
  and (_11511_, _08759_, _07667_);
  or (_11512_, _11452_, _08777_);
  or (_11513_, _11512_, _11511_);
  and (_11514_, _11513_, _08782_);
  and (_11515_, _11514_, _11510_);
  or (_11516_, _11515_, _11455_);
  and (_11517_, _11516_, _06718_);
  and (_11518_, _11463_, _06316_);
  or (_11519_, _11518_, _06047_);
  or (_11520_, _11519_, _11517_);
  and (_11521_, _08279_, _07667_);
  or (_11522_, _11452_, _06048_);
  or (_11523_, _11522_, _11521_);
  and (_11524_, _11523_, _01336_);
  and (_11525_, _11524_, _11520_);
  or (_11526_, _11525_, _11450_);
  and (_40760_, _11526_, _42882_);
  and (_11527_, _01340_, \oc8051_golden_model_1.TL0 [7]);
  not (_11528_, _07659_);
  and (_11529_, _11528_, \oc8051_golden_model_1.TL0 [7]);
  nor (_11530_, _08767_, _11528_);
  or (_11531_, _11530_, _11529_);
  and (_11532_, _11531_, _06292_);
  and (_11533_, _08768_, _07659_);
  or (_11534_, _11533_, _11529_);
  and (_11535_, _11534_, _06284_);
  and (_11536_, _08549_, _07659_);
  or (_11537_, _11536_, _11529_);
  or (_11538_, _11537_, _06020_);
  and (_11539_, _08498_, _07659_);
  or (_11540_, _11539_, _11529_);
  or (_11541_, _11540_, _06954_);
  and (_11542_, _07659_, \oc8051_golden_model_1.ACC [7]);
  or (_11543_, _11542_, _11529_);
  and (_11544_, _11543_, _06938_);
  and (_11545_, _06939_, \oc8051_golden_model_1.TL0 [7]);
  or (_11546_, _11545_, _06102_);
  or (_11547_, _11546_, _11544_);
  and (_11548_, _11547_, _06848_);
  and (_11549_, _11548_, _11541_);
  nor (_11550_, _07785_, _11528_);
  or (_11551_, _11550_, _11529_);
  and (_11552_, _11551_, _06239_);
  or (_11553_, _11552_, _11549_);
  and (_11554_, _11553_, _06220_);
  and (_11555_, _11543_, _06219_);
  or (_11556_, _11555_, _09818_);
  or (_11557_, _11556_, _11554_);
  and (_11558_, _08485_, _07659_);
  or (_11559_, _11529_, _07012_);
  or (_11560_, _11559_, _11558_);
  or (_11561_, _11551_, _09827_);
  and (_11562_, _11561_, _05669_);
  and (_11563_, _11562_, _11560_);
  and (_11564_, _11563_, _11557_);
  and (_11565_, _08738_, _07659_);
  or (_11566_, _11565_, _11529_);
  and (_11567_, _11566_, _09833_);
  or (_11568_, _11567_, _06019_);
  or (_11569_, _11568_, _11564_);
  and (_11570_, _11569_, _11538_);
  or (_11571_, _11570_, _06112_);
  and (_11572_, _08760_, _07659_);
  or (_11573_, _11529_, _08751_);
  or (_11574_, _11573_, _11572_);
  and (_11575_, _11574_, _08756_);
  and (_11576_, _11575_, _11571_);
  or (_11577_, _11576_, _11535_);
  and (_11578_, _11577_, _07032_);
  or (_11579_, _11529_, _07788_);
  and (_11580_, _11537_, _06108_);
  and (_11581_, _11580_, _11579_);
  or (_11582_, _11581_, _11578_);
  and (_11583_, _11582_, _06278_);
  and (_11584_, _11543_, _06277_);
  and (_11585_, _11584_, _11579_);
  or (_11586_, _11585_, _06130_);
  or (_11587_, _11586_, _11583_);
  and (_11588_, _08759_, _07659_);
  or (_11589_, _11529_, _08777_);
  or (_11590_, _11589_, _11588_);
  and (_11591_, _11590_, _08782_);
  and (_11592_, _11591_, _11587_);
  or (_11593_, _11592_, _11532_);
  and (_11594_, _11593_, _06718_);
  and (_11595_, _11540_, _06316_);
  or (_11596_, _11595_, _06047_);
  or (_11597_, _11596_, _11594_);
  and (_11598_, _08279_, _07659_);
  or (_11599_, _11529_, _06048_);
  or (_11600_, _11599_, _11598_);
  and (_11601_, _11600_, _01336_);
  and (_11602_, _11601_, _11597_);
  or (_11603_, _11602_, _11527_);
  and (_40762_, _11603_, _42882_);
  and (_11604_, _01340_, \oc8051_golden_model_1.TCON [7]);
  not (_11605_, _07648_);
  and (_11606_, _11605_, \oc8051_golden_model_1.TCON [7]);
  and (_11607_, _08768_, _07648_);
  or (_11608_, _11607_, _11606_);
  and (_11609_, _11608_, _06284_);
  and (_11610_, _08549_, _07648_);
  or (_11611_, _11610_, _11606_);
  or (_11612_, _11611_, _06020_);
  and (_11613_, _08498_, _07648_);
  or (_11614_, _11613_, _11606_);
  or (_11615_, _11614_, _06954_);
  and (_11616_, _07648_, \oc8051_golden_model_1.ACC [7]);
  or (_11617_, _11616_, _11606_);
  and (_11618_, _11617_, _06938_);
  and (_11619_, _06939_, \oc8051_golden_model_1.TCON [7]);
  or (_11620_, _11619_, _06102_);
  or (_11621_, _11620_, _11618_);
  and (_11622_, _11621_, _06044_);
  and (_11623_, _11622_, _11615_);
  not (_11624_, _08341_);
  and (_11625_, _11624_, \oc8051_golden_model_1.TCON [7]);
  and (_11626_, _08503_, _08341_);
  or (_11627_, _11626_, _11625_);
  and (_11628_, _11627_, _06043_);
  or (_11629_, _11628_, _06239_);
  or (_11630_, _11629_, _11623_);
  nor (_11631_, _07785_, _11605_);
  or (_11632_, _11631_, _11606_);
  or (_11633_, _11632_, _06848_);
  and (_11634_, _11633_, _11630_);
  or (_11635_, _11634_, _06219_);
  or (_11636_, _11617_, _06220_);
  and (_11637_, _11636_, _06040_);
  and (_11638_, _11637_, _11635_);
  and (_11639_, _08374_, _08341_);
  or (_11640_, _11639_, _11625_);
  and (_11641_, _11640_, _06039_);
  or (_11642_, _11641_, _06032_);
  or (_11643_, _11642_, _11638_);
  or (_11644_, _11625_, _08519_);
  and (_11645_, _11644_, _11627_);
  or (_11646_, _11645_, _06033_);
  and (_11647_, _11646_, _06027_);
  and (_11648_, _11647_, _11643_);
  and (_11649_, _08376_, _08341_);
  or (_11650_, _11649_, _11625_);
  and (_11651_, _11650_, _06026_);
  or (_11652_, _11651_, _09818_);
  or (_11653_, _11652_, _11648_);
  and (_11654_, _08485_, _07648_);
  or (_11655_, _11606_, _07012_);
  or (_11656_, _11655_, _11654_);
  or (_11657_, _11632_, _09827_);
  and (_11658_, _11657_, _05669_);
  and (_11659_, _11658_, _11656_);
  and (_11660_, _11659_, _11653_);
  and (_11661_, _08738_, _07648_);
  or (_11662_, _11661_, _11606_);
  and (_11663_, _11662_, _09833_);
  or (_11664_, _11663_, _06019_);
  or (_11665_, _11664_, _11660_);
  and (_11666_, _11665_, _11612_);
  or (_11667_, _11666_, _06112_);
  and (_11668_, _08760_, _07648_);
  or (_11669_, _11606_, _08751_);
  or (_11670_, _11669_, _11668_);
  and (_11671_, _11670_, _08756_);
  and (_11672_, _11671_, _11667_);
  or (_11673_, _11672_, _11609_);
  and (_11674_, _11673_, _07032_);
  or (_11675_, _11606_, _07788_);
  and (_11676_, _11611_, _06108_);
  and (_11677_, _11676_, _11675_);
  or (_11678_, _11677_, _11674_);
  and (_11679_, _11678_, _06278_);
  and (_11680_, _11617_, _06277_);
  and (_11681_, _11680_, _11675_);
  or (_11682_, _11681_, _06130_);
  or (_11683_, _11682_, _11679_);
  and (_11684_, _08759_, _07648_);
  or (_11685_, _11606_, _08777_);
  or (_11686_, _11685_, _11684_);
  and (_11687_, _11686_, _08782_);
  and (_11688_, _11687_, _11683_);
  nor (_11689_, _08767_, _11605_);
  or (_11690_, _11689_, _11606_);
  and (_11691_, _11690_, _06292_);
  or (_11692_, _11691_, _06316_);
  or (_11693_, _11692_, _11688_);
  or (_11694_, _11614_, _06718_);
  and (_11695_, _11694_, _05653_);
  and (_11696_, _11695_, _11693_);
  and (_11697_, _11640_, _05652_);
  or (_11698_, _11697_, _06047_);
  or (_11699_, _11698_, _11696_);
  and (_11700_, _08279_, _07648_);
  or (_11701_, _11606_, _06048_);
  or (_11702_, _11701_, _11700_);
  and (_11703_, _11702_, _01336_);
  and (_11704_, _11703_, _11699_);
  or (_11705_, _11704_, _11604_);
  and (_40763_, _11705_, _42882_);
  and (_11706_, _01340_, \oc8051_golden_model_1.TH1 [7]);
  not (_11707_, _07670_);
  and (_11708_, _11707_, \oc8051_golden_model_1.TH1 [7]);
  nor (_11709_, _08767_, _11707_);
  or (_11710_, _11709_, _11708_);
  and (_11711_, _11710_, _06292_);
  or (_11712_, _11708_, _07788_);
  and (_11713_, _08549_, _07670_);
  or (_11714_, _11713_, _11708_);
  and (_11715_, _11714_, _06108_);
  and (_11716_, _11715_, _11712_);
  and (_11717_, _08768_, _07670_);
  or (_11718_, _11717_, _11708_);
  and (_11719_, _11718_, _06284_);
  or (_11720_, _11714_, _06020_);
  and (_11721_, _08498_, _07670_);
  or (_11722_, _11721_, _11708_);
  or (_11723_, _11722_, _06954_);
  and (_11724_, _07670_, \oc8051_golden_model_1.ACC [7]);
  or (_11725_, _11724_, _11708_);
  and (_11726_, _11725_, _06938_);
  and (_11727_, _06939_, \oc8051_golden_model_1.TH1 [7]);
  or (_11728_, _11727_, _06102_);
  or (_11729_, _11728_, _11726_);
  and (_11730_, _11729_, _06848_);
  and (_11731_, _11730_, _11723_);
  nor (_11732_, _07785_, _11707_);
  or (_11733_, _11732_, _11708_);
  and (_11734_, _11733_, _06239_);
  or (_11735_, _11734_, _11731_);
  and (_11736_, _11735_, _06220_);
  and (_11737_, _11725_, _06219_);
  or (_11738_, _11737_, _09818_);
  or (_11739_, _11738_, _11736_);
  and (_11740_, _08485_, _07670_);
  or (_11741_, _11708_, _07012_);
  or (_11742_, _11741_, _11740_);
  or (_11743_, _11733_, _09827_);
  and (_11744_, _11743_, _05669_);
  and (_11745_, _11744_, _11742_);
  and (_11746_, _11745_, _11739_);
  and (_11747_, _08738_, _07670_);
  or (_11748_, _11747_, _11708_);
  and (_11749_, _11748_, _09833_);
  or (_11750_, _11749_, _06019_);
  or (_11751_, _11750_, _11746_);
  and (_11752_, _11751_, _11720_);
  or (_11753_, _11752_, _06112_);
  and (_11754_, _08760_, _07670_);
  or (_11755_, _11754_, _11708_);
  or (_11756_, _11755_, _08751_);
  and (_11757_, _11756_, _08756_);
  and (_11758_, _11757_, _11753_);
  or (_11759_, _11758_, _11719_);
  and (_11760_, _11759_, _07032_);
  or (_11761_, _11760_, _11716_);
  and (_11762_, _11761_, _06278_);
  and (_11763_, _11725_, _06277_);
  and (_11764_, _11763_, _11712_);
  or (_11765_, _11764_, _06130_);
  or (_11766_, _11765_, _11762_);
  and (_11767_, _08759_, _07670_);
  or (_11768_, _11708_, _08777_);
  or (_11769_, _11768_, _11767_);
  and (_11770_, _11769_, _08782_);
  and (_11771_, _11770_, _11766_);
  or (_11772_, _11771_, _11711_);
  and (_11773_, _11772_, _06718_);
  and (_11774_, _11722_, _06316_);
  or (_11775_, _11774_, _06047_);
  or (_11776_, _11775_, _11773_);
  and (_11777_, _08279_, _07670_);
  or (_11778_, _11708_, _06048_);
  or (_11779_, _11778_, _11777_);
  and (_11780_, _11779_, _01336_);
  and (_11781_, _11780_, _11776_);
  or (_11782_, _11781_, _11706_);
  and (_40764_, _11782_, _42882_);
  and (_11783_, _01340_, \oc8051_golden_model_1.TH0 [7]);
  not (_11784_, _07663_);
  and (_11785_, _11784_, \oc8051_golden_model_1.TH0 [7]);
  nor (_11786_, _08767_, _11784_);
  or (_11787_, _11786_, _11785_);
  and (_11788_, _11787_, _06292_);
  and (_11789_, _08768_, _07663_);
  or (_11790_, _11789_, _11785_);
  and (_11791_, _11790_, _06284_);
  and (_11792_, _08549_, _07663_);
  or (_11793_, _11792_, _11785_);
  or (_11794_, _11793_, _06020_);
  and (_11795_, _08498_, _07663_);
  or (_11796_, _11795_, _11785_);
  or (_11797_, _11796_, _06954_);
  and (_11798_, _07663_, \oc8051_golden_model_1.ACC [7]);
  or (_11799_, _11798_, _11785_);
  and (_11800_, _11799_, _06938_);
  and (_11801_, _06939_, \oc8051_golden_model_1.TH0 [7]);
  or (_11802_, _11801_, _06102_);
  or (_11803_, _11802_, _11800_);
  and (_11804_, _11803_, _06848_);
  and (_11805_, _11804_, _11797_);
  nor (_11806_, _07785_, _11784_);
  or (_11807_, _11806_, _11785_);
  and (_11808_, _11807_, _06239_);
  or (_11809_, _11808_, _11805_);
  and (_11810_, _11809_, _06220_);
  and (_11811_, _11799_, _06219_);
  or (_11812_, _11811_, _09818_);
  or (_11813_, _11812_, _11810_);
  and (_11814_, _08485_, _07663_);
  or (_11815_, _11785_, _07012_);
  or (_11816_, _11815_, _11814_);
  or (_11817_, _11807_, _09827_);
  and (_11818_, _11817_, _05669_);
  and (_11819_, _11818_, _11816_);
  and (_11820_, _11819_, _11813_);
  and (_11821_, _08738_, _07663_);
  or (_11822_, _11821_, _11785_);
  and (_11823_, _11822_, _09833_);
  or (_11824_, _11823_, _06019_);
  or (_11825_, _11824_, _11820_);
  and (_11826_, _11825_, _11794_);
  or (_11827_, _11826_, _06112_);
  and (_11828_, _08760_, _07663_);
  or (_11829_, _11785_, _08751_);
  or (_11830_, _11829_, _11828_);
  and (_11831_, _11830_, _08756_);
  and (_11832_, _11831_, _11827_);
  or (_11833_, _11832_, _11791_);
  and (_11834_, _11833_, _07032_);
  or (_11835_, _11785_, _07788_);
  and (_11836_, _11793_, _06108_);
  and (_11837_, _11836_, _11835_);
  or (_11838_, _11837_, _11834_);
  and (_11839_, _11838_, _06278_);
  and (_11840_, _11799_, _06277_);
  and (_11841_, _11840_, _11835_);
  or (_11842_, _11841_, _06130_);
  or (_11843_, _11842_, _11839_);
  and (_11844_, _08759_, _07663_);
  or (_11845_, _11785_, _08777_);
  or (_11846_, _11845_, _11844_);
  and (_11847_, _11846_, _08782_);
  and (_11848_, _11847_, _11843_);
  or (_11849_, _11848_, _11788_);
  and (_11850_, _11849_, _06718_);
  and (_11851_, _11796_, _06316_);
  or (_11852_, _11851_, _06047_);
  or (_11853_, _11852_, _11850_);
  and (_11854_, _08279_, _07663_);
  or (_11855_, _11785_, _06048_);
  or (_11856_, _11855_, _11854_);
  and (_11857_, _11856_, _01336_);
  and (_11858_, _11857_, _11853_);
  or (_11859_, _11858_, _11783_);
  and (_40765_, _11859_, _42882_);
  not (_11860_, _05331_);
  and (_11861_, _08387_, _11860_);
  and (_11862_, _11861_, \oc8051_golden_model_1.PC [7]);
  and (_11863_, _11862_, _09201_);
  and (_11864_, _11863_, \oc8051_golden_model_1.PC [10]);
  and (_11865_, _11864_, \oc8051_golden_model_1.PC [11]);
  and (_11866_, _11865_, \oc8051_golden_model_1.PC [12]);
  and (_11867_, _11866_, \oc8051_golden_model_1.PC [13]);
  and (_11868_, _11867_, \oc8051_golden_model_1.PC [14]);
  or (_11869_, _11868_, \oc8051_golden_model_1.PC [15]);
  nand (_11870_, _11868_, \oc8051_golden_model_1.PC [15]);
  and (_11871_, _11870_, _11869_);
  and (_11872_, _10934_, _10890_);
  or (_11873_, _11872_, _11871_);
  nor (_11874_, _09206_, \oc8051_golden_model_1.PC [14]);
  nor (_11875_, _11874_, _09207_);
  and (_11876_, _11875_, _05952_);
  nor (_11877_, _11875_, _05952_);
  nor (_11878_, _11877_, _11876_);
  nor (_11879_, _09205_, \oc8051_golden_model_1.PC [13]);
  nor (_11880_, _11879_, _09206_);
  and (_11881_, _11880_, _05952_);
  nor (_11882_, _11880_, _05952_);
  nor (_11883_, _09204_, \oc8051_golden_model_1.PC [12]);
  nor (_11884_, _11883_, _09205_);
  and (_11885_, _11884_, _05952_);
  nor (_11886_, _09209_, \oc8051_golden_model_1.PC [10]);
  nor (_11887_, _11886_, _09210_);
  and (_11888_, _11887_, _05952_);
  not (_11889_, _11888_);
  nor (_11890_, _09210_, \oc8051_golden_model_1.PC [11]);
  nor (_11891_, _11890_, _09211_);
  and (_11892_, _11891_, _05952_);
  nor (_11893_, _11891_, _05952_);
  nor (_11894_, _11893_, _11892_);
  nor (_11895_, _11887_, _05952_);
  nor (_11896_, _11895_, _11888_);
  and (_11897_, _11896_, _11894_);
  and (_11898_, _08389_, \oc8051_golden_model_1.PC [8]);
  nor (_11899_, _11898_, \oc8051_golden_model_1.PC [9]);
  nor (_11900_, _11899_, _09209_);
  and (_11901_, _11900_, _05952_);
  nor (_11902_, _11900_, _05952_);
  nor (_11903_, _11902_, _11901_);
  and (_11904_, _08391_, _05952_);
  nor (_11905_, _08391_, _05952_);
  and (_11906_, _08386_, _05850_);
  nor (_11907_, _11906_, \oc8051_golden_model_1.PC [6]);
  nor (_11908_, _11907_, _08388_);
  not (_11909_, _11908_);
  nor (_11910_, _11909_, _06084_);
  and (_11911_, _11909_, _06084_);
  nor (_11912_, _11911_, _11910_);
  not (_11913_, _11912_);
  and (_11914_, _05850_, \oc8051_golden_model_1.PC [4]);
  nor (_11915_, _11914_, \oc8051_golden_model_1.PC [5]);
  nor (_11916_, _11915_, _11906_);
  not (_11917_, _11916_);
  nor (_11918_, _11917_, _06359_);
  and (_11919_, _11917_, _06359_);
  nor (_11920_, _05850_, \oc8051_golden_model_1.PC [4]);
  nor (_11921_, _11920_, _11914_);
  not (_11922_, _11921_);
  nor (_11923_, _11922_, _06758_);
  nor (_11924_, _05983_, _06148_);
  and (_11925_, _05983_, _06148_);
  nor (_11926_, _06403_, _05804_);
  nor (_11927_, _06799_, \oc8051_golden_model_1.PC [1]);
  nor (_11928_, _06016_, _05346_);
  and (_11929_, _06799_, \oc8051_golden_model_1.PC [1]);
  nor (_11930_, _11929_, _11927_);
  and (_11931_, _11930_, _11928_);
  nor (_11932_, _11931_, _11927_);
  and (_11933_, _06403_, _05804_);
  nor (_11934_, _11933_, _11926_);
  not (_11935_, _11934_);
  nor (_11936_, _11935_, _11932_);
  nor (_11937_, _11936_, _11926_);
  nor (_11938_, _11937_, _11925_);
  nor (_11939_, _11938_, _11924_);
  and (_11940_, _11922_, _06758_);
  nor (_11941_, _11940_, _11923_);
  not (_11942_, _11941_);
  nor (_11943_, _11942_, _11939_);
  nor (_11944_, _11943_, _11923_);
  nor (_11945_, _11944_, _11919_);
  nor (_11946_, _11945_, _11918_);
  nor (_11947_, _11946_, _11913_);
  nor (_11948_, _11947_, _11910_);
  nor (_11949_, _11948_, _11905_);
  or (_11950_, _11949_, _11904_);
  nor (_11951_, _08389_, \oc8051_golden_model_1.PC [8]);
  nor (_11952_, _11951_, _11898_);
  and (_11953_, _11952_, _05952_);
  nor (_11954_, _11952_, _05952_);
  nor (_11955_, _11954_, _11953_);
  and (_11956_, _11955_, _11950_);
  and (_11957_, _11956_, _11903_);
  and (_11958_, _11957_, _11897_);
  nor (_11959_, _11953_, _11901_);
  not (_11960_, _11959_);
  and (_11961_, _11960_, _11897_);
  or (_11962_, _11961_, _11892_);
  nor (_11963_, _11962_, _11958_);
  and (_11964_, _11963_, _11889_);
  nor (_11965_, _11884_, _05952_);
  nor (_11966_, _11965_, _11885_);
  not (_11967_, _11966_);
  nor (_11968_, _11967_, _11964_);
  nor (_11969_, _11968_, _11885_);
  nor (_11970_, _11969_, _11882_);
  nor (_11971_, _11970_, _11881_);
  not (_11972_, _11971_);
  and (_11973_, _11972_, _11878_);
  nor (_11974_, _11973_, _11876_);
  nor (_11975_, _09216_, _05952_);
  and (_11976_, _09216_, _05952_);
  nor (_11977_, _11976_, _11975_);
  and (_11978_, _11977_, _11974_);
  nor (_11979_, _11977_, _11974_);
  or (_11980_, _11979_, _11978_);
  or (_11981_, _11980_, _10606_);
  and (_11982_, _05739_, _05650_);
  or (_11983_, _09216_, \oc8051_golden_model_1.PSW [7]);
  and (_11984_, _11983_, _11982_);
  and (_11985_, _11984_, _11981_);
  nor (_11986_, _10781_, _06290_);
  not (_11987_, _11986_);
  or (_11988_, _06093_, _06135_);
  and (_11989_, _11988_, _05739_);
  not (_11990_, _11989_);
  and (_11991_, _07002_, _05739_);
  nor (_11992_, _10775_, _11991_);
  and (_11993_, _11992_, _11990_);
  or (_11994_, _11993_, _11871_);
  nor (_11995_, _06093_, _06229_);
  nor (_11996_, _11995_, _06656_);
  not (_11997_, _11996_);
  and (_11998_, _06227_, _05735_);
  and (_11999_, _07002_, _05735_);
  or (_12000_, _11999_, _10731_);
  nor (_12001_, _12000_, _11998_);
  and (_12002_, _12001_, _11997_);
  or (_12003_, _12002_, _11871_);
  not (_12004_, _07248_);
  nor (_12005_, _11988_, _12004_);
  nor (_12006_, _12005_, _06644_);
  not (_12007_, _12006_);
  or (_12008_, _12007_, _11871_);
  or (_12009_, _09216_, _08742_);
  not (_12010_, _09227_);
  nor (_12011_, _12010_, _05669_);
  nor (_12012_, _05685_, _05662_);
  not (_12013_, _12012_);
  and (_12014_, _09202_, _09139_);
  and (_12015_, _12014_, \oc8051_golden_model_1.PC [11]);
  and (_12016_, _12015_, \oc8051_golden_model_1.PC [12]);
  and (_12017_, _12016_, \oc8051_golden_model_1.PC [13]);
  and (_12018_, _12017_, \oc8051_golden_model_1.PC [14]);
  nor (_12019_, _12017_, \oc8051_golden_model_1.PC [14]);
  nor (_12020_, _12019_, _12018_);
  not (_12021_, _12020_);
  nor (_12022_, _12021_, _08332_);
  and (_12023_, _12021_, _08332_);
  nor (_12024_, _12023_, _12022_);
  not (_12025_, _12024_);
  nor (_12026_, _12016_, \oc8051_golden_model_1.PC [13]);
  nor (_12027_, _12026_, _12017_);
  not (_12028_, _12027_);
  nor (_12029_, _12028_, _08332_);
  and (_12030_, _12028_, _08332_);
  nor (_12031_, _12015_, \oc8051_golden_model_1.PC [12]);
  nor (_12032_, _12031_, _12016_);
  not (_12033_, _12032_);
  nor (_12034_, _12033_, _08332_);
  nor (_12035_, _12014_, \oc8051_golden_model_1.PC [11]);
  nor (_12036_, _12035_, _12015_);
  not (_12037_, _12036_);
  nor (_12038_, _12037_, _08332_);
  and (_12039_, _12037_, _08332_);
  nor (_12040_, _12039_, _12038_);
  and (_12041_, _09201_, _09139_);
  nor (_12042_, _12041_, \oc8051_golden_model_1.PC [10]);
  nor (_12043_, _12042_, _12014_);
  not (_12044_, _12043_);
  nor (_12045_, _12044_, _08332_);
  and (_12046_, _12044_, _08332_);
  nor (_12047_, _12046_, _12045_);
  and (_12048_, _12047_, _12040_);
  and (_12049_, _09139_, \oc8051_golden_model_1.PC [8]);
  nor (_12050_, _12049_, \oc8051_golden_model_1.PC [9]);
  nor (_12051_, _12050_, _12041_);
  not (_12052_, _12051_);
  nor (_12053_, _12052_, _08332_);
  and (_12054_, _12052_, _08332_);
  nor (_12055_, _12054_, _12053_);
  nor (_12056_, _09142_, _08332_);
  and (_12057_, _09142_, _08332_);
  nor (_12058_, _12057_, _12056_);
  not (_12059_, _12058_);
  and (_12060_, _09137_, _08386_);
  nor (_12061_, _12060_, \oc8051_golden_model_1.PC [6]);
  nor (_12062_, _12061_, _09138_);
  not (_12063_, _12062_);
  nor (_12064_, _12063_, _08647_);
  and (_12065_, _12063_, _08647_);
  nor (_12066_, _12065_, _12064_);
  and (_12067_, _09137_, \oc8051_golden_model_1.PC [4]);
  nor (_12068_, _12067_, \oc8051_golden_model_1.PC [5]);
  nor (_12069_, _12068_, _12060_);
  not (_12070_, _12069_);
  nor (_12071_, _12070_, _08612_);
  and (_12072_, _12070_, _08612_);
  nor (_12073_, _09137_, \oc8051_golden_model_1.PC [4]);
  nor (_12074_, _12073_, _12067_);
  not (_12075_, _12074_);
  nor (_12076_, _12075_, _08581_);
  nor (_12077_, _09136_, \oc8051_golden_model_1.PC [3]);
  nor (_12078_, _12077_, _09137_);
  not (_12079_, _12078_);
  nor (_12080_, _12079_, _06215_);
  and (_12081_, _12079_, _06215_);
  nor (_12082_, _05350_, \oc8051_golden_model_1.PC [2]);
  nor (_12083_, _12082_, _09136_);
  not (_12084_, _12083_);
  nor (_12085_, _12084_, _06445_);
  not (_12086_, _05777_);
  nor (_12087_, _06832_, _12086_);
  nor (_12088_, _06633_, \oc8051_golden_model_1.PC [0]);
  and (_12089_, _06832_, _12086_);
  nor (_12090_, _12089_, _12087_);
  and (_12091_, _12090_, _12088_);
  nor (_12092_, _12091_, _12087_);
  and (_12093_, _12084_, _06445_);
  nor (_12094_, _12093_, _12085_);
  not (_12095_, _12094_);
  nor (_12096_, _12095_, _12092_);
  nor (_12097_, _12096_, _12085_);
  nor (_12098_, _12097_, _12081_);
  nor (_12099_, _12098_, _12080_);
  and (_12100_, _12075_, _08581_);
  nor (_12101_, _12100_, _12076_);
  not (_12102_, _12101_);
  nor (_12103_, _12102_, _12099_);
  nor (_12104_, _12103_, _12076_);
  nor (_12105_, _12104_, _12072_);
  or (_12106_, _12105_, _12071_);
  and (_12107_, _12106_, _12066_);
  nor (_12108_, _12107_, _12064_);
  nor (_12109_, _12108_, _12059_);
  nor (_12110_, _12109_, _12056_);
  nor (_12111_, _09139_, \oc8051_golden_model_1.PC [8]);
  nor (_12112_, _12111_, _12049_);
  not (_12113_, _12112_);
  nor (_12114_, _12113_, _08332_);
  and (_12115_, _12113_, _08332_);
  nor (_12116_, _12115_, _12114_);
  not (_12117_, _12116_);
  nor (_12118_, _12117_, _12110_);
  and (_12119_, _12118_, _12055_);
  and (_12120_, _12119_, _12048_);
  nor (_12121_, _12114_, _12053_);
  not (_12122_, _12121_);
  and (_12123_, _12122_, _12048_);
  or (_12124_, _12123_, _12045_);
  or (_12125_, _12124_, _12120_);
  nor (_12126_, _12125_, _12038_);
  and (_12127_, _12033_, _08332_);
  nor (_12128_, _12127_, _12034_);
  not (_12129_, _12128_);
  nor (_12130_, _12129_, _12126_);
  nor (_12131_, _12130_, _12034_);
  nor (_12132_, _12131_, _12030_);
  nor (_12133_, _12132_, _12029_);
  nor (_12134_, _12133_, _12025_);
  nor (_12135_, _12134_, _12022_);
  and (_12136_, _12010_, _08332_);
  nor (_12137_, _12010_, _08332_);
  nor (_12138_, _12137_, _12136_);
  and (_12139_, _12138_, _12135_);
  nor (_12140_, _12138_, _12135_);
  or (_12141_, _12140_, _12139_);
  or (_12142_, _09181_, _05983_);
  or (_12143_, _08985_, _06299_);
  and (_12144_, _12143_, _12142_);
  or (_12145_, _09182_, _06403_);
  or (_12146_, _09030_, _07477_);
  and (_12147_, _12146_, _12145_);
  and (_12148_, _12147_, _12144_);
  nand (_12149_, _09120_, _06016_);
  nand (_12150_, _09074_, _09052_);
  or (_12151_, _12150_, _07076_);
  or (_12152_, _09075_, _06799_);
  and (_12153_, _12152_, _12151_);
  and (_12154_, _12153_, _12149_);
  and (_12155_, _12154_, _12148_);
  or (_12156_, _09120_, _06016_);
  and (_12157_, _08798_, _05952_);
  nor (_12158_, _12157_, _08531_);
  or (_12159_, _09178_, _06084_);
  or (_12160_, _08843_, _07414_);
  and (_12161_, _12160_, _12159_);
  and (_12162_, _12161_, _12158_);
  or (_12163_, _09179_, _06359_);
  or (_12164_, _08888_, _07683_);
  and (_12165_, _12164_, _12163_);
  or (_12166_, _09180_, _06758_);
  or (_12167_, _08937_, _07674_);
  and (_12168_, _12167_, _12166_);
  and (_12169_, _12168_, _12165_);
  and (_12170_, _12169_, _12162_);
  and (_12171_, _12170_, _12156_);
  and (_12172_, _12171_, _12155_);
  or (_12173_, _12172_, _12141_);
  nand (_12174_, _12171_, _12155_);
  or (_12175_, _12174_, _09227_);
  and (_12176_, _12175_, _06104_);
  and (_12177_, _12176_, _12173_);
  and (_12178_, _09216_, _06219_);
  and (_12179_, _06244_, _05690_);
  or (_12180_, _12179_, _09216_);
  nor (_12181_, _05689_, _05662_);
  nor (_12182_, _12181_, _10412_);
  and (_12183_, _07885_, _07787_);
  and (_12184_, _12183_, _08489_);
  and (_12185_, _08127_, _08077_);
  and (_12186_, _08492_, _12185_);
  nand (_12187_, _12186_, _12184_);
  or (_12188_, _12187_, _09227_);
  and (_12189_, _12186_, _12184_);
  or (_12190_, _12189_, _12141_);
  and (_12191_, _12190_, _06102_);
  and (_12192_, _12191_, _12188_);
  and (_12193_, _07132_, _06931_);
  and (_12194_, _07883_, _07785_);
  and (_12195_, _12194_, _12193_);
  and (_12196_, _08290_, _08289_);
  and (_12197_, _12196_, _12195_);
  and (_12198_, _12197_, _09216_);
  nand (_12199_, _12196_, _12195_);
  and (_12200_, _12199_, _11980_);
  or (_12201_, _12200_, _08383_);
  or (_12202_, _12201_, _12198_);
  nor (_12203_, _06933_, _05697_);
  not (_12204_, _12203_);
  and (_12205_, _12204_, _10400_);
  nor (_12206_, _06938_, _06943_);
  or (_12207_, _12206_, _09216_);
  or (_12208_, _06530_, _06943_);
  or (_12209_, _06938_, \oc8051_golden_model_1.PC [15]);
  or (_12210_, _12209_, _12208_);
  or (_12211_, _12210_, _07250_);
  nand (_12212_, _12211_, _12207_);
  nand (_12213_, _12212_, _12205_);
  nor (_12214_, _07250_, _06530_);
  and (_12215_, _12214_, _12205_);
  or (_12216_, _12215_, _11871_);
  and (_12217_, _12216_, _12213_);
  or (_12218_, _12217_, _08384_);
  nor (_12219_, _06948_, _06102_);
  and (_12220_, _12219_, _12218_);
  and (_12221_, _12220_, _12202_);
  or (_12222_, _12221_, _12192_);
  and (_12223_, _12222_, _12182_);
  not (_12224_, _12179_);
  and (_12225_, _12182_, _06949_);
  not (_12226_, _12225_);
  and (_12227_, _12226_, _11871_);
  or (_12228_, _12227_, _12224_);
  or (_12229_, _12228_, _12223_);
  and (_12230_, _12229_, _12180_);
  nor (_12231_, _10378_, _06970_);
  not (_12232_, _12231_);
  or (_12233_, _12232_, _12230_);
  or (_12234_, _12231_, _11871_);
  and (_12235_, _12234_, _06220_);
  and (_12236_, _12235_, _12233_);
  or (_12237_, _12236_, _12178_);
  nor (_12238_, _05693_, _05662_);
  nor (_12239_, _12238_, _10376_);
  and (_12240_, _12239_, _12237_);
  not (_12241_, _12239_);
  and (_12242_, _12241_, _11871_);
  not (_12243_, _05694_);
  nor (_12244_, _06038_, _12243_);
  and (_12245_, _12244_, _06040_);
  not (_12246_, _12245_);
  or (_12247_, _12246_, _12242_);
  or (_12248_, _12247_, _12240_);
  or (_12249_, _12245_, _09216_);
  and (_12250_, _12249_, _12248_);
  not (_12251_, _06138_);
  and (_12252_, _07002_, _06031_);
  and (_12253_, _07005_, _06031_);
  nor (_12254_, _12253_, _12252_);
  and (_12255_, _12254_, _12251_);
  not (_12256_, _12255_);
  or (_12257_, _12256_, _12250_);
  not (_12258_, _06104_);
  not (_12259_, _07786_);
  and (_12260_, _07785_, _05952_);
  nor (_12261_, _12260_, _12259_);
  nor (_12262_, _07883_, _07414_);
  and (_12263_, _07883_, _07414_);
  nor (_12264_, _12263_, _12262_);
  and (_12265_, _12264_, _12261_);
  nor (_12266_, _07977_, _07683_);
  and (_12267_, _07977_, _07683_);
  nor (_12268_, _12267_, _12266_);
  and (_12269_, _08270_, _07674_);
  nor (_12270_, _08270_, _07674_);
  nor (_12271_, _12270_, _12269_);
  and (_12272_, _12271_, _12268_);
  and (_12273_, _12272_, _12265_);
  and (_12274_, _07353_, _06299_);
  nor (_12275_, _07353_, _06299_);
  nor (_12276_, _12275_, _12274_);
  and (_12277_, _07530_, _07477_);
  nor (_12278_, _07530_, _07477_);
  nor (_12279_, _12278_, _12277_);
  and (_12280_, _12279_, _12276_);
  nor (_12281_, _07132_, _07076_);
  and (_12282_, _07132_, _07076_);
  nor (_12283_, _12282_, _12281_);
  and (_12284_, _06931_, _06016_);
  nor (_12285_, _06931_, _06016_);
  nor (_12286_, _12285_, _12284_);
  and (_12287_, _12286_, _12283_);
  and (_12288_, _12287_, _12280_);
  and (_12289_, _12288_, _12273_);
  or (_12290_, _12289_, _12141_);
  nand (_12291_, _12289_, _12010_);
  and (_12292_, _12291_, _12290_);
  or (_12293_, _12292_, _12255_);
  and (_12294_, _12293_, _12258_);
  and (_12295_, _12294_, _12257_);
  or (_12296_, _12295_, _06121_);
  or (_12297_, _12296_, _12177_);
  not (_12298_, _06115_);
  nor (_12299_, _10988_, _10987_);
  nor (_12300_, _12299_, _10991_);
  not (_12301_, _10994_);
  nor (_12302_, _08127_, \oc8051_golden_model_1.ACC [0]);
  or (_12303_, _12302_, _10995_);
  and (_12304_, _12303_, _12301_);
  and (_12305_, _12304_, _12300_);
  nor (_12306_, _10981_, _10982_);
  nor (_12307_, _12306_, _10986_);
  nor (_12308_, _10980_, _08768_);
  and (_12309_, _12308_, _12307_);
  and (_12310_, _12309_, _12305_);
  and (_12311_, _12310_, _09227_);
  not (_12312_, _12310_);
  and (_12313_, _12312_, _12141_);
  or (_12314_, _12313_, _06509_);
  or (_12315_, _12314_, _12311_);
  and (_12316_, _12315_, _12298_);
  and (_12317_, _12316_, _12297_);
  not (_12318_, _11032_);
  nor (_12319_, _11028_, _11029_);
  nor (_12320_, _12319_, _12318_);
  and (_12321_, _06016_, _05758_);
  nor (_12322_, _12321_, _11036_);
  nor (_12323_, _12322_, _11035_);
  and (_12324_, _12323_, _12320_);
  nor (_12325_, _11021_, _11022_);
  nor (_12326_, _12325_, _11027_);
  nor (_12327_, _11020_, _10705_);
  and (_12328_, _12327_, _12326_);
  and (_12329_, _12328_, _12324_);
  or (_12330_, _12329_, _12141_);
  nand (_12331_, _12329_, _12010_);
  and (_12332_, _12331_, _06115_);
  and (_12333_, _12332_, _12330_);
  or (_12334_, _12333_, _12317_);
  and (_12335_, _12334_, _12013_);
  nand (_12336_, _12012_, _11871_);
  nor (_12337_, _06032_, _07355_);
  and (_12338_, _06222_, _05609_);
  nor (_12339_, _12338_, _06253_);
  and (_12340_, _12339_, _06231_);
  and (_12341_, _06460_, _06221_);
  nor (_12342_, _07248_, _05701_);
  nor (_12343_, _12342_, _12341_);
  and (_12344_, _12343_, _12340_);
  and (_12345_, _12344_, _12337_);
  nand (_12346_, _12345_, _12336_);
  or (_12347_, _12346_, _12335_);
  nor (_12348_, _05701_, _05668_);
  not (_12349_, _12348_);
  nor (_12350_, _11290_, _09269_);
  and (_12351_, _12350_, _12349_);
  or (_12352_, _12345_, _09216_);
  and (_12353_, _12352_, _12351_);
  and (_12354_, _12353_, _12347_);
  not (_12355_, _12351_);
  and (_12356_, _12355_, _11871_);
  and (_12357_, _06252_, _05702_);
  not (_12358_, _12357_);
  or (_12359_, _12358_, _12356_);
  or (_12360_, _12359_, _12354_);
  and (_12361_, _06103_, _05671_);
  nor (_12362_, _10468_, _12361_);
  or (_12363_, _12357_, _09216_);
  and (_12364_, _12363_, _12362_);
  and (_12365_, _12364_, _12360_);
  nor (_12366_, _10306_, _06261_);
  not (_12367_, _12366_);
  not (_12368_, _12362_);
  and (_12369_, _12368_, _11871_);
  or (_12370_, _12369_, _12367_);
  or (_12371_, _12370_, _12365_);
  or (_12372_, _12366_, _09216_);
  and (_12373_, _12372_, _05675_);
  and (_12374_, _12373_, _12371_);
  nand (_12375_, _11871_, _05676_);
  nor (_12376_, _06026_, _06023_);
  nand (_12377_, _12376_, _12375_);
  or (_12378_, _12377_, _12374_);
  or (_12379_, _12376_, _09216_);
  and (_12380_, _12379_, _06111_);
  and (_12381_, _12380_, _12378_);
  nand (_12382_, _09227_, _06110_);
  nand (_12383_, _12382_, _09817_);
  or (_12384_, _12383_, _12381_);
  or (_12385_, _09817_, _09216_);
  and (_12386_, _12385_, _05669_);
  and (_12387_, _12386_, _12384_);
  or (_12388_, _12387_, _12011_);
  nor (_12389_, _09832_, _05663_);
  and (_12390_, _12389_, _12388_);
  nor (_12391_, _06089_, _05719_);
  not (_12392_, _12391_);
  not (_12393_, _12389_);
  and (_12394_, _12393_, _11871_);
  or (_12395_, _12394_, _12392_);
  or (_12396_, _12395_, _12390_);
  and (_12397_, _05659_, _05650_);
  not (_12398_, _12397_);
  or (_12399_, _12391_, _09216_);
  and (_12400_, _12399_, _12398_);
  and (_12401_, _12400_, _12396_);
  and (_12402_, _12397_, _11980_);
  or (_12403_, _12402_, _08743_);
  or (_12404_, _12403_, _12401_);
  and (_12405_, _12404_, _12009_);
  or (_12406_, _12405_, _06019_);
  nand (_12407_, _12010_, _06019_);
  and (_12408_, _12407_, _10662_);
  and (_12409_, _12408_, _12406_);
  and (_12410_, _10661_, _09216_);
  or (_12411_, _12410_, _12409_);
  and (_12412_, _05723_, _06107_);
  not (_12413_, _12412_);
  and (_12414_, _12413_, _12411_);
  nor (_12415_, _06088_, _05724_);
  not (_12416_, _12415_);
  and (_12417_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_12418_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_12419_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_12420_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_12421_, _12420_, _12419_);
  not (_12422_, _12421_);
  and (_12423_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_12424_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_12425_, _12424_, _12423_);
  not (_12426_, _12425_);
  and (_12427_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_12428_, _05862_, _05857_);
  nor (_12429_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_12430_, _12429_, _12427_);
  not (_12431_, _12430_);
  nor (_12432_, _12431_, _12428_);
  nor (_12433_, _12432_, _12427_);
  nor (_12434_, _12433_, _12426_);
  nor (_12435_, _12434_, _12423_);
  nor (_12436_, _12435_, _12422_);
  nor (_12437_, _12436_, _12419_);
  nor (_12438_, _12437_, _12418_);
  or (_12439_, _12438_, _12417_);
  and (_12440_, _12439_, \oc8051_golden_model_1.DPH [0]);
  and (_12441_, _12440_, \oc8051_golden_model_1.DPH [1]);
  and (_12442_, _12441_, \oc8051_golden_model_1.DPH [2]);
  and (_12443_, _12442_, \oc8051_golden_model_1.DPH [3]);
  and (_12444_, _12443_, \oc8051_golden_model_1.DPH [4]);
  and (_12445_, _12444_, \oc8051_golden_model_1.DPH [5]);
  and (_12446_, _12445_, \oc8051_golden_model_1.DPH [6]);
  nand (_12447_, _12446_, \oc8051_golden_model_1.DPH [7]);
  or (_12448_, _12446_, \oc8051_golden_model_1.DPH [7]);
  and (_12449_, _12448_, _12412_);
  and (_12450_, _12449_, _12447_);
  or (_12451_, _12450_, _12416_);
  or (_12452_, _12451_, _12414_);
  and (_12453_, _05723_, _05650_);
  not (_12454_, _12453_);
  or (_12455_, _12415_, _09216_);
  and (_12456_, _12455_, _12454_);
  and (_12457_, _12456_, _12452_);
  or (_12458_, _11980_, _11071_);
  not (_12459_, _11071_);
  or (_12460_, _12459_, _09216_);
  and (_12461_, _12460_, _12453_);
  and (_12462_, _12461_, _12458_);
  or (_12463_, _12462_, _12006_);
  or (_12464_, _12463_, _12457_);
  and (_12465_, _12464_, _12008_);
  nor (_12466_, _10698_, _06282_);
  not (_12467_, _12466_);
  or (_12468_, _12467_, _12465_);
  or (_12469_, _12466_, _09216_);
  and (_12470_, _12469_, _08751_);
  and (_12471_, _12470_, _12468_);
  nand (_12472_, _09227_, _06112_);
  nor (_12473_, _06284_, _05727_);
  nand (_12474_, _12473_, _12472_);
  or (_12475_, _12474_, _12471_);
  and (_12476_, _05726_, _05650_);
  not (_12477_, _12476_);
  or (_12478_, _12473_, _09216_);
  and (_12479_, _12478_, _12477_);
  and (_12480_, _12479_, _12475_);
  not (_12481_, _12002_);
  or (_12482_, _11980_, _12459_);
  or (_12483_, _11071_, _09216_);
  and (_12484_, _12483_, _12476_);
  and (_12485_, _12484_, _12482_);
  or (_12486_, _12485_, _12481_);
  or (_12487_, _12486_, _12480_);
  and (_12488_, _12487_, _12003_);
  or (_12489_, _12488_, _10743_);
  or (_12490_, _10742_, _09216_);
  and (_12491_, _12490_, _07032_);
  and (_12492_, _12491_, _12489_);
  nand (_12493_, _09227_, _06108_);
  nor (_12494_, _06277_, _05736_);
  nand (_12495_, _12494_, _12493_);
  or (_12496_, _12495_, _12492_);
  and (_12497_, _05735_, _05650_);
  not (_12498_, _12497_);
  or (_12499_, _12494_, _09216_);
  and (_12500_, _12499_, _12498_);
  and (_12501_, _12500_, _12496_);
  not (_12502_, _11993_);
  or (_12503_, _11980_, \oc8051_golden_model_1.PSW [7]);
  or (_12504_, _09216_, _10606_);
  and (_12505_, _12504_, _12497_);
  and (_12506_, _12505_, _12503_);
  or (_12507_, _12506_, _12502_);
  or (_12508_, _12507_, _12501_);
  and (_12509_, _12508_, _11994_);
  or (_12510_, _12509_, _11987_);
  or (_12511_, _11986_, _09216_);
  and (_12512_, _12511_, _08777_);
  and (_12513_, _12512_, _12510_);
  nand (_12514_, _09227_, _06130_);
  nor (_12515_, _06292_, _05740_);
  nand (_12516_, _12515_, _12514_);
  or (_12517_, _12516_, _12513_);
  not (_12518_, _11982_);
  or (_12519_, _12515_, _09216_);
  and (_12520_, _12519_, _12518_);
  and (_12521_, _12520_, _12517_);
  or (_12522_, _12521_, _11985_);
  nor (_12523_, _10794_, _10303_);
  and (_12524_, _12523_, _12522_);
  not (_12525_, _12523_);
  and (_12526_, _12525_, _11871_);
  or (_12527_, _12526_, _10826_);
  or (_12528_, _12527_, _12524_);
  or (_12529_, _10825_, _09216_);
  and (_12530_, _12529_, _10855_);
  and (_12531_, _12530_, _12528_);
  and (_12532_, _11871_, _10854_);
  or (_12533_, _12532_, _06298_);
  or (_12534_, _12533_, _12531_);
  nand (_12535_, _07785_, _06298_);
  and (_12536_, _12535_, _12534_);
  or (_12537_, _12536_, _05732_);
  or (_12538_, _09216_, _05734_);
  and (_12539_, _12538_, _06306_);
  and (_12540_, _12539_, _12537_);
  not (_12541_, _11872_);
  not (_12542_, _07732_);
  and (_12543_, _07638_, \oc8051_golden_model_1.P0 [2]);
  and (_12544_, _08341_, \oc8051_golden_model_1.TCON [2]);
  and (_12545_, _08345_, \oc8051_golden_model_1.P1 [2]);
  and (_12546_, _08347_, \oc8051_golden_model_1.SCON [2]);
  and (_12547_, _08349_, \oc8051_golden_model_1.P2 [2]);
  and (_12548_, _08351_, \oc8051_golden_model_1.IE [2]);
  and (_12549_, _08353_, \oc8051_golden_model_1.P3 [2]);
  and (_12550_, _08357_, \oc8051_golden_model_1.IP [2]);
  and (_12551_, _08355_, \oc8051_golden_model_1.PSW [2]);
  and (_12552_, _08359_, \oc8051_golden_model_1.ACC [2]);
  and (_12553_, _08361_, \oc8051_golden_model_1.B [2]);
  or (_12554_, _12553_, _12552_);
  or (_12555_, _12554_, _12551_);
  or (_12556_, _12555_, _12550_);
  or (_12557_, _12556_, _12549_);
  or (_12558_, _12557_, _12548_);
  or (_12559_, _12558_, _12547_);
  or (_12560_, _12559_, _12546_);
  or (_12561_, _12560_, _12545_);
  or (_12562_, _12561_, _12544_);
  nor (_12563_, _12562_, _12543_);
  and (_12564_, _12563_, _08175_);
  nor (_12565_, _12564_, _12542_);
  not (_12566_, _07726_);
  and (_12567_, _08357_, \oc8051_golden_model_1.IP [1]);
  and (_12568_, _08355_, \oc8051_golden_model_1.PSW [1]);
  and (_12569_, _08359_, \oc8051_golden_model_1.ACC [1]);
  and (_12570_, _08361_, \oc8051_golden_model_1.B [1]);
  or (_12571_, _12570_, _12569_);
  or (_12572_, _12571_, _12568_);
  and (_12573_, _08341_, \oc8051_golden_model_1.TCON [1]);
  and (_12574_, _07638_, \oc8051_golden_model_1.P0 [1]);
  and (_12575_, _08345_, \oc8051_golden_model_1.P1 [1]);
  or (_12576_, _12575_, _12574_);
  or (_12577_, _12576_, _12573_);
  and (_12578_, _08353_, \oc8051_golden_model_1.P3 [1]);
  and (_12579_, _08351_, \oc8051_golden_model_1.IE [1]);
  or (_12580_, _12579_, _12578_);
  and (_12581_, _08347_, \oc8051_golden_model_1.SCON [1]);
  and (_12582_, _08349_, \oc8051_golden_model_1.P2 [1]);
  or (_12583_, _12582_, _12581_);
  or (_12584_, _12583_, _12580_);
  or (_12585_, _12584_, _12577_);
  or (_12586_, _12585_, _12572_);
  nor (_12587_, _12586_, _12567_);
  and (_12588_, _12587_, _08076_);
  nor (_12589_, _12588_, _12566_);
  nor (_12590_, _12589_, _12565_);
  and (_12591_, _07644_, _06403_);
  not (_12592_, _12591_);
  and (_12593_, _07638_, \oc8051_golden_model_1.P0 [0]);
  and (_12594_, _08341_, \oc8051_golden_model_1.TCON [0]);
  and (_12595_, _08345_, \oc8051_golden_model_1.P1 [0]);
  and (_12596_, _08347_, \oc8051_golden_model_1.SCON [0]);
  and (_12597_, _08349_, \oc8051_golden_model_1.P2 [0]);
  and (_12598_, _08351_, \oc8051_golden_model_1.IE [0]);
  and (_12599_, _08353_, \oc8051_golden_model_1.P3 [0]);
  and (_12600_, _08357_, \oc8051_golden_model_1.IP [0]);
  and (_12601_, _08355_, \oc8051_golden_model_1.PSW [0]);
  and (_12602_, _08359_, \oc8051_golden_model_1.ACC [0]);
  and (_12603_, _08361_, \oc8051_golden_model_1.B [0]);
  or (_12604_, _12603_, _12602_);
  or (_12605_, _12604_, _12601_);
  or (_12606_, _12605_, _12600_);
  or (_12607_, _12606_, _12599_);
  or (_12608_, _12607_, _12598_);
  or (_12609_, _12608_, _12597_);
  or (_12610_, _12609_, _12596_);
  or (_12611_, _12610_, _12595_);
  or (_12612_, _12611_, _12594_);
  nor (_12613_, _12612_, _12593_);
  not (_12614_, _12613_);
  nor (_12615_, _12614_, _08126_);
  nor (_12616_, _12615_, _12592_);
  and (_12617_, _07638_, \oc8051_golden_model_1.P0 [5]);
  and (_12618_, _08341_, \oc8051_golden_model_1.TCON [5]);
  and (_12619_, _08345_, \oc8051_golden_model_1.P1 [5]);
  and (_12620_, _08347_, \oc8051_golden_model_1.SCON [5]);
  and (_12621_, _08349_, \oc8051_golden_model_1.P2 [5]);
  and (_12622_, _08351_, \oc8051_golden_model_1.IE [5]);
  and (_12623_, _08353_, \oc8051_golden_model_1.P3 [5]);
  and (_12624_, _08357_, \oc8051_golden_model_1.IP [5]);
  and (_12625_, _08355_, \oc8051_golden_model_1.PSW [5]);
  and (_12626_, _08359_, \oc8051_golden_model_1.ACC [5]);
  and (_12627_, _08361_, \oc8051_golden_model_1.B [5]);
  or (_12628_, _12627_, _12626_);
  or (_12629_, _12628_, _12625_);
  or (_12630_, _12629_, _12624_);
  or (_12631_, _12630_, _12623_);
  or (_12632_, _12631_, _12622_);
  or (_12633_, _12632_, _12621_);
  or (_12634_, _12633_, _12620_);
  or (_12635_, _12634_, _12619_);
  or (_12636_, _12635_, _12618_);
  nor (_12637_, _12636_, _12617_);
  and (_12638_, _12637_, _07978_);
  and (_12639_, _07650_, _07477_);
  not (_12640_, _12639_);
  nor (_12641_, _12640_, _12638_);
  nor (_12642_, _12641_, _12616_);
  and (_12643_, _12642_, _12590_);
  not (_12644_, _07723_);
  and (_12645_, _08357_, \oc8051_golden_model_1.IP [3]);
  and (_12646_, _08355_, \oc8051_golden_model_1.PSW [3]);
  and (_12647_, _08361_, \oc8051_golden_model_1.B [3]);
  and (_12648_, _08359_, \oc8051_golden_model_1.ACC [3]);
  or (_12649_, _12648_, _12647_);
  or (_12650_, _12649_, _12646_);
  and (_12651_, _08341_, \oc8051_golden_model_1.TCON [3]);
  and (_12652_, _07638_, \oc8051_golden_model_1.P0 [3]);
  and (_12653_, _08345_, \oc8051_golden_model_1.P1 [3]);
  or (_12654_, _12653_, _12652_);
  or (_12655_, _12654_, _12651_);
  and (_12656_, _08353_, \oc8051_golden_model_1.P3 [3]);
  and (_12657_, _08351_, \oc8051_golden_model_1.IE [3]);
  or (_12658_, _12657_, _12656_);
  and (_12659_, _08347_, \oc8051_golden_model_1.SCON [3]);
  and (_12660_, _08349_, \oc8051_golden_model_1.P2 [3]);
  or (_12661_, _12660_, _12659_);
  or (_12662_, _12661_, _12658_);
  or (_12663_, _12662_, _12655_);
  or (_12664_, _12663_, _12650_);
  nor (_12665_, _12664_, _12645_);
  and (_12666_, _12665_, _08027_);
  nor (_12667_, _12666_, _12644_);
  nor (_12668_, _12667_, _08518_);
  and (_12669_, _07638_, \oc8051_golden_model_1.P0 [6]);
  and (_12670_, _08341_, \oc8051_golden_model_1.TCON [6]);
  and (_12671_, _08345_, \oc8051_golden_model_1.P1 [6]);
  and (_12672_, _08347_, \oc8051_golden_model_1.SCON [6]);
  and (_12673_, _08349_, \oc8051_golden_model_1.P2 [6]);
  and (_12674_, _08351_, \oc8051_golden_model_1.IE [6]);
  and (_12675_, _08353_, \oc8051_golden_model_1.P3 [6]);
  and (_12676_, _08357_, \oc8051_golden_model_1.IP [6]);
  and (_12677_, _08355_, \oc8051_golden_model_1.PSW [6]);
  and (_12678_, _08359_, \oc8051_golden_model_1.ACC [6]);
  and (_12679_, _08361_, \oc8051_golden_model_1.B [6]);
  or (_12680_, _12679_, _12678_);
  or (_12681_, _12680_, _12677_);
  or (_12682_, _12681_, _12676_);
  or (_12683_, _12682_, _12675_);
  or (_12684_, _12683_, _12674_);
  or (_12685_, _12684_, _12673_);
  or (_12686_, _12685_, _12672_);
  or (_12687_, _12686_, _12671_);
  or (_12688_, _12687_, _12670_);
  nor (_12689_, _12688_, _12669_);
  and (_12690_, _12689_, _07884_);
  and (_12691_, _07656_, _07477_);
  not (_12692_, _12691_);
  nor (_12693_, _12692_, _12690_);
  and (_12694_, _08349_, \oc8051_golden_model_1.P2 [4]);
  and (_12695_, _08351_, \oc8051_golden_model_1.IE [4]);
  and (_12696_, _08353_, \oc8051_golden_model_1.P3 [4]);
  or (_12697_, _12696_, _12695_);
  nor (_12698_, _12697_, _12694_);
  and (_12699_, _08341_, \oc8051_golden_model_1.TCON [4]);
  and (_12700_, _08345_, \oc8051_golden_model_1.P1 [4]);
  and (_12701_, _07638_, \oc8051_golden_model_1.P0 [4]);
  or (_12702_, _12701_, _12700_);
  nor (_12703_, _12702_, _12699_);
  and (_12704_, _08357_, \oc8051_golden_model_1.IP [4]);
  and (_12705_, _08361_, \oc8051_golden_model_1.B [4]);
  and (_12706_, _08359_, \oc8051_golden_model_1.ACC [4]);
  or (_12707_, _12706_, _12705_);
  nor (_12708_, _12707_, _12704_);
  and (_12709_, _08347_, \oc8051_golden_model_1.SCON [4]);
  and (_12710_, _08355_, \oc8051_golden_model_1.PSW [4]);
  nor (_12711_, _12710_, _12709_);
  and (_12712_, _12711_, _12708_);
  and (_12714_, _12712_, _12703_);
  and (_12715_, _12714_, _12698_);
  and (_12716_, _12715_, _08271_);
  and (_12717_, _07644_, _07477_);
  not (_12718_, _12717_);
  nor (_12719_, _12718_, _12716_);
  nor (_12720_, _12719_, _12693_);
  and (_12721_, _12720_, _12668_);
  and (_12722_, _12721_, _12643_);
  not (_12723_, _12722_);
  or (_12724_, _12141_, _12723_);
  or (_12725_, _09227_, _12722_);
  and (_12726_, _12725_, _06129_);
  and (_12727_, _12726_, _12724_);
  or (_12728_, _12727_, _12541_);
  or (_12729_, _12728_, _12540_);
  and (_12730_, _12729_, _11873_);
  or (_12731_, _12730_, _10976_);
  or (_12732_, _10975_, _09216_);
  and (_12733_, _12732_, _11016_);
  and (_12735_, _12733_, _12731_);
  and (_12736_, _11871_, _11015_);
  or (_12737_, _12736_, _06049_);
  or (_12738_, _12737_, _12735_);
  nand (_12739_, _07785_, _06049_);
  and (_12740_, _12739_, _12738_);
  or (_12741_, _12740_, _05747_);
  or (_12742_, _09216_, _05748_);
  and (_12743_, _12742_, _06704_);
  and (_12744_, _12743_, _12741_);
  or (_12745_, _12141_, _12722_);
  nand (_12746_, _12010_, _12722_);
  and (_12747_, _12746_, _12745_);
  and (_12748_, _12747_, _06126_);
  and (_12749_, _08287_, _07052_);
  not (_12750_, _12749_);
  or (_12751_, _12750_, _12748_);
  or (_12752_, _12751_, _12744_);
  or (_12753_, _12749_, _11871_);
  and (_12754_, _12753_, _06718_);
  and (_12755_, _12754_, _12752_);
  nor (_12756_, _11064_, _11059_);
  nand (_12757_, _09216_, _06316_);
  nand (_12758_, _12757_, _12756_);
  or (_12759_, _12758_, _12755_);
  or (_12760_, _11871_, _12756_);
  and (_12761_, _12760_, _09200_);
  and (_12762_, _12761_, _12759_);
  and (_12763_, _06127_, _05952_);
  or (_12764_, _12763_, _05752_);
  or (_12765_, _12764_, _12762_);
  not (_12766_, _05752_);
  or (_12767_, _09216_, _12766_);
  and (_12768_, _12767_, _05653_);
  and (_12769_, _12768_, _12765_);
  and (_12770_, _12747_, _05652_);
  and (_12771_, _09154_, _07069_);
  not (_12772_, _12771_);
  or (_12773_, _12772_, _12770_);
  or (_12774_, _12773_, _12769_);
  or (_12775_, _12771_, _11871_);
  and (_12776_, _12775_, _06048_);
  and (_12777_, _12776_, _12774_);
  nand (_12778_, _09216_, _06047_);
  nor (_12779_, _11089_, _11082_);
  nand (_12780_, _12779_, _12778_);
  or (_12781_, _12780_, _12777_);
  not (_12782_, _06119_);
  or (_12783_, _12779_, _11871_);
  and (_12784_, _12783_, _12782_);
  and (_12785_, _12784_, _12781_);
  and (_12786_, _06119_, _05952_);
  or (_12787_, _12786_, _05751_);
  or (_12788_, _12787_, _12785_);
  and (_12789_, _05750_, _05650_);
  not (_12790_, _12789_);
  not (_12791_, _05751_);
  or (_12792_, _09216_, _12791_);
  and (_12793_, _12792_, _12790_);
  and (_12794_, _12793_, _12788_);
  and (_12795_, _12789_, _11871_);
  or (_12796_, _12795_, _12794_);
  or (_12797_, _12796_, _01340_);
  or (_12798_, _01336_, \oc8051_golden_model_1.PC [15]);
  and (_12799_, _12798_, _42882_);
  and (_40766_, _12799_, _12797_);
  not (_12800_, _07686_);
  and (_12801_, _12800_, \oc8051_golden_model_1.P2 [7]);
  and (_12802_, _08768_, _07686_);
  or (_12803_, _12802_, _12801_);
  and (_12804_, _12803_, _06284_);
  and (_12805_, _08549_, _07686_);
  or (_12806_, _12805_, _12801_);
  or (_12807_, _12806_, _06020_);
  and (_12808_, _08498_, _07686_);
  or (_12809_, _12808_, _12801_);
  or (_12810_, _12809_, _06954_);
  and (_12811_, _07686_, \oc8051_golden_model_1.ACC [7]);
  or (_12812_, _12811_, _12801_);
  and (_12813_, _12812_, _06938_);
  and (_12814_, _06939_, \oc8051_golden_model_1.P2 [7]);
  or (_12815_, _12814_, _06102_);
  or (_12816_, _12815_, _12813_);
  and (_12817_, _12816_, _06044_);
  and (_12818_, _12817_, _12810_);
  not (_12819_, _08349_);
  and (_12820_, _12819_, \oc8051_golden_model_1.P2 [7]);
  and (_12821_, _08503_, _08349_);
  or (_12822_, _12821_, _12820_);
  and (_12823_, _12822_, _06043_);
  or (_12824_, _12823_, _06239_);
  or (_12825_, _12824_, _12818_);
  nor (_12826_, _07785_, _12800_);
  or (_12827_, _12826_, _12801_);
  or (_12828_, _12827_, _06848_);
  and (_12829_, _12828_, _12825_);
  or (_12830_, _12829_, _06219_);
  or (_12831_, _12812_, _06220_);
  and (_12832_, _12831_, _06040_);
  and (_12833_, _12832_, _12830_);
  and (_12834_, _08374_, _08349_);
  or (_12835_, _12834_, _12820_);
  and (_12836_, _12835_, _06039_);
  or (_12837_, _12836_, _06032_);
  or (_12838_, _12837_, _12833_);
  or (_12839_, _12820_, _08519_);
  and (_12840_, _12839_, _12822_);
  or (_12841_, _12840_, _06033_);
  and (_12842_, _12841_, _06027_);
  and (_12843_, _12842_, _12838_);
  and (_12844_, _08376_, _08349_);
  or (_12845_, _12844_, _12820_);
  and (_12846_, _12845_, _06026_);
  or (_12847_, _12846_, _09818_);
  or (_12848_, _12847_, _12843_);
  and (_12849_, _08485_, _07686_);
  or (_12850_, _12801_, _07012_);
  or (_12851_, _12850_, _12849_);
  or (_12852_, _12827_, _09827_);
  and (_12853_, _12852_, _05669_);
  and (_12854_, _12853_, _12851_);
  and (_12855_, _12854_, _12848_);
  and (_12856_, _08738_, _07686_);
  or (_12857_, _12856_, _12801_);
  and (_12858_, _12857_, _09833_);
  or (_12859_, _12858_, _06019_);
  or (_12860_, _12859_, _12855_);
  and (_12861_, _12860_, _12807_);
  or (_12862_, _12861_, _06112_);
  and (_12863_, _08760_, _07686_);
  or (_12864_, _12801_, _08751_);
  or (_12865_, _12864_, _12863_);
  and (_12866_, _12865_, _08756_);
  and (_12867_, _12866_, _12862_);
  or (_12868_, _12867_, _12804_);
  and (_12869_, _12868_, _07032_);
  or (_12870_, _12801_, _07788_);
  and (_12871_, _12806_, _06108_);
  and (_12872_, _12871_, _12870_);
  or (_12873_, _12872_, _12869_);
  and (_12874_, _12873_, _06278_);
  and (_12875_, _12812_, _06277_);
  and (_12876_, _12875_, _12870_);
  or (_12877_, _12876_, _06130_);
  or (_12878_, _12877_, _12874_);
  and (_12879_, _08759_, _07686_);
  or (_12880_, _12801_, _08777_);
  or (_12881_, _12880_, _12879_);
  and (_12882_, _12881_, _08782_);
  and (_12883_, _12882_, _12878_);
  nor (_12884_, _08767_, _12800_);
  or (_12885_, _12884_, _12801_);
  and (_12886_, _12885_, _06292_);
  or (_12887_, _12886_, _06316_);
  or (_12888_, _12887_, _12883_);
  or (_12889_, _12809_, _06718_);
  and (_12890_, _12889_, _05653_);
  and (_12891_, _12890_, _12888_);
  and (_12892_, _12835_, _05652_);
  or (_12893_, _12892_, _06047_);
  or (_12894_, _12893_, _12891_);
  and (_12895_, _08279_, _07686_);
  or (_12896_, _12801_, _06048_);
  or (_12897_, _12896_, _12895_);
  and (_12898_, _12897_, _01336_);
  and (_12899_, _12898_, _12894_);
  nor (_12900_, \oc8051_golden_model_1.P2 [7], rst);
  nor (_12901_, _12900_, _00000_);
  or (_40768_, _12901_, _12899_);
  not (_12902_, _07692_);
  and (_12903_, _12902_, \oc8051_golden_model_1.P3 [7]);
  and (_12904_, _08768_, _07692_);
  or (_12905_, _12904_, _12903_);
  and (_12906_, _12905_, _06284_);
  and (_12907_, _08549_, _07692_);
  or (_12908_, _12907_, _12903_);
  or (_12909_, _12908_, _06020_);
  and (_12910_, _08498_, _07692_);
  or (_12911_, _12910_, _12903_);
  or (_12912_, _12911_, _06954_);
  and (_12913_, _07692_, \oc8051_golden_model_1.ACC [7]);
  or (_12914_, _12913_, _12903_);
  and (_12915_, _12914_, _06938_);
  and (_12916_, _06939_, \oc8051_golden_model_1.P3 [7]);
  or (_12917_, _12916_, _06102_);
  or (_12918_, _12917_, _12915_);
  and (_12919_, _12918_, _06044_);
  and (_12920_, _12919_, _12912_);
  not (_12921_, _08353_);
  and (_12922_, _12921_, \oc8051_golden_model_1.P3 [7]);
  and (_12923_, _08503_, _08353_);
  or (_12924_, _12923_, _12922_);
  and (_12925_, _12924_, _06043_);
  or (_12926_, _12925_, _06239_);
  or (_12927_, _12926_, _12920_);
  nor (_12928_, _07785_, _12902_);
  or (_12929_, _12928_, _12903_);
  or (_12930_, _12929_, _06848_);
  and (_12931_, _12930_, _12927_);
  or (_12932_, _12931_, _06219_);
  or (_12933_, _12914_, _06220_);
  and (_12934_, _12933_, _06040_);
  and (_12935_, _12934_, _12932_);
  and (_12936_, _08374_, _08353_);
  or (_12937_, _12936_, _12922_);
  and (_12938_, _12937_, _06039_);
  or (_12939_, _12938_, _06032_);
  or (_12940_, _12939_, _12935_);
  or (_12941_, _12922_, _08519_);
  and (_12942_, _12941_, _12924_);
  or (_12943_, _12942_, _06033_);
  and (_12944_, _12943_, _06027_);
  and (_12945_, _12944_, _12940_);
  and (_12946_, _08376_, _08353_);
  or (_12947_, _12946_, _12922_);
  and (_12948_, _12947_, _06026_);
  or (_12949_, _12948_, _09818_);
  or (_12950_, _12949_, _12945_);
  and (_12951_, _08485_, _07692_);
  or (_12952_, _12903_, _07012_);
  or (_12953_, _12952_, _12951_);
  or (_12954_, _12929_, _09827_);
  and (_12955_, _12954_, _05669_);
  and (_12956_, _12955_, _12953_);
  and (_12957_, _12956_, _12950_);
  and (_12958_, _08738_, _07692_);
  or (_12959_, _12958_, _12903_);
  and (_12960_, _12959_, _09833_);
  or (_12961_, _12960_, _06019_);
  or (_12962_, _12961_, _12957_);
  and (_12963_, _12962_, _12909_);
  or (_12964_, _12963_, _06112_);
  and (_12965_, _08760_, _07692_);
  or (_12966_, _12965_, _12903_);
  or (_12967_, _12966_, _08751_);
  and (_12968_, _12967_, _08756_);
  and (_12969_, _12968_, _12964_);
  or (_12970_, _12969_, _12906_);
  and (_12971_, _12970_, _07032_);
  or (_12972_, _12903_, _07788_);
  and (_12973_, _12908_, _06108_);
  and (_12974_, _12973_, _12972_);
  or (_12975_, _12974_, _12971_);
  and (_12976_, _12975_, _06278_);
  and (_12977_, _12914_, _06277_);
  and (_12978_, _12977_, _12972_);
  or (_12979_, _12978_, _06130_);
  or (_12980_, _12979_, _12976_);
  and (_12981_, _08759_, _07692_);
  or (_12982_, _12903_, _08777_);
  or (_12983_, _12982_, _12981_);
  and (_12984_, _12983_, _08782_);
  and (_12985_, _12984_, _12980_);
  nor (_12986_, _08767_, _12902_);
  or (_12987_, _12986_, _12903_);
  and (_12988_, _12987_, _06292_);
  or (_12989_, _12988_, _06316_);
  or (_12990_, _12989_, _12985_);
  or (_12991_, _12911_, _06718_);
  and (_12992_, _12991_, _05653_);
  and (_12993_, _12992_, _12990_);
  and (_12994_, _12937_, _05652_);
  or (_12995_, _12994_, _06047_);
  or (_12996_, _12995_, _12993_);
  and (_12997_, _08279_, _07692_);
  or (_12998_, _12903_, _06048_);
  or (_12999_, _12998_, _12997_);
  and (_13000_, _12999_, _01336_);
  and (_13001_, _13000_, _12996_);
  nor (_13002_, \oc8051_golden_model_1.P3 [7], rst);
  nor (_13003_, _13002_, _00000_);
  or (_40769_, _13003_, _13001_);
  nor (_13004_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_13005_, _13004_, _00000_);
  not (_13006_, _07730_);
  and (_13007_, _13006_, \oc8051_golden_model_1.P0 [7]);
  and (_13008_, _08768_, _07730_);
  or (_13009_, _13008_, _13007_);
  and (_13010_, _13009_, _06284_);
  and (_13011_, _08549_, _07730_);
  or (_13012_, _13011_, _13007_);
  or (_13013_, _13012_, _06020_);
  and (_13014_, _08498_, _07730_);
  or (_13015_, _13014_, _13007_);
  or (_13016_, _13015_, _06954_);
  and (_13017_, _07730_, \oc8051_golden_model_1.ACC [7]);
  or (_13018_, _13017_, _13007_);
  and (_13019_, _13018_, _06938_);
  and (_13020_, _06939_, \oc8051_golden_model_1.P0 [7]);
  or (_13021_, _13020_, _06102_);
  or (_13022_, _13021_, _13019_);
  and (_13023_, _13022_, _06044_);
  and (_13024_, _13023_, _13016_);
  not (_13025_, _07638_);
  and (_13026_, _13025_, \oc8051_golden_model_1.P0 [7]);
  and (_13027_, _08503_, _07638_);
  or (_13028_, _13027_, _13026_);
  and (_13029_, _13028_, _06043_);
  or (_13030_, _13029_, _06239_);
  or (_13031_, _13030_, _13024_);
  nor (_13032_, _07785_, _13006_);
  or (_13033_, _13032_, _13007_);
  or (_13034_, _13033_, _06848_);
  and (_13035_, _13034_, _13031_);
  or (_13036_, _13035_, _06219_);
  or (_13037_, _13018_, _06220_);
  and (_13038_, _13037_, _06040_);
  and (_13039_, _13038_, _13036_);
  and (_13040_, _08374_, _07638_);
  or (_13041_, _13040_, _13026_);
  and (_13042_, _13041_, _06039_);
  or (_13043_, _13042_, _06032_);
  or (_13044_, _13043_, _13039_);
  or (_13045_, _13026_, _08519_);
  and (_13046_, _13045_, _13028_);
  or (_13047_, _13046_, _06033_);
  and (_13048_, _13047_, _06027_);
  and (_13049_, _13048_, _13044_);
  and (_13050_, _08376_, _07638_);
  or (_13051_, _13050_, _13026_);
  and (_13052_, _13051_, _06026_);
  or (_13053_, _13052_, _09818_);
  or (_13054_, _13053_, _13049_);
  and (_13055_, _08485_, _07730_);
  or (_13056_, _13007_, _07012_);
  or (_13057_, _13056_, _13055_);
  or (_13058_, _13033_, _09827_);
  and (_13059_, _13058_, _05669_);
  and (_13060_, _13059_, _13057_);
  and (_13061_, _13060_, _13054_);
  and (_13062_, _08738_, _07730_);
  or (_13063_, _13062_, _13007_);
  and (_13064_, _13063_, _09833_);
  or (_13065_, _13064_, _06019_);
  or (_13066_, _13065_, _13061_);
  and (_13067_, _13066_, _13013_);
  or (_13068_, _13067_, _06112_);
  and (_13069_, _08760_, _07730_);
  or (_13070_, _13007_, _08751_);
  or (_13071_, _13070_, _13069_);
  and (_13072_, _13071_, _08756_);
  and (_13073_, _13072_, _13068_);
  or (_13074_, _13073_, _13010_);
  and (_13075_, _13074_, _07032_);
  or (_13076_, _13007_, _07788_);
  and (_13077_, _13012_, _06108_);
  and (_13078_, _13077_, _13076_);
  or (_13079_, _13078_, _13075_);
  and (_13080_, _13079_, _06278_);
  and (_13081_, _13018_, _06277_);
  and (_13082_, _13081_, _13076_);
  or (_13083_, _13082_, _06130_);
  or (_13084_, _13083_, _13080_);
  and (_13085_, _08759_, _07730_);
  or (_13086_, _13007_, _08777_);
  or (_13087_, _13086_, _13085_);
  and (_13088_, _13087_, _08782_);
  and (_13089_, _13088_, _13084_);
  nor (_13090_, _08767_, _13006_);
  or (_13091_, _13090_, _13007_);
  and (_13092_, _13091_, _06292_);
  or (_13093_, _13092_, _06316_);
  or (_13094_, _13093_, _13089_);
  or (_13095_, _13015_, _06718_);
  and (_13096_, _13095_, _05653_);
  and (_13097_, _13096_, _13094_);
  and (_13098_, _13041_, _05652_);
  or (_13099_, _13098_, _06047_);
  or (_13100_, _13099_, _13097_);
  and (_13101_, _08279_, _07730_);
  or (_13102_, _13007_, _06048_);
  or (_13103_, _13102_, _13101_);
  and (_13104_, _13103_, _01336_);
  and (_13105_, _13104_, _13100_);
  or (_40770_, _13105_, _13005_);
  nor (_13106_, \oc8051_golden_model_1.P1 [7], rst);
  nor (_13107_, _13106_, _00000_);
  not (_13108_, _07677_);
  and (_13109_, _13108_, \oc8051_golden_model_1.P1 [7]);
  and (_13110_, _08768_, _07677_);
  or (_13111_, _13110_, _13109_);
  and (_13112_, _13111_, _06284_);
  and (_13113_, _08549_, _07677_);
  or (_13114_, _13113_, _13109_);
  or (_13115_, _13114_, _06020_);
  and (_13116_, _08498_, _07677_);
  or (_13117_, _13116_, _13109_);
  or (_13118_, _13117_, _06954_);
  and (_13119_, _07677_, \oc8051_golden_model_1.ACC [7]);
  or (_13120_, _13119_, _13109_);
  and (_13121_, _13120_, _06938_);
  and (_13122_, _06939_, \oc8051_golden_model_1.P1 [7]);
  or (_13123_, _13122_, _06102_);
  or (_13124_, _13123_, _13121_);
  and (_13125_, _13124_, _06044_);
  and (_13126_, _13125_, _13118_);
  not (_13127_, _08345_);
  and (_13128_, _13127_, \oc8051_golden_model_1.P1 [7]);
  and (_13129_, _08503_, _08345_);
  or (_13130_, _13129_, _13128_);
  and (_13131_, _13130_, _06043_);
  or (_13132_, _13131_, _06239_);
  or (_13133_, _13132_, _13126_);
  nor (_13134_, _07785_, _13108_);
  or (_13135_, _13134_, _13109_);
  or (_13136_, _13135_, _06848_);
  and (_13137_, _13136_, _13133_);
  or (_13138_, _13137_, _06219_);
  or (_13139_, _13120_, _06220_);
  and (_13140_, _13139_, _06040_);
  and (_13141_, _13140_, _13138_);
  and (_13142_, _08374_, _08345_);
  or (_13143_, _13142_, _13128_);
  and (_13144_, _13143_, _06039_);
  or (_13145_, _13144_, _06032_);
  or (_13146_, _13145_, _13141_);
  or (_13147_, _13128_, _08519_);
  and (_13148_, _13147_, _13130_);
  or (_13149_, _13148_, _06033_);
  and (_13150_, _13149_, _06027_);
  and (_13151_, _13150_, _13146_);
  and (_13152_, _08376_, _08345_);
  or (_13153_, _13152_, _13128_);
  and (_13154_, _13153_, _06026_);
  or (_13155_, _13154_, _09818_);
  or (_13156_, _13155_, _13151_);
  and (_13157_, _08485_, _07677_);
  or (_13158_, _13109_, _07012_);
  or (_13159_, _13158_, _13157_);
  or (_13160_, _13135_, _09827_);
  and (_13161_, _13160_, _05669_);
  and (_13162_, _13161_, _13159_);
  and (_13163_, _13162_, _13156_);
  and (_13164_, _08738_, _07677_);
  or (_13165_, _13164_, _13109_);
  and (_13166_, _13165_, _09833_);
  or (_13167_, _13166_, _06019_);
  or (_13168_, _13167_, _13163_);
  and (_13169_, _13168_, _13115_);
  or (_13170_, _13169_, _06112_);
  and (_13171_, _08760_, _07677_);
  or (_13172_, _13171_, _13109_);
  or (_13173_, _13172_, _08751_);
  and (_13174_, _13173_, _08756_);
  and (_13175_, _13174_, _13170_);
  or (_13176_, _13175_, _13112_);
  and (_13177_, _13176_, _07032_);
  or (_13178_, _13109_, _07788_);
  and (_13179_, _13114_, _06108_);
  and (_13180_, _13179_, _13178_);
  or (_13181_, _13180_, _13177_);
  and (_13182_, _13181_, _06278_);
  and (_13183_, _13120_, _06277_);
  and (_13184_, _13183_, _13178_);
  or (_13185_, _13184_, _06130_);
  or (_13186_, _13185_, _13182_);
  and (_13187_, _08759_, _07677_);
  or (_13188_, _13109_, _08777_);
  or (_13189_, _13188_, _13187_);
  and (_13190_, _13189_, _08782_);
  and (_13191_, _13190_, _13186_);
  nor (_13192_, _08767_, _13108_);
  or (_13193_, _13192_, _13109_);
  and (_13194_, _13193_, _06292_);
  or (_13195_, _13194_, _06316_);
  or (_13196_, _13195_, _13191_);
  or (_13197_, _13117_, _06718_);
  and (_13198_, _13197_, _05653_);
  and (_13199_, _13198_, _13196_);
  and (_13200_, _13143_, _05652_);
  or (_13201_, _13200_, _06047_);
  or (_13202_, _13201_, _13199_);
  and (_13203_, _08279_, _07677_);
  or (_13204_, _13109_, _06048_);
  or (_13205_, _13204_, _13203_);
  and (_13206_, _13205_, _01336_);
  and (_13207_, _13206_, _13202_);
  or (_40771_, _13207_, _13107_);
  and (_13208_, _01340_, \oc8051_golden_model_1.IP [7]);
  not (_13209_, _07694_);
  and (_13210_, _13209_, \oc8051_golden_model_1.IP [7]);
  and (_13211_, _08768_, _07694_);
  or (_13212_, _13211_, _13210_);
  and (_13213_, _13212_, _06284_);
  and (_13214_, _08549_, _07694_);
  or (_13215_, _13214_, _13210_);
  or (_13216_, _13215_, _06020_);
  and (_13217_, _08498_, _07694_);
  or (_13218_, _13217_, _13210_);
  or (_13219_, _13218_, _06954_);
  and (_13220_, _07694_, \oc8051_golden_model_1.ACC [7]);
  or (_13221_, _13220_, _13210_);
  and (_13222_, _13221_, _06938_);
  and (_13223_, _06939_, \oc8051_golden_model_1.IP [7]);
  or (_13224_, _13223_, _06102_);
  or (_13225_, _13224_, _13222_);
  and (_13226_, _13225_, _06044_);
  and (_13227_, _13226_, _13219_);
  not (_13228_, _08357_);
  and (_13229_, _13228_, \oc8051_golden_model_1.IP [7]);
  and (_13230_, _08503_, _08357_);
  or (_13231_, _13230_, _13229_);
  and (_13232_, _13231_, _06043_);
  or (_13233_, _13232_, _06239_);
  or (_13234_, _13233_, _13227_);
  nor (_13235_, _07785_, _13209_);
  or (_13236_, _13235_, _13210_);
  or (_13237_, _13236_, _06848_);
  and (_13238_, _13237_, _13234_);
  or (_13239_, _13238_, _06219_);
  or (_13240_, _13221_, _06220_);
  and (_13241_, _13240_, _06040_);
  and (_13242_, _13241_, _13239_);
  and (_13243_, _08374_, _08357_);
  or (_13244_, _13243_, _13229_);
  and (_13245_, _13244_, _06039_);
  or (_13246_, _13245_, _06032_);
  or (_13247_, _13246_, _13242_);
  or (_13248_, _13229_, _08519_);
  and (_13249_, _13248_, _13231_);
  or (_13250_, _13249_, _06033_);
  and (_13251_, _13250_, _06027_);
  and (_13252_, _13251_, _13247_);
  and (_13253_, _08376_, _08357_);
  or (_13254_, _13253_, _13229_);
  and (_13255_, _13254_, _06026_);
  or (_13256_, _13255_, _09818_);
  or (_13257_, _13256_, _13252_);
  and (_13258_, _08485_, _07694_);
  or (_13259_, _13210_, _07012_);
  or (_13260_, _13259_, _13258_);
  or (_13261_, _13236_, _09827_);
  and (_13262_, _13261_, _05669_);
  and (_13263_, _13262_, _13260_);
  and (_13264_, _13263_, _13257_);
  and (_13265_, _08738_, _07694_);
  or (_13266_, _13265_, _13210_);
  and (_13267_, _13266_, _09833_);
  or (_13268_, _13267_, _06019_);
  or (_13269_, _13268_, _13264_);
  and (_13270_, _13269_, _13216_);
  or (_13271_, _13270_, _06112_);
  and (_13272_, _08760_, _07694_);
  or (_13273_, _13210_, _08751_);
  or (_13274_, _13273_, _13272_);
  and (_13275_, _13274_, _08756_);
  and (_13276_, _13275_, _13271_);
  or (_13277_, _13276_, _13213_);
  and (_13278_, _13277_, _07032_);
  or (_13279_, _13210_, _07788_);
  and (_13280_, _13215_, _06108_);
  and (_13281_, _13280_, _13279_);
  or (_13282_, _13281_, _13278_);
  and (_13283_, _13282_, _06278_);
  and (_13284_, _13221_, _06277_);
  and (_13285_, _13284_, _13279_);
  or (_13286_, _13285_, _06130_);
  or (_13287_, _13286_, _13283_);
  and (_13288_, _08759_, _07694_);
  or (_13289_, _13210_, _08777_);
  or (_13290_, _13289_, _13288_);
  and (_13291_, _13290_, _08782_);
  and (_13292_, _13291_, _13287_);
  nor (_13293_, _08767_, _13209_);
  or (_13294_, _13293_, _13210_);
  and (_13295_, _13294_, _06292_);
  or (_13296_, _13295_, _06316_);
  or (_13297_, _13296_, _13292_);
  or (_13298_, _13218_, _06718_);
  and (_13299_, _13298_, _05653_);
  and (_13300_, _13299_, _13297_);
  and (_13301_, _13244_, _05652_);
  or (_13302_, _13301_, _06047_);
  or (_13303_, _13302_, _13300_);
  and (_13304_, _08279_, _07694_);
  or (_13305_, _13210_, _06048_);
  or (_13306_, _13305_, _13304_);
  and (_13307_, _13306_, _01336_);
  and (_13308_, _13307_, _13303_);
  or (_13309_, _13308_, _13208_);
  and (_40772_, _13309_, _42882_);
  and (_13310_, _01340_, \oc8051_golden_model_1.IE [7]);
  not (_13311_, _07688_);
  and (_13312_, _13311_, \oc8051_golden_model_1.IE [7]);
  and (_13313_, _08768_, _07688_);
  or (_13314_, _13313_, _13312_);
  and (_13315_, _13314_, _06284_);
  and (_13316_, _08549_, _07688_);
  or (_13317_, _13316_, _13312_);
  or (_13318_, _13317_, _06020_);
  and (_13319_, _08498_, _07688_);
  or (_13320_, _13319_, _13312_);
  or (_13321_, _13320_, _06954_);
  and (_13322_, _07688_, \oc8051_golden_model_1.ACC [7]);
  or (_13323_, _13322_, _13312_);
  and (_13324_, _13323_, _06938_);
  and (_13325_, _06939_, \oc8051_golden_model_1.IE [7]);
  or (_13326_, _13325_, _06102_);
  or (_13327_, _13326_, _13324_);
  and (_13328_, _13327_, _06044_);
  and (_13329_, _13328_, _13321_);
  not (_13330_, _08351_);
  and (_13331_, _13330_, \oc8051_golden_model_1.IE [7]);
  and (_13332_, _08503_, _08351_);
  or (_13333_, _13332_, _13331_);
  and (_13334_, _13333_, _06043_);
  or (_13335_, _13334_, _06239_);
  or (_13336_, _13335_, _13329_);
  nor (_13337_, _07785_, _13311_);
  or (_13338_, _13337_, _13312_);
  or (_13339_, _13338_, _06848_);
  and (_13340_, _13339_, _13336_);
  or (_13341_, _13340_, _06219_);
  or (_13342_, _13323_, _06220_);
  and (_13343_, _13342_, _06040_);
  and (_13344_, _13343_, _13341_);
  and (_13345_, _08374_, _08351_);
  or (_13346_, _13345_, _13331_);
  and (_13347_, _13346_, _06039_);
  or (_13348_, _13347_, _06032_);
  or (_13349_, _13348_, _13344_);
  or (_13350_, _13331_, _08519_);
  and (_13351_, _13350_, _13333_);
  or (_13352_, _13351_, _06033_);
  and (_13353_, _13352_, _06027_);
  and (_13354_, _13353_, _13349_);
  and (_13355_, _08376_, _08351_);
  or (_13356_, _13355_, _13331_);
  and (_13357_, _13356_, _06026_);
  or (_13358_, _13357_, _09818_);
  or (_13359_, _13358_, _13354_);
  and (_13360_, _08485_, _07688_);
  or (_13361_, _13312_, _07012_);
  or (_13362_, _13361_, _13360_);
  or (_13363_, _13338_, _09827_);
  and (_13364_, _13363_, _05669_);
  and (_13365_, _13364_, _13362_);
  and (_13366_, _13365_, _13359_);
  and (_13367_, _08738_, _07688_);
  or (_13368_, _13367_, _13312_);
  and (_13369_, _13368_, _09833_);
  or (_13370_, _13369_, _06019_);
  or (_13371_, _13370_, _13366_);
  and (_13372_, _13371_, _13318_);
  or (_13373_, _13372_, _06112_);
  and (_13374_, _08760_, _07688_);
  or (_13375_, _13374_, _13312_);
  or (_13376_, _13375_, _08751_);
  and (_13377_, _13376_, _08756_);
  and (_13378_, _13377_, _13373_);
  or (_13379_, _13378_, _13315_);
  and (_13380_, _13379_, _07032_);
  or (_13381_, _13312_, _07788_);
  and (_13382_, _13317_, _06108_);
  and (_13383_, _13382_, _13381_);
  or (_13384_, _13383_, _13380_);
  and (_13385_, _13384_, _06278_);
  and (_13386_, _13323_, _06277_);
  and (_13387_, _13386_, _13381_);
  or (_13388_, _13387_, _06130_);
  or (_13389_, _13388_, _13385_);
  and (_13390_, _08759_, _07688_);
  or (_13391_, _13312_, _08777_);
  or (_13392_, _13391_, _13390_);
  and (_13393_, _13392_, _08782_);
  and (_13394_, _13393_, _13389_);
  nor (_13395_, _08767_, _13311_);
  or (_13396_, _13395_, _13312_);
  and (_13397_, _13396_, _06292_);
  or (_13398_, _13397_, _06316_);
  or (_13399_, _13398_, _13394_);
  or (_13400_, _13320_, _06718_);
  and (_13401_, _13400_, _05653_);
  and (_13402_, _13401_, _13399_);
  and (_13403_, _13346_, _05652_);
  or (_13404_, _13403_, _06047_);
  or (_13405_, _13404_, _13402_);
  and (_13406_, _08279_, _07688_);
  or (_13407_, _13312_, _06048_);
  or (_13408_, _13407_, _13406_);
  and (_13409_, _13408_, _01336_);
  and (_13410_, _13409_, _13405_);
  or (_13411_, _13410_, _13310_);
  and (_40774_, _13411_, _42882_);
  and (_13412_, _01340_, \oc8051_golden_model_1.SCON [7]);
  not (_13413_, _07679_);
  and (_13414_, _13413_, \oc8051_golden_model_1.SCON [7]);
  and (_13415_, _08768_, _07679_);
  or (_13416_, _13415_, _13414_);
  and (_13417_, _13416_, _06284_);
  and (_13418_, _08549_, _07679_);
  or (_13419_, _13418_, _13414_);
  or (_13420_, _13419_, _06020_);
  and (_13421_, _08498_, _07679_);
  or (_13422_, _13421_, _13414_);
  or (_13423_, _13422_, _06954_);
  and (_13424_, _07679_, \oc8051_golden_model_1.ACC [7]);
  or (_13425_, _13424_, _13414_);
  and (_13426_, _13425_, _06938_);
  and (_13427_, _06939_, \oc8051_golden_model_1.SCON [7]);
  or (_13428_, _13427_, _06102_);
  or (_13429_, _13428_, _13426_);
  and (_13430_, _13429_, _06044_);
  and (_13431_, _13430_, _13423_);
  not (_13432_, _08347_);
  and (_13433_, _13432_, \oc8051_golden_model_1.SCON [7]);
  and (_13434_, _08503_, _08347_);
  or (_13435_, _13434_, _13433_);
  and (_13436_, _13435_, _06043_);
  or (_13437_, _13436_, _06239_);
  or (_13438_, _13437_, _13431_);
  nor (_13439_, _07785_, _13413_);
  or (_13440_, _13439_, _13414_);
  or (_13441_, _13440_, _06848_);
  and (_13442_, _13441_, _13438_);
  or (_13443_, _13442_, _06219_);
  or (_13444_, _13425_, _06220_);
  and (_13445_, _13444_, _06040_);
  and (_13446_, _13445_, _13443_);
  and (_13447_, _08374_, _08347_);
  or (_13448_, _13447_, _13433_);
  and (_13449_, _13448_, _06039_);
  or (_13450_, _13449_, _06032_);
  or (_13451_, _13450_, _13446_);
  or (_13452_, _13433_, _08519_);
  and (_13453_, _13452_, _13435_);
  or (_13454_, _13453_, _06033_);
  and (_13455_, _13454_, _06027_);
  and (_13456_, _13455_, _13451_);
  and (_13457_, _08376_, _08347_);
  or (_13458_, _13457_, _13433_);
  and (_13459_, _13458_, _06026_);
  or (_13460_, _13459_, _09818_);
  or (_13461_, _13460_, _13456_);
  and (_13462_, _08485_, _07679_);
  or (_13463_, _13414_, _07012_);
  or (_13464_, _13463_, _13462_);
  or (_13465_, _13440_, _09827_);
  and (_13466_, _13465_, _05669_);
  and (_13467_, _13466_, _13464_);
  and (_13468_, _13467_, _13461_);
  and (_13469_, _08738_, _07679_);
  or (_13470_, _13469_, _13414_);
  and (_13471_, _13470_, _09833_);
  or (_13472_, _13471_, _06019_);
  or (_13473_, _13472_, _13468_);
  and (_13474_, _13473_, _13420_);
  or (_13475_, _13474_, _06112_);
  and (_13476_, _08760_, _07679_);
  or (_13477_, _13476_, _13414_);
  or (_13478_, _13477_, _08751_);
  and (_13479_, _13478_, _08756_);
  and (_13480_, _13479_, _13475_);
  or (_13481_, _13480_, _13417_);
  and (_13482_, _13481_, _07032_);
  or (_13483_, _13414_, _07788_);
  and (_13484_, _13419_, _06108_);
  and (_13485_, _13484_, _13483_);
  or (_13486_, _13485_, _13482_);
  and (_13487_, _13486_, _06278_);
  and (_13488_, _13425_, _06277_);
  and (_13489_, _13488_, _13483_);
  or (_13490_, _13489_, _06130_);
  or (_13491_, _13490_, _13487_);
  and (_13492_, _08759_, _07679_);
  or (_13493_, _13414_, _08777_);
  or (_13494_, _13493_, _13492_);
  and (_13495_, _13494_, _08782_);
  and (_13496_, _13495_, _13491_);
  nor (_13497_, _08767_, _13413_);
  or (_13498_, _13497_, _13414_);
  and (_13499_, _13498_, _06292_);
  or (_13500_, _13499_, _06316_);
  or (_13501_, _13500_, _13496_);
  or (_13502_, _13422_, _06718_);
  and (_13503_, _13502_, _05653_);
  and (_13504_, _13503_, _13501_);
  and (_13505_, _13448_, _05652_);
  or (_13506_, _13505_, _06047_);
  or (_13507_, _13506_, _13504_);
  and (_13508_, _08279_, _07679_);
  or (_13509_, _13414_, _06048_);
  or (_13510_, _13509_, _13508_);
  and (_13511_, _13510_, _01336_);
  and (_13512_, _13511_, _13507_);
  or (_13513_, _13512_, _13412_);
  and (_40775_, _13513_, _42882_);
  not (_13514_, \oc8051_golden_model_1.SP [7]);
  nor (_13515_, _01336_, _13514_);
  and (_13516_, _07360_, \oc8051_golden_model_1.SP [4]);
  and (_13517_, _13516_, \oc8051_golden_model_1.SP [5]);
  and (_13518_, _13517_, \oc8051_golden_model_1.SP [6]);
  or (_13519_, _13518_, \oc8051_golden_model_1.SP [7]);
  nand (_13520_, _13518_, \oc8051_golden_model_1.SP [7]);
  and (_13521_, _13520_, _13519_);
  or (_13522_, _13521_, _07059_);
  nor (_13523_, _07727_, _13514_);
  and (_13524_, _08768_, _07727_);
  or (_13525_, _13524_, _13523_);
  and (_13526_, _13525_, _06284_);
  and (_13527_, _13517_, \oc8051_golden_model_1.SP [0]);
  and (_13528_, _13527_, \oc8051_golden_model_1.SP [6]);
  nor (_13529_, _13528_, _13514_);
  and (_13530_, _13528_, _13514_);
  or (_13531_, _13530_, _13529_);
  and (_13532_, _13531_, _06038_);
  and (_13533_, _08498_, _07727_);
  or (_13534_, _13533_, _13523_);
  or (_13535_, _13534_, _06954_);
  and (_13536_, _07833_, \oc8051_golden_model_1.ACC [7]);
  or (_13537_, _13536_, _13523_);
  or (_13538_, _13537_, _06939_);
  or (_13539_, _06938_, \oc8051_golden_model_1.SP [7]);
  and (_13540_, _13539_, _07233_);
  and (_13541_, _13540_, _13538_);
  and (_13542_, _13521_, _06943_);
  or (_13543_, _13542_, _06102_);
  or (_13544_, _13543_, _13541_);
  and (_13545_, _13544_, _05690_);
  and (_13546_, _13545_, _13535_);
  and (_13547_, _13521_, _07272_);
  or (_13548_, _13547_, _06239_);
  or (_13549_, _13548_, _13546_);
  not (_13550_, \oc8051_golden_model_1.SP [6]);
  not (_13551_, \oc8051_golden_model_1.SP [5]);
  not (_13552_, \oc8051_golden_model_1.SP [4]);
  and (_13553_, _08403_, _13552_);
  and (_13554_, _13553_, _13551_);
  and (_13555_, _13554_, _13550_);
  and (_13556_, _13555_, _06029_);
  nor (_13557_, _13556_, _13514_);
  and (_13558_, _13556_, _13514_);
  nor (_13559_, _13558_, _13557_);
  nand (_13560_, _13559_, _06239_);
  and (_13561_, _13560_, _13549_);
  or (_13562_, _13561_, _06219_);
  or (_13563_, _13537_, _06220_);
  and (_13564_, _13563_, _07364_);
  and (_13565_, _13564_, _13562_);
  or (_13566_, _13565_, _13532_);
  and (_13567_, _13566_, _07271_);
  not (_13568_, _07271_);
  and (_13569_, _13521_, _13568_);
  or (_13570_, _13569_, _09818_);
  or (_13571_, _13570_, _13567_);
  or (_13572_, _13523_, _07012_);
  and (_13573_, _08485_, _07833_);
  or (_13574_, _13573_, _13572_);
  not (_13575_, _07727_);
  nor (_13576_, _07785_, _13575_);
  or (_13577_, _13523_, _09827_);
  or (_13578_, _13577_, _13576_);
  and (_13579_, _13578_, _05669_);
  and (_13580_, _13579_, _13574_);
  and (_13581_, _13580_, _13571_);
  and (_13582_, _08738_, _07727_);
  or (_13583_, _13582_, _13523_);
  and (_13584_, _13583_, _09833_);
  or (_13585_, _13584_, _06019_);
  or (_13586_, _13585_, _13581_);
  not (_13587_, _05724_);
  and (_13588_, _08549_, _07833_);
  or (_13589_, _13588_, _13523_);
  or (_13590_, _13589_, _06020_);
  and (_13591_, _13590_, _13587_);
  and (_13592_, _13591_, _13586_);
  and (_13593_, _13521_, _05724_);
  or (_13594_, _13593_, _06112_);
  or (_13595_, _13594_, _13592_);
  and (_13596_, _08760_, _07833_);
  or (_13597_, _13596_, _13523_);
  or (_13598_, _13597_, _08751_);
  and (_13599_, _13598_, _08756_);
  and (_13600_, _13599_, _13595_);
  or (_13601_, _13600_, _13526_);
  and (_13602_, _13601_, _07032_);
  or (_13603_, _13523_, _07788_);
  and (_13604_, _13589_, _06108_);
  and (_13605_, _13604_, _13603_);
  or (_13606_, _13605_, _13602_);
  and (_13607_, _13606_, _12494_);
  and (_13608_, _13521_, _05736_);
  or (_13609_, _13608_, _06130_);
  and (_13610_, _13537_, _06277_);
  and (_13611_, _13610_, _13603_);
  or (_13612_, _13611_, _13609_);
  or (_13613_, _13612_, _13607_);
  and (_13614_, _08759_, _07727_);
  or (_13615_, _13523_, _08777_);
  or (_13616_, _13615_, _13614_);
  and (_13617_, _13616_, _13613_);
  or (_13618_, _13617_, _06292_);
  not (_13619_, _06298_);
  nor (_13620_, _08767_, _13575_);
  or (_13621_, _13523_, _08782_);
  or (_13622_, _13621_, _13620_);
  and (_13623_, _13622_, _13619_);
  and (_13624_, _13623_, _13618_);
  or (_13625_, _13555_, \oc8051_golden_model_1.SP [7]);
  nand (_13626_, _13555_, \oc8051_golden_model_1.SP [7]);
  and (_13627_, _13626_, _13625_);
  and (_13628_, _13627_, _06298_);
  or (_13629_, _13628_, _05732_);
  or (_13630_, _13629_, _13624_);
  or (_13631_, _13521_, _05734_);
  and (_13632_, _13631_, _13630_);
  or (_13633_, _13632_, _06049_);
  or (_13634_, _13627_, _06050_);
  and (_13635_, _13634_, _06718_);
  and (_13636_, _13635_, _13633_);
  and (_13637_, _13534_, _06316_);
  or (_13638_, _13637_, _07458_);
  or (_13639_, _13638_, _13636_);
  and (_13640_, _13639_, _13522_);
  or (_13641_, _13640_, _06047_);
  and (_13642_, _08279_, _07727_);
  or (_13643_, _13523_, _06048_);
  or (_13644_, _13643_, _13642_);
  and (_13645_, _13644_, _01336_);
  and (_13646_, _13645_, _13641_);
  or (_13648_, _13646_, _13515_);
  and (_40776_, _13648_, _42882_);
  and (_13649_, _01340_, \oc8051_golden_model_1.SBUF [7]);
  not (_13650_, _07681_);
  and (_13651_, _13650_, \oc8051_golden_model_1.SBUF [7]);
  nor (_13652_, _08767_, _13650_);
  or (_13653_, _13652_, _13651_);
  and (_13654_, _13653_, _06292_);
  or (_13655_, _13651_, _07788_);
  and (_13656_, _08549_, _07681_);
  or (_13658_, _13656_, _13651_);
  and (_13659_, _13658_, _06108_);
  and (_13660_, _13659_, _13655_);
  and (_13661_, _08768_, _07681_);
  or (_13662_, _13661_, _13651_);
  and (_13663_, _13662_, _06284_);
  or (_13664_, _13658_, _06020_);
  and (_13665_, _08498_, _07681_);
  or (_13666_, _13665_, _13651_);
  or (_13667_, _13666_, _06954_);
  and (_13669_, _07681_, \oc8051_golden_model_1.ACC [7]);
  or (_13670_, _13669_, _13651_);
  and (_13671_, _13670_, _06938_);
  and (_13672_, _06939_, \oc8051_golden_model_1.SBUF [7]);
  or (_13673_, _13672_, _06102_);
  or (_13674_, _13673_, _13671_);
  and (_13675_, _13674_, _06848_);
  and (_13676_, _13675_, _13667_);
  nor (_13677_, _07785_, _13650_);
  or (_13678_, _13677_, _13651_);
  and (_13680_, _13678_, _06239_);
  or (_13681_, _13680_, _13676_);
  and (_13682_, _13681_, _06220_);
  and (_13683_, _13670_, _06219_);
  or (_13684_, _13683_, _09818_);
  or (_13685_, _13684_, _13682_);
  and (_13686_, _08485_, _07681_);
  or (_13687_, _13651_, _07012_);
  or (_13688_, _13687_, _13686_);
  or (_13689_, _13678_, _09827_);
  and (_13691_, _13689_, _05669_);
  and (_13692_, _13691_, _13688_);
  and (_13693_, _13692_, _13685_);
  and (_13694_, _08738_, _07681_);
  or (_13695_, _13694_, _13651_);
  and (_13696_, _13695_, _09833_);
  or (_13697_, _13696_, _06019_);
  or (_13698_, _13697_, _13693_);
  and (_13699_, _13698_, _13664_);
  or (_13700_, _13699_, _06112_);
  and (_13702_, _08760_, _07681_);
  or (_13703_, _13651_, _08751_);
  or (_13704_, _13703_, _13702_);
  and (_13705_, _13704_, _08756_);
  and (_13706_, _13705_, _13700_);
  or (_13707_, _13706_, _13663_);
  and (_13708_, _13707_, _07032_);
  or (_13709_, _13708_, _13660_);
  and (_13710_, _13709_, _06278_);
  and (_13711_, _13670_, _06277_);
  and (_13713_, _13711_, _13655_);
  or (_13714_, _13713_, _06130_);
  or (_13715_, _13714_, _13710_);
  and (_13716_, _08759_, _07681_);
  or (_13717_, _13651_, _08777_);
  or (_13718_, _13717_, _13716_);
  and (_13719_, _13718_, _08782_);
  and (_13720_, _13719_, _13715_);
  or (_13721_, _13720_, _13654_);
  and (_13722_, _13721_, _06718_);
  and (_13724_, _13666_, _06316_);
  or (_13725_, _13724_, _06047_);
  or (_13726_, _13725_, _13722_);
  and (_13727_, _08279_, _07681_);
  or (_13728_, _13651_, _06048_);
  or (_13729_, _13728_, _13727_);
  and (_13730_, _13729_, _01336_);
  and (_13731_, _13730_, _13726_);
  or (_13732_, _13731_, _13649_);
  and (_40777_, _13732_, _42882_);
  nor (_13734_, _01336_, _10606_);
  nor (_13735_, _08355_, _10606_);
  and (_13736_, _08374_, _08355_);
  or (_13737_, _13736_, _13735_);
  or (_13738_, _13737_, _05653_);
  not (_13739_, _10704_);
  or (_13740_, _11048_, _10703_);
  and (_13741_, _13740_, _10974_);
  nand (_13742_, _13741_, _13739_);
  nor (_13743_, _07705_, _10606_);
  not (_13745_, _07705_);
  nor (_13746_, _08767_, _13745_);
  or (_13747_, _13746_, _13743_);
  and (_13748_, _13747_, _06292_);
  and (_13749_, _08768_, _07705_);
  or (_13750_, _13749_, _13743_);
  and (_13751_, _13750_, _06284_);
  and (_13752_, _08738_, _07705_);
  or (_13753_, _13752_, _13743_);
  and (_13754_, _13753_, _09833_);
  and (_13756_, _10314_, _07788_);
  and (_13757_, _10324_, _10320_);
  nor (_13758_, _13757_, _10318_);
  nand (_13759_, _10367_, _10320_);
  or (_13760_, _13759_, _10365_);
  and (_13761_, _13760_, _13758_);
  or (_13762_, _13761_, _13756_);
  and (_13763_, _13762_, _06261_);
  not (_13764_, _06250_);
  not (_13765_, _06251_);
  nor (_13767_, _12722_, _13765_);
  nand (_13768_, _07979_, \oc8051_golden_model_1.ACC [5]);
  nor (_13769_, _07979_, \oc8051_golden_model_1.ACC [5]);
  nor (_13770_, _08272_, \oc8051_golden_model_1.ACC [4]);
  or (_13771_, _13770_, _13769_);
  and (_13772_, _13771_, _13768_);
  and (_13773_, _13772_, _12308_);
  nor (_13774_, _07787_, \oc8051_golden_model_1.ACC [7]);
  or (_13775_, _07885_, \oc8051_golden_model_1.ACC [6]);
  nor (_13776_, _13775_, _08768_);
  or (_13778_, _13776_, _13774_);
  or (_13779_, _13778_, _13773_);
  nand (_13780_, _08028_, \oc8051_golden_model_1.ACC [3]);
  nor (_13781_, _08028_, \oc8051_golden_model_1.ACC [3]);
  nor (_13782_, _08176_, \oc8051_golden_model_1.ACC [2]);
  or (_13783_, _13782_, _13781_);
  and (_13784_, _13783_, _13780_);
  nor (_13785_, _08077_, \oc8051_golden_model_1.ACC [1]);
  nor (_13786_, _08127_, _05758_);
  nor (_13787_, _13786_, _10994_);
  or (_13789_, _13787_, _13785_);
  and (_13790_, _13789_, _12300_);
  or (_13791_, _13790_, _13784_);
  and (_13792_, _13791_, _12309_);
  or (_13793_, _13792_, _13779_);
  nor (_13794_, _12310_, _06509_);
  and (_13795_, _13794_, _13793_);
  and (_13796_, _08498_, _07705_);
  or (_13797_, _13796_, _13743_);
  or (_13798_, _13797_, _06954_);
  and (_13799_, _07705_, \oc8051_golden_model_1.ACC [7]);
  or (_13800_, _13799_, _13743_);
  and (_13801_, _13800_, _06938_);
  nor (_13802_, _06938_, _10606_);
  or (_13803_, _13802_, _06102_);
  or (_13804_, _13803_, _13801_);
  and (_13805_, _13804_, _10413_);
  and (_13806_, _13805_, _13798_);
  nor (_13807_, _10431_, _10413_);
  not (_13808_, _12181_);
  nand (_13809_, _13808_, _06244_);
  or (_13810_, _13809_, _13807_);
  or (_13811_, _13810_, _13806_);
  and (_13812_, _08503_, _08355_);
  or (_13813_, _13812_, _13735_);
  or (_13814_, _13813_, _06044_);
  nor (_13815_, _07785_, _13745_);
  or (_13816_, _13815_, _13743_);
  or (_13817_, _13816_, _06848_);
  and (_13818_, _13817_, _13814_);
  and (_13819_, _13818_, _13811_);
  or (_13820_, _13819_, _06219_);
  or (_13821_, _13800_, _06220_);
  nor (_13822_, _12238_, _06039_);
  and (_13823_, _13822_, _13821_);
  and (_13824_, _13823_, _13820_);
  and (_13825_, _13737_, _06039_);
  or (_13826_, _13825_, _12256_);
  or (_13827_, _13826_, _13824_);
  not (_13828_, _12289_);
  nor (_13829_, _12284_, _12281_);
  or (_13830_, _12282_, _13829_);
  and (_13831_, _13830_, _12280_);
  nor (_13832_, _12277_, _12274_);
  nor (_13833_, _12275_, _13832_);
  or (_13834_, _13833_, _13831_);
  and (_13835_, _13834_, _12273_);
  and (_13836_, _12268_, _12269_);
  or (_13837_, _13836_, _12267_);
  and (_13838_, _13837_, _12265_);
  and (_13839_, _12263_, _07786_);
  or (_13840_, _13839_, _12260_);
  or (_13841_, _13840_, _13838_);
  or (_13842_, _13841_, _13835_);
  and (_13843_, _13842_, _13828_);
  or (_13844_, _13843_, _12255_);
  and (_13845_, _13844_, _12258_);
  and (_13846_, _13845_, _13827_);
  and (_13847_, _06513_, _06031_);
  and (_13848_, _10394_, _06031_);
  nor (_13849_, _13848_, _13847_);
  not (_13850_, _13849_);
  not (_13851_, _12145_);
  nand (_13852_, _12143_, _13851_);
  nand (_13853_, _13852_, _12142_);
  not (_13854_, _12152_);
  or (_13855_, _12154_, _13854_);
  and (_13856_, _13855_, _12148_);
  or (_13857_, _13856_, _13853_);
  and (_13858_, _13857_, _12170_);
  nand (_13859_, _12166_, _12163_);
  and (_13860_, _12164_, _13859_);
  and (_13861_, _13860_, _12162_);
  not (_13862_, _12157_);
  and (_13863_, _12159_, _13862_);
  nor (_13864_, _13863_, _08531_);
  or (_13865_, _13864_, _13861_);
  or (_13866_, _13865_, _13858_);
  and (_13867_, _13866_, _12174_);
  and (_13868_, _13867_, _13850_);
  or (_13869_, _13868_, _13846_);
  and (_13870_, _13869_, _06509_);
  or (_13871_, _13870_, _13795_);
  and (_13872_, _13871_, _12298_);
  nor (_13873_, _06799_, \oc8051_golden_model_1.ACC [1]);
  and (_13874_, _06799_, \oc8051_golden_model_1.ACC [1]);
  and (_13875_, _06016_, \oc8051_golden_model_1.ACC [0]);
  nor (_13876_, _13875_, _13874_);
  or (_13877_, _13876_, _13873_);
  and (_13878_, _13877_, _12320_);
  nand (_13879_, _05983_, \oc8051_golden_model_1.ACC [3]);
  nor (_13880_, _05983_, \oc8051_golden_model_1.ACC [3]);
  nor (_13881_, _06403_, \oc8051_golden_model_1.ACC [2]);
  or (_13882_, _13881_, _13880_);
  and (_13883_, _13882_, _13879_);
  or (_13884_, _13883_, _13878_);
  and (_13885_, _13884_, _12328_);
  nand (_13886_, _06359_, \oc8051_golden_model_1.ACC [5]);
  nor (_13887_, _06359_, \oc8051_golden_model_1.ACC [5]);
  nor (_13888_, _06758_, \oc8051_golden_model_1.ACC [4]);
  or (_13889_, _13888_, _13887_);
  and (_13890_, _13889_, _13886_);
  and (_13891_, _13890_, _12327_);
  and (_13892_, _05952_, _08393_);
  or (_13893_, _06084_, \oc8051_golden_model_1.ACC [6]);
  nor (_13894_, _13893_, _10705_);
  or (_13895_, _13894_, _13892_);
  or (_13896_, _13895_, _13891_);
  or (_13897_, _13896_, _13885_);
  nor (_13898_, _12329_, _12298_);
  and (_13899_, _13898_, _13897_);
  or (_13900_, _13899_, _12012_);
  or (_13901_, _13900_, _13872_);
  nand (_13902_, _12012_, \oc8051_golden_model_1.PSW [7]);
  and (_13903_, _13902_, _06033_);
  and (_13904_, _13903_, _13901_);
  and (_13905_, _08520_, _08355_);
  or (_13906_, _13905_, _13735_);
  and (_13907_, _13906_, _06032_);
  nor (_13908_, _13907_, _13904_);
  nor (_13909_, _13908_, _06253_);
  and (_13910_, _06253_, \oc8051_golden_model_1.PSW [7]);
  and (_13911_, _13910_, _12722_);
  or (_13912_, _13911_, _13909_);
  nor (_13913_, _09269_, _06251_);
  and (_13914_, _13913_, _13912_);
  or (_13915_, _13914_, _13767_);
  and (_13916_, _13915_, _13764_);
  or (_13917_, _12722_, \oc8051_golden_model_1.PSW [7]);
  and (_13918_, _13917_, _06250_);
  or (_13919_, _13918_, _10468_);
  or (_13920_, _13919_, _13916_);
  and (_13921_, _10250_, _10246_);
  nor (_13922_, _13921_, _10244_);
  nand (_13923_, _10252_, _10246_);
  or (_13924_, _13923_, _10485_);
  and (_13925_, _13924_, _13922_);
  or (_13926_, _10469_, _10241_);
  or (_13927_, _13926_, _13925_);
  and (_13928_, _13927_, _13920_);
  or (_13929_, _13928_, _12361_);
  and (_13930_, _10506_, _10501_);
  nor (_13931_, _13930_, _10499_);
  nand (_13932_, _10553_, _10501_);
  or (_13933_, _13932_, _10551_);
  and (_13934_, _13933_, _13931_);
  not (_13935_, _12361_);
  and (_13936_, _10495_, _08485_);
  or (_13937_, _13936_, _13935_);
  or (_13938_, _13937_, _13934_);
  and (_13939_, _13938_, _06267_);
  and (_13940_, _13939_, _13929_);
  or (_13941_, _13940_, _13763_);
  and (_13942_, _13941_, _10307_);
  and (_13943_, _10578_, _10575_);
  nor (_13944_, _13943_, _10573_);
  nand (_13945_, _10625_, _10575_);
  or (_13946_, _13945_, _10623_);
  and (_13947_, _13946_, _13944_);
  or (_13948_, _13947_, _10568_);
  and (_13949_, _13948_, _10306_);
  or (_13950_, _13949_, _09818_);
  or (_13951_, _13950_, _13942_);
  and (_13952_, _08485_, _07705_);
  or (_13953_, _13743_, _07012_);
  or (_13954_, _13953_, _13952_);
  or (_13955_, _13816_, _09827_);
  and (_13956_, _13955_, _05669_);
  and (_13957_, _13956_, _13954_);
  and (_13958_, _13957_, _13951_);
  or (_13959_, _13958_, _13754_);
  nor (_13960_, _09832_, _06089_);
  and (_13961_, _13960_, _13959_);
  nor (_13962_, _12722_, _10606_);
  and (_13963_, _13962_, _06089_);
  or (_13964_, _13963_, _06019_);
  or (_13965_, _13964_, _13961_);
  and (_13966_, _08549_, _07705_);
  or (_13967_, _13966_, _13743_);
  or (_13968_, _13967_, _06020_);
  and (_13969_, _13968_, _13965_);
  or (_13970_, _13969_, _06088_);
  nand (_13971_, _12722_, _10606_);
  or (_13972_, _13971_, _06636_);
  and (_13973_, _13972_, _13970_);
  or (_13974_, _13973_, _06112_);
  and (_13975_, _08760_, _07705_);
  or (_13976_, _13975_, _13743_);
  or (_13977_, _13976_, _08751_);
  and (_13978_, _13977_, _08756_);
  and (_13979_, _13978_, _13974_);
  or (_13980_, _13979_, _13751_);
  and (_13981_, _13980_, _07032_);
  or (_13982_, _13743_, _07788_);
  and (_13983_, _13967_, _06108_);
  and (_13984_, _13983_, _13982_);
  or (_13985_, _13984_, _13981_);
  and (_13986_, _13985_, _06278_);
  and (_13987_, _13800_, _06277_);
  and (_13988_, _13987_, _13982_);
  or (_13989_, _13988_, _06130_);
  or (_13990_, _13989_, _13986_);
  and (_13991_, _08759_, _07705_);
  or (_13992_, _13743_, _08777_);
  or (_13993_, _13992_, _13991_);
  and (_13994_, _13993_, _08782_);
  and (_13995_, _13994_, _13990_);
  or (_13996_, _13995_, _13748_);
  and (_13997_, _13996_, _10304_);
  nor (_13998_, _10243_, _08393_);
  or (_13999_, _13998_, _10300_);
  or (_14000_, _13999_, _10241_);
  and (_14001_, _14000_, _10303_);
  or (_14002_, _14001_, _10794_);
  or (_14003_, _14002_, _13997_);
  or (_14004_, _10796_, _13936_);
  nor (_14005_, _10498_, _08393_);
  or (_14006_, _14005_, _10818_);
  or (_14007_, _14006_, _14004_);
  and (_14008_, _14007_, _06289_);
  and (_14009_, _14008_, _14003_);
  nor (_14010_, _10317_, _08393_);
  or (_14011_, _14010_, _10848_);
  or (_14012_, _10824_, _13756_);
  or (_14013_, _14012_, _14011_);
  and (_14014_, _14013_, _10826_);
  or (_14015_, _14014_, _14009_);
  and (_14016_, _10572_, \oc8051_golden_model_1.ACC [7]);
  or (_14017_, _14016_, _10878_);
  or (_14018_, _10856_, _10568_);
  or (_14019_, _14018_, _14017_);
  and (_14020_, _14019_, _10855_);
  and (_14021_, _14020_, _14015_);
  nand (_14022_, _10885_, _06545_);
  and (_14023_, _14022_, _10889_);
  nand (_14024_, _10854_, \oc8051_golden_model_1.ACC [7]);
  nand (_14025_, _14024_, _14023_);
  or (_14026_, _14025_, _14021_);
  or (_14027_, _10926_, _10672_);
  nand (_14028_, _14027_, _10719_);
  nor (_14029_, _14028_, _14023_);
  nor (_14030_, _14029_, _06693_);
  and (_14031_, _14030_, _14026_);
  and (_14032_, _14028_, _06693_);
  or (_14033_, _14032_, _10932_);
  or (_14034_, _14033_, _14031_);
  and (_14035_, _10966_, _10693_);
  nor (_14036_, _10935_, _10692_);
  nor (_14037_, _14036_, _10691_);
  or (_14038_, _14037_, _10934_);
  or (_14039_, _14038_, _14035_);
  and (_14040_, _14039_, _06052_);
  and (_14041_, _14040_, _14034_);
  not (_14042_, _08767_);
  not (_14043_, _08766_);
  nand (_14044_, _11008_, _14043_);
  and (_14045_, _14044_, _06051_);
  and (_14046_, _14045_, _14042_);
  or (_14047_, _14046_, _10974_);
  or (_14048_, _14047_, _14041_);
  and (_14049_, _14048_, _13742_);
  or (_14050_, _14049_, _06316_);
  nor (_14051_, _13797_, _06718_);
  nor (_14052_, _14051_, _11064_);
  and (_14053_, _14052_, _14050_);
  and (_14054_, _11064_, \oc8051_golden_model_1.ACC [0]);
  or (_14055_, _14054_, _05652_);
  or (_14056_, _14055_, _14053_);
  and (_14057_, _14056_, _13738_);
  or (_14058_, _14057_, _06047_);
  and (_14059_, _08279_, _07705_);
  or (_14060_, _13743_, _06048_);
  or (_14061_, _14060_, _14059_);
  and (_14062_, _14061_, _01336_);
  and (_14063_, _14062_, _14058_);
  or (_14064_, _14063_, _13734_);
  and (_40778_, _14064_, _42882_);
  and (_14065_, _12112_, _06127_);
  not (_14066_, _11952_);
  nor (_14067_, _14066_, _06127_);
  or (_14068_, _14067_, _14065_);
  nor (_14069_, _08403_, _07360_);
  not (_14070_, _14069_);
  and (_14071_, _14070_, _07628_);
  and (_14072_, _14071_, _07081_);
  not (_14073_, _14072_);
  or (_14074_, _14073_, _14068_);
  nor (_14075_, _07476_, _07305_);
  nor (_14076_, _14075_, _07615_);
  nor (_14077_, _07305_, _07074_);
  nor (_14078_, _14077_, _07306_);
  and (_14079_, _14078_, _07304_);
  and (_14080_, _14079_, _14076_);
  nand (_14081_, _06127_, \oc8051_golden_model_1.PC [0]);
  nand (_14082_, _12302_, _08783_);
  or (_14083_, _08127_, _08672_);
  and (_14084_, _08127_, _08672_);
  not (_14085_, _14084_);
  and (_14086_, _14085_, _14083_);
  and (_14087_, _14086_, _08752_);
  or (_14088_, _07009_, _06931_);
  or (_14089_, _08127_, _06233_);
  nor (_14090_, _12615_, _12591_);
  or (_14091_, _14090_, _08378_);
  nor (_14092_, _08127_, _08381_);
  nand (_14093_, _08384_, _06931_);
  nand (_14094_, _06943_, _05346_);
  or (_14095_, _06943_, \oc8051_golden_model_1.ACC [0]);
  and (_14096_, _14095_, _14094_);
  nor (_14097_, _14096_, _08384_);
  nor (_14098_, _14097_, _06955_);
  and (_14099_, _14098_, _14093_);
  or (_14100_, _14099_, _14092_);
  and (_14101_, _14100_, _08380_);
  nand (_14102_, _12615_, _12592_);
  and (_14103_, _14102_, _06953_);
  or (_14104_, _14103_, _07272_);
  or (_14105_, _14104_, _14101_);
  nor (_14106_, _05690_, \oc8051_golden_model_1.PC [0]);
  nor (_14107_, _14106_, _06963_);
  and (_14108_, _14107_, _14105_);
  and (_14109_, _06963_, _06931_);
  or (_14110_, _14109_, _06975_);
  or (_14111_, _14110_, _14108_);
  and (_14112_, _14111_, _14091_);
  or (_14113_, _14112_, _06038_);
  or (_14114_, _08127_, _07364_);
  and (_14115_, _14114_, _06036_);
  and (_14116_, _14115_, _14113_);
  nor (_14117_, _12616_, _06036_);
  and (_14118_, _14117_, _14102_);
  or (_14119_, _14118_, _14116_);
  and (_14120_, _14119_, _05686_);
  or (_14121_, _05686_, _05346_);
  nand (_14122_, _06233_, _14121_);
  or (_14123_, _14122_, _14120_);
  and (_14124_, _14123_, _14089_);
  or (_14125_, _14124_, _06992_);
  and (_14126_, _09120_, _06053_);
  nand (_14127_, _08124_, _06992_);
  or (_14128_, _14127_, _14126_);
  and (_14129_, _14128_, _14125_);
  or (_14130_, _14129_, _06991_);
  nand (_14131_, _12591_, _10606_);
  and (_14132_, _14131_, _14102_);
  or (_14133_, _14132_, _07308_);
  and (_14134_, _14133_, _05673_);
  and (_14135_, _14134_, _14130_);
  or (_14136_, _05673_, _05346_);
  nand (_14137_, _07009_, _14136_);
  or (_14138_, _14137_, _14135_);
  and (_14139_, _14138_, _14088_);
  or (_14140_, _14139_, _07013_);
  or (_14141_, _09120_, _07231_);
  and (_14142_, _14141_, _08545_);
  and (_14143_, _14142_, _14140_);
  and (_14144_, _08332_, _06931_);
  and (_14145_, _08668_, \oc8051_golden_model_1.SCON [0]);
  and (_14146_, _08677_, \oc8051_golden_model_1.SBUF [0]);
  or (_14147_, _14146_, _14145_);
  and (_14148_, _08660_, \oc8051_golden_model_1.P0 [0]);
  and (_14149_, _08682_, \oc8051_golden_model_1.P1 [0]);
  or (_14150_, _14149_, _14148_);
  or (_14151_, _14150_, _14147_);
  and (_14152_, _08680_, \oc8051_golden_model_1.TCON [0]);
  and (_14153_, _08654_, \oc8051_golden_model_1.ACC [0]);
  or (_14154_, _14153_, _14152_);
  and (_14155_, _08675_, \oc8051_golden_model_1.TMOD [0]);
  and (_14156_, _08702_, \oc8051_golden_model_1.TL0 [0]);
  or (_14157_, _14156_, _14155_);
  or (_14158_, _14157_, _14154_);
  and (_14159_, _08693_, \oc8051_golden_model_1.IE [0]);
  and (_14160_, _08695_, \oc8051_golden_model_1.P3 [0]);
  or (_14161_, _14160_, _14159_);
  and (_14162_, _08687_, \oc8051_golden_model_1.P2 [0]);
  and (_14163_, _08690_, \oc8051_golden_model_1.IP [0]);
  or (_14164_, _14163_, _14162_);
  or (_14165_, _14164_, _14161_);
  and (_14166_, _08650_, \oc8051_golden_model_1.B [0]);
  and (_14167_, _08704_, \oc8051_golden_model_1.PSW [0]);
  or (_14168_, _14167_, _14166_);
  or (_14169_, _14168_, _14165_);
  or (_14170_, _14169_, _14158_);
  or (_14171_, _14170_, _14151_);
  and (_14172_, _08732_, \oc8051_golden_model_1.PCON [0]);
  and (_14173_, _08725_, \oc8051_golden_model_1.TH1 [0]);
  and (_14174_, _08712_, \oc8051_golden_model_1.TH0 [0]);
  or (_14175_, _14174_, _14173_);
  or (_14176_, _14175_, _14172_);
  and (_14177_, _08716_, \oc8051_golden_model_1.TL1 [0]);
  and (_14178_, _08723_, \oc8051_golden_model_1.DPH [0]);
  or (_14179_, _14178_, _14177_);
  and (_14180_, _08728_, \oc8051_golden_model_1.DPL [0]);
  and (_14181_, _08719_, \oc8051_golden_model_1.SP [0]);
  or (_14182_, _14181_, _14180_);
  or (_14183_, _14182_, _14179_);
  or (_14184_, _14183_, _14176_);
  or (_14185_, _14184_, _14171_);
  or (_14186_, _14185_, _14144_);
  and (_14187_, _14186_, _07010_);
  or (_14188_, _14187_, _08743_);
  or (_14189_, _14188_, _14143_);
  and (_14190_, _08743_, _06016_);
  nor (_14191_, _14190_, _06021_);
  and (_14192_, _14191_, _14189_);
  and (_14193_, _08672_, _06021_);
  or (_14194_, _14193_, _05724_);
  or (_14195_, _14194_, _14192_);
  and (_14196_, _05724_, _05346_);
  nor (_14197_, _14196_, _08752_);
  and (_14198_, _14197_, _14195_);
  or (_14199_, _14198_, _14087_);
  and (_14200_, _14199_, _08765_);
  nor (_14201_, _12303_, _08765_);
  or (_14202_, _14201_, _14200_);
  and (_14203_, _14202_, _08764_);
  and (_14204_, _14084_, _08301_);
  or (_14205_, _14204_, _14203_);
  and (_14206_, _14205_, _08300_);
  and (_14207_, _10995_, _07031_);
  or (_14208_, _14207_, _05736_);
  or (_14209_, _14208_, _14206_);
  and (_14210_, _05736_, _05346_);
  nor (_14211_, _14210_, _08778_);
  and (_14212_, _14211_, _14209_);
  and (_14213_, _14083_, _08778_);
  or (_14214_, _14213_, _08783_);
  or (_14215_, _14214_, _14212_);
  and (_14216_, _14215_, _14082_);
  or (_14217_, _14216_, _05732_);
  nand (_14218_, _05732_, _05346_);
  and (_14219_, _14218_, _08287_);
  and (_14220_, _14219_, _14217_);
  nand (_14221_, _07052_, _06931_);
  and (_14222_, _14221_, _12750_);
  or (_14223_, _14222_, _14220_);
  nand (_14224_, _09120_, _07051_);
  and (_14225_, _14224_, _08797_);
  and (_14226_, _14225_, _14223_);
  nor (_14227_, _08127_, _08797_);
  or (_14228_, _14227_, _06127_);
  or (_14229_, _14228_, _14226_);
  and (_14230_, _14229_, _14081_);
  or (_14231_, _14230_, _05752_);
  and (_14232_, _05752_, _05346_);
  nor (_14233_, _14232_, _07058_);
  and (_14234_, _14233_, _14231_);
  not (_14235_, _09154_);
  and (_14236_, _14090_, _07058_);
  or (_14237_, _14236_, _14235_);
  or (_14238_, _14237_, _14234_);
  nand (_14239_, _14235_, _06931_);
  and (_14240_, _14239_, _07069_);
  and (_14241_, _14240_, _14238_);
  nor (_14242_, _09120_, _07069_);
  or (_14243_, _14242_, _07067_);
  or (_14244_, _14243_, _14241_);
  nand (_14245_, _08127_, _07067_);
  and (_14246_, _14245_, _07304_);
  and (_14247_, _14246_, _14244_);
  and (_14248_, _14247_, _14080_);
  or (_14249_, _14080_, _06505_);
  nand (_14250_, _14249_, _14073_);
  or (_14251_, _14250_, _14248_);
  and (_40792_, _14251_, _14074_);
  or (_14252_, _14080_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_14253_, _14252_, _14073_);
  not (_14254_, _14080_);
  nor (_14255_, _09162_, _08291_);
  and (_14256_, _14255_, _14235_);
  nor (_14257_, _14255_, _06866_);
  or (_14258_, _14257_, _07210_);
  and (_14259_, _05732_, _05312_);
  nand (_14260_, _08077_, _06832_);
  nor (_14261_, _08077_, _06832_);
  not (_14262_, _14261_);
  and (_14263_, _14262_, _14260_);
  and (_14264_, _14263_, _08752_);
  nand (_14265_, _07132_, _08541_);
  nand (_14266_, _12588_, _12566_);
  nand (_14267_, _07726_, _10606_);
  and (_14268_, _14267_, _06991_);
  and (_14269_, _14268_, _14266_);
  or (_14270_, _12150_, _05952_);
  nand (_14271_, _14270_, _08075_);
  and (_14272_, _14271_, _06992_);
  nor (_14273_, _12588_, _07726_);
  or (_14274_, _14273_, _08378_);
  nand (_14275_, _14255_, _08384_);
  and (_14276_, _06943_, _05312_);
  and (_14277_, _11988_, _06042_);
  nor (_14278_, _06943_, _05784_);
  or (_14279_, _14278_, _14277_);
  or (_14280_, _14279_, _07139_);
  or (_14281_, _14280_, _14276_);
  and (_14282_, _14281_, _14275_);
  and (_14283_, _14282_, _08381_);
  nor (_14284_, _08491_, _08128_);
  nor (_14285_, _14284_, _08381_);
  or (_14286_, _14285_, _14283_);
  or (_14287_, _14286_, _06953_);
  or (_14288_, _14266_, _08380_);
  and (_14289_, _14288_, _14287_);
  or (_14290_, _14289_, _07272_);
  nor (_14291_, _05690_, _05312_);
  nor (_14292_, _14291_, _06963_);
  and (_14293_, _14292_, _14290_);
  and (_14294_, _09161_, _06963_);
  or (_14295_, _14294_, _06975_);
  or (_14296_, _14295_, _14293_);
  and (_14297_, _14296_, _14274_);
  or (_14298_, _14297_, _06038_);
  nand (_14299_, _08077_, _06038_);
  and (_14300_, _14299_, _06036_);
  and (_14301_, _14300_, _14298_);
  not (_14302_, _12589_);
  and (_14303_, _14266_, _14302_);
  and (_14304_, _14303_, _06035_);
  or (_14305_, _14304_, _14301_);
  and (_14306_, _14305_, _05686_);
  or (_14307_, _05686_, \oc8051_golden_model_1.PC [1]);
  nand (_14308_, _06233_, _14307_);
  or (_14309_, _14308_, _14306_);
  nand (_14310_, _08077_, _06573_);
  and (_14311_, _14310_, _06993_);
  and (_14312_, _14311_, _14309_);
  or (_14313_, _14312_, _14272_);
  and (_14314_, _14313_, _07308_);
  or (_14315_, _14314_, _14269_);
  and (_14316_, _14315_, _05673_);
  or (_14317_, _05673_, \oc8051_golden_model_1.PC [1]);
  nand (_14318_, _07009_, _14317_);
  or (_14319_, _14318_, _14316_);
  and (_14320_, _14319_, _14265_);
  or (_14321_, _14320_, _07013_);
  or (_14322_, _09075_, _07231_);
  and (_14323_, _14322_, _08545_);
  and (_14324_, _14323_, _14321_);
  nor (_14325_, _08549_, _07132_);
  and (_14326_, _08675_, \oc8051_golden_model_1.TMOD [1]);
  and (_14327_, _08682_, \oc8051_golden_model_1.P1 [1]);
  or (_14328_, _14327_, _14326_);
  and (_14329_, _08702_, \oc8051_golden_model_1.TL0 [1]);
  and (_14330_, _08650_, \oc8051_golden_model_1.B [1]);
  or (_14331_, _14330_, _14329_);
  or (_14332_, _14331_, _14328_);
  and (_14333_, _08660_, \oc8051_golden_model_1.P0 [1]);
  and (_14334_, _08680_, \oc8051_golden_model_1.TCON [1]);
  or (_14335_, _14334_, _14333_);
  and (_14336_, _08668_, \oc8051_golden_model_1.SCON [1]);
  and (_14337_, _08704_, \oc8051_golden_model_1.PSW [1]);
  or (_14338_, _14337_, _14336_);
  or (_14339_, _14338_, _14335_);
  and (_14340_, _08693_, \oc8051_golden_model_1.IE [1]);
  and (_14341_, _08690_, \oc8051_golden_model_1.IP [1]);
  or (_14342_, _14341_, _14340_);
  and (_14343_, _08687_, \oc8051_golden_model_1.P2 [1]);
  and (_14344_, _08695_, \oc8051_golden_model_1.P3 [1]);
  or (_14345_, _14344_, _14343_);
  or (_14346_, _14345_, _14342_);
  and (_14347_, _08677_, \oc8051_golden_model_1.SBUF [1]);
  and (_14348_, _08654_, \oc8051_golden_model_1.ACC [1]);
  or (_14349_, _14348_, _14347_);
  or (_14350_, _14349_, _14346_);
  or (_14351_, _14350_, _14339_);
  or (_14352_, _14351_, _14332_);
  and (_14353_, _08716_, \oc8051_golden_model_1.TL1 [1]);
  and (_14354_, _08732_, \oc8051_golden_model_1.PCON [1]);
  and (_14355_, _08725_, \oc8051_golden_model_1.TH1 [1]);
  or (_14356_, _14355_, _14354_);
  or (_14357_, _14356_, _14353_);
  and (_14358_, _08712_, \oc8051_golden_model_1.TH0 [1]);
  and (_14359_, _08719_, \oc8051_golden_model_1.SP [1]);
  or (_14360_, _14359_, _14358_);
  and (_14361_, _08728_, \oc8051_golden_model_1.DPL [1]);
  and (_14362_, _08723_, \oc8051_golden_model_1.DPH [1]);
  or (_14363_, _14362_, _14361_);
  or (_14364_, _14363_, _14360_);
  or (_14365_, _14364_, _14357_);
  or (_14366_, _14365_, _14352_);
  or (_14367_, _14366_, _14325_);
  and (_14368_, _14367_, _07010_);
  or (_14369_, _14368_, _08743_);
  or (_14370_, _14369_, _14324_);
  and (_14371_, _08743_, _06799_);
  nor (_14372_, _14371_, _06021_);
  and (_14373_, _14372_, _14370_);
  and (_14374_, _08699_, _06021_);
  or (_14375_, _14374_, _05724_);
  or (_14376_, _14375_, _14373_);
  and (_14377_, _05724_, \oc8051_golden_model_1.PC [1]);
  nor (_14378_, _14377_, _08752_);
  and (_14379_, _14378_, _14376_);
  or (_14380_, _14379_, _14264_);
  and (_14381_, _14380_, _08765_);
  and (_14382_, _10994_, _08757_);
  or (_14383_, _14382_, _08301_);
  or (_14384_, _14383_, _14381_);
  or (_14385_, _14261_, _08764_);
  and (_14386_, _14385_, _08300_);
  and (_14387_, _14386_, _14384_);
  and (_14388_, _10992_, _07031_);
  or (_14389_, _14388_, _05736_);
  or (_14390_, _14389_, _14387_);
  and (_14391_, _05736_, \oc8051_golden_model_1.PC [1]);
  nor (_14392_, _14391_, _08778_);
  and (_14393_, _14392_, _14390_);
  and (_14394_, _14260_, _08778_);
  or (_14395_, _14394_, _08783_);
  or (_14396_, _14395_, _14393_);
  nand (_14397_, _10993_, _08783_);
  and (_14398_, _14397_, _05734_);
  and (_14399_, _14398_, _14396_);
  nor (_14400_, _14399_, _14259_);
  nor (_14401_, _14400_, _07278_);
  not (_14402_, _14255_);
  nand (_14403_, _14402_, _07278_);
  nand (_14404_, _14403_, _06459_);
  or (_14405_, _14404_, _14401_);
  or (_14406_, _14402_, _06459_);
  and (_14407_, _14406_, _06866_);
  and (_14408_, _14407_, _14405_);
  or (_14409_, _14408_, _14258_);
  nand (_14410_, _14255_, _07210_);
  and (_14411_, _14410_, _07052_);
  and (_14412_, _14411_, _14409_);
  nor (_14413_, _09183_, _09121_);
  nor (_14414_, _14413_, _07052_);
  or (_14415_, _14414_, _14412_);
  and (_14416_, _14415_, _08797_);
  nor (_14417_, _14284_, _08797_);
  or (_14418_, _14417_, _06127_);
  or (_14419_, _14418_, _14416_);
  nand (_14420_, _06127_, _12086_);
  and (_14421_, _14420_, _12766_);
  and (_14422_, _14421_, _14419_);
  and (_14423_, _05752_, _05312_);
  or (_14424_, _07058_, _14423_);
  or (_14425_, _14424_, _14422_);
  or (_14426_, _14273_, _07295_);
  and (_14427_, _14426_, _09154_);
  and (_14428_, _14427_, _14425_);
  or (_14429_, _14428_, _14256_);
  and (_14430_, _14429_, _07069_);
  and (_14431_, _14413_, _07068_);
  or (_14432_, _14431_, _07067_);
  or (_14433_, _14432_, _14430_);
  or (_14434_, _14284_, _07232_);
  and (_14435_, _14434_, _07304_);
  and (_14436_, _14435_, _14433_);
  or (_14437_, _14436_, _14254_);
  and (_14438_, _14437_, _14253_);
  nor (_14439_, _07627_, _01340_);
  and (_14440_, _14439_, _42882_);
  nor (_14441_, _07627_, _06029_);
  and (_14442_, _14441_, _01336_);
  and (_14443_, _14442_, _42882_);
  not (_14444_, _14443_);
  or (_14445_, _07627_, \oc8051_golden_model_1.SP [1]);
  or (_14446_, _14445_, _01340_);
  or (_14447_, _14446_, rst);
  and (_14448_, _14447_, _14444_);
  not (_14449_, _07622_);
  or (_14450_, _07627_, _14449_);
  or (_14451_, _14450_, _01340_);
  or (_14452_, _14451_, rst);
  not (_14453_, _07625_);
  or (_14454_, _07627_, _14453_);
  or (_14455_, _14454_, _01340_);
  or (_14456_, _14455_, rst);
  and (_14457_, _14456_, _14452_);
  and (_14458_, _14457_, _14448_);
  and (_14459_, _14458_, _14440_);
  not (_14460_, _07627_);
  not (_14461_, _11900_);
  nor (_14462_, _14461_, _06127_);
  and (_14463_, _12051_, _06127_);
  or (_14464_, _14463_, _14462_);
  and (_14465_, _14464_, _14460_);
  and (_14466_, _14465_, _01336_);
  and (_14467_, _14466_, _42882_);
  and (_14468_, _14467_, _14459_);
  or (_40793_, _14468_, _14438_);
  or (_14469_, _14080_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_14470_, _14469_, _14073_);
  nor (_14471_, _09162_, _09160_);
  nor (_14472_, _14471_, _09163_);
  and (_14473_, _14472_, _14235_);
  and (_14474_, _05803_, _05732_);
  nand (_14475_, _07530_, _08541_);
  or (_14476_, _09030_, _05952_);
  nand (_14477_, _14476_, _08174_);
  and (_14478_, _14477_, _06992_);
  nor (_14479_, _12564_, _07732_);
  or (_14480_, _14479_, _08378_);
  and (_14481_, _08291_, _07530_);
  nor (_14482_, _08291_, _07530_);
  or (_14483_, _14482_, _14481_);
  or (_14484_, _14483_, _08383_);
  nor (_14485_, _06943_, _09956_);
  and (_14486_, _06943_, _05803_);
  or (_14487_, _14486_, _08384_);
  or (_14488_, _14487_, _14485_);
  and (_14489_, _14488_, _14484_);
  and (_14490_, _14489_, _08381_);
  nand (_14491_, _08491_, _08176_);
  or (_14492_, _08491_, _08176_);
  nand (_14493_, _14492_, _14491_);
  and (_14494_, _14493_, _06955_);
  or (_14495_, _14494_, _14490_);
  and (_14496_, _14495_, _08380_);
  nand (_14497_, _12564_, _12542_);
  and (_14498_, _14497_, _06953_);
  or (_14499_, _14498_, _07272_);
  or (_14500_, _14499_, _14496_);
  nor (_14501_, _05803_, _05690_);
  nor (_14502_, _14501_, _06963_);
  and (_14503_, _14502_, _14500_);
  and (_14504_, _09160_, _06963_);
  or (_14505_, _14504_, _06975_);
  or (_14506_, _14505_, _14503_);
  and (_14507_, _14506_, _14480_);
  or (_14508_, _14507_, _06038_);
  nand (_14509_, _08176_, _06038_);
  and (_14510_, _14509_, _06036_);
  and (_14511_, _14510_, _14508_);
  not (_14512_, _12565_);
  and (_14513_, _14497_, _14512_);
  and (_14514_, _14513_, _06035_);
  or (_14515_, _14514_, _14511_);
  and (_14516_, _14515_, _05686_);
  or (_14517_, _05804_, _05686_);
  nand (_14518_, _06233_, _14517_);
  or (_14519_, _14518_, _14516_);
  nand (_14520_, _08176_, _06573_);
  and (_14521_, _14520_, _06993_);
  and (_14522_, _14521_, _14519_);
  or (_14523_, _14522_, _14478_);
  and (_14524_, _14523_, _07308_);
  nand (_14525_, _07732_, _10606_);
  and (_14526_, _14525_, _06991_);
  and (_14527_, _14526_, _14497_);
  or (_14528_, _14527_, _14524_);
  and (_14529_, _14528_, _05673_);
  or (_14530_, _05804_, _05673_);
  nand (_14531_, _07009_, _14530_);
  or (_14532_, _14531_, _14529_);
  and (_14533_, _14532_, _14475_);
  or (_14534_, _14533_, _07013_);
  or (_14535_, _09182_, _07231_);
  and (_14536_, _14535_, _08545_);
  and (_14537_, _14536_, _14534_);
  nor (_14538_, _08549_, _07530_);
  and (_14539_, _08668_, \oc8051_golden_model_1.SCON [2]);
  and (_14540_, _08650_, \oc8051_golden_model_1.B [2]);
  or (_14541_, _14540_, _14539_);
  and (_14542_, _08702_, \oc8051_golden_model_1.TL0 [2]);
  and (_14543_, _08704_, \oc8051_golden_model_1.PSW [2]);
  or (_14544_, _14543_, _14542_);
  or (_14545_, _14544_, _14541_);
  and (_14546_, _08675_, \oc8051_golden_model_1.TMOD [2]);
  and (_14547_, _08682_, \oc8051_golden_model_1.P1 [2]);
  or (_14548_, _14547_, _14546_);
  and (_14549_, _08680_, \oc8051_golden_model_1.TCON [2]);
  and (_14550_, _08677_, \oc8051_golden_model_1.SBUF [2]);
  or (_14551_, _14550_, _14549_);
  or (_14552_, _14551_, _14548_);
  and (_14553_, _08687_, \oc8051_golden_model_1.P2 [2]);
  and (_14554_, _08690_, \oc8051_golden_model_1.IP [2]);
  or (_14555_, _14554_, _14553_);
  and (_14556_, _08693_, \oc8051_golden_model_1.IE [2]);
  and (_14557_, _08695_, \oc8051_golden_model_1.P3 [2]);
  or (_14558_, _14557_, _14556_);
  or (_14559_, _14558_, _14555_);
  and (_14560_, _08660_, \oc8051_golden_model_1.P0 [2]);
  and (_14561_, _08654_, \oc8051_golden_model_1.ACC [2]);
  or (_14562_, _14561_, _14560_);
  or (_14563_, _14562_, _14559_);
  or (_14564_, _14563_, _14552_);
  or (_14565_, _14564_, _14545_);
  and (_14566_, _08725_, \oc8051_golden_model_1.TH1 [2]);
  and (_14567_, _08716_, \oc8051_golden_model_1.TL1 [2]);
  and (_14568_, _08719_, \oc8051_golden_model_1.SP [2]);
  or (_14569_, _14568_, _14567_);
  or (_14570_, _14569_, _14566_);
  and (_14571_, _08728_, \oc8051_golden_model_1.DPL [2]);
  and (_14572_, _08732_, \oc8051_golden_model_1.PCON [2]);
  or (_14573_, _14572_, _14571_);
  and (_14574_, _08723_, \oc8051_golden_model_1.DPH [2]);
  and (_14575_, _08712_, \oc8051_golden_model_1.TH0 [2]);
  or (_14576_, _14575_, _14574_);
  or (_14577_, _14576_, _14573_);
  or (_14578_, _14577_, _14570_);
  or (_14579_, _14578_, _14565_);
  or (_14580_, _14579_, _14538_);
  and (_14581_, _14580_, _07010_);
  or (_14582_, _14581_, _08743_);
  or (_14583_, _14582_, _14537_);
  and (_14584_, _08743_, _06403_);
  nor (_14585_, _14584_, _06021_);
  and (_14586_, _14585_, _14583_);
  and (_14587_, _08730_, _06021_);
  or (_14588_, _14587_, _05724_);
  or (_14589_, _14588_, _14586_);
  and (_14590_, _05804_, _05724_);
  nor (_14591_, _14590_, _08752_);
  and (_14592_, _14591_, _14589_);
  nand (_14593_, _08176_, _06445_);
  nor (_14594_, _08176_, _06445_);
  not (_14595_, _14594_);
  and (_14596_, _14595_, _14593_);
  and (_14597_, _14596_, _08752_);
  or (_14598_, _14597_, _14592_);
  and (_14599_, _14598_, _08765_);
  and (_14600_, _10991_, _08757_);
  or (_14601_, _14600_, _14599_);
  and (_14602_, _14601_, _08764_);
  and (_14603_, _14594_, _08301_);
  or (_14604_, _14603_, _14602_);
  and (_14605_, _14604_, _08300_);
  and (_14606_, _10989_, _07031_);
  or (_14607_, _14606_, _05736_);
  or (_14608_, _14607_, _14605_);
  and (_14609_, _05804_, _05736_);
  nor (_14610_, _14609_, _08778_);
  and (_14611_, _14610_, _14608_);
  and (_14612_, _14593_, _08778_);
  or (_14613_, _14612_, _08783_);
  or (_14614_, _14613_, _14611_);
  nand (_14615_, _10990_, _08783_);
  and (_14616_, _14615_, _05734_);
  and (_14617_, _14616_, _14614_);
  or (_14618_, _14617_, _14474_);
  and (_14619_, _14618_, _08283_);
  and (_14620_, _06133_, _05495_);
  not (_14621_, _14620_);
  and (_14622_, _08285_, _14621_);
  not (_14623_, _14622_);
  or (_14624_, _14623_, _06708_);
  and (_14625_, _14483_, _08282_);
  or (_14626_, _14625_, _14624_);
  or (_14627_, _14626_, _14619_);
  not (_14628_, _14624_);
  or (_14629_, _14628_, _14483_);
  and (_14630_, _14629_, _07052_);
  and (_14631_, _14630_, _14627_);
  nor (_14632_, _09121_, _09030_);
  or (_14633_, _14632_, _09122_);
  and (_14634_, _14633_, _07051_);
  or (_14635_, _14634_, _14631_);
  and (_14636_, _14635_, _08797_);
  and (_14637_, _14493_, _07050_);
  or (_14638_, _14637_, _06127_);
  or (_14639_, _14638_, _14636_);
  nand (_14640_, _12084_, _06127_);
  and (_14641_, _14640_, _12766_);
  and (_14642_, _14641_, _14639_);
  and (_14643_, _05803_, _05752_);
  or (_14644_, _07058_, _14643_);
  or (_14645_, _14644_, _14642_);
  or (_14646_, _14479_, _07295_);
  and (_14647_, _14646_, _09154_);
  and (_14648_, _14647_, _14645_);
  or (_14649_, _14648_, _14473_);
  and (_14650_, _14649_, _07069_);
  or (_14651_, _09183_, _09182_);
  nor (_14652_, _09184_, _07069_);
  and (_14653_, _14652_, _14651_);
  or (_14654_, _14653_, _07067_);
  or (_14655_, _14654_, _14650_);
  nor (_14656_, _08177_, _08128_);
  nor (_14657_, _14656_, _08178_);
  or (_14658_, _14657_, _07232_);
  and (_14659_, _14658_, _07304_);
  and (_14660_, _14659_, _14655_);
  or (_14661_, _14660_, _14254_);
  and (_14662_, _14661_, _14470_);
  and (_14663_, _12043_, _06127_);
  not (_14664_, _11887_);
  nor (_14665_, _14664_, _06127_);
  or (_14666_, _14665_, _14663_);
  and (_14667_, _14666_, _14460_);
  and (_14668_, _14667_, _01336_);
  and (_14669_, _14668_, _42882_);
  and (_14670_, _14669_, _14459_);
  or (_40794_, _14670_, _14662_);
  and (_14671_, _14491_, _08029_);
  or (_14672_, _14671_, _08493_);
  or (_14673_, _14672_, _08797_);
  nor (_14674_, _14481_, _07353_);
  or (_14675_, _14674_, _08292_);
  or (_14676_, _14675_, _08286_);
  nor (_14677_, _08028_, _06215_);
  and (_14678_, _14677_, _08301_);
  nor (_14679_, _06148_, _05673_);
  nand (_14680_, _08028_, _06573_);
  nor (_14681_, _12666_, _07723_);
  or (_14682_, _14681_, _08378_);
  nand (_14683_, _12666_, _12644_);
  or (_14684_, _14683_, _08380_);
  and (_14685_, _14672_, _06955_);
  or (_14686_, _14675_, _08383_);
  and (_14687_, _06943_, _05853_);
  nor (_14688_, _06943_, _10010_);
  or (_14689_, _14688_, _14687_);
  nor (_14690_, _14689_, _08384_);
  nor (_14691_, _14690_, _06955_);
  and (_14692_, _14691_, _14686_);
  or (_14693_, _14692_, _06953_);
  or (_14694_, _14693_, _14685_);
  and (_14695_, _14694_, _14684_);
  or (_14696_, _14695_, _07272_);
  nor (_14697_, _05853_, _05690_);
  nor (_14698_, _14697_, _06963_);
  and (_14699_, _14698_, _14696_);
  and (_14700_, _09159_, _06963_);
  or (_14701_, _14700_, _06975_);
  or (_14702_, _14701_, _14699_);
  and (_14703_, _14702_, _14682_);
  or (_14704_, _14703_, _06038_);
  nand (_14705_, _08028_, _06038_);
  and (_14706_, _14705_, _06036_);
  and (_14707_, _14706_, _14704_);
  not (_14708_, _12667_);
  and (_14709_, _14683_, _14708_);
  and (_14710_, _14709_, _06035_);
  or (_14711_, _14710_, _14707_);
  and (_14712_, _14711_, _05686_);
  or (_14713_, _06148_, _05686_);
  nand (_14714_, _06233_, _14713_);
  or (_14715_, _14714_, _14712_);
  and (_14716_, _14715_, _14680_);
  or (_14717_, _14716_, _06992_);
  and (_14718_, _09181_, _06053_);
  nand (_14719_, _08026_, _06992_);
  or (_14720_, _14719_, _14718_);
  and (_14721_, _14720_, _14717_);
  or (_14722_, _14721_, _06991_);
  and (_14723_, _07723_, \oc8051_golden_model_1.PSW [7]);
  or (_14724_, _14681_, _14723_);
  or (_14725_, _14724_, _07308_);
  and (_14726_, _14725_, _05673_);
  and (_14727_, _14726_, _14722_);
  or (_14728_, _14727_, _14679_);
  and (_14729_, _14728_, _07009_);
  nor (_14730_, _07353_, _07009_);
  or (_14731_, _14730_, _07013_);
  or (_14732_, _14731_, _14729_);
  or (_14733_, _09181_, _07231_);
  and (_14734_, _14733_, _08545_);
  and (_14735_, _14734_, _14732_);
  nor (_14736_, _08549_, _07353_);
  and (_14737_, _08654_, \oc8051_golden_model_1.ACC [3]);
  and (_14738_, _08650_, \oc8051_golden_model_1.B [3]);
  or (_14739_, _14738_, _14737_);
  and (_14740_, _08660_, \oc8051_golden_model_1.P0 [3]);
  and (_14741_, _08704_, \oc8051_golden_model_1.PSW [3]);
  or (_14742_, _14741_, _14740_);
  or (_14743_, _14742_, _14739_);
  and (_14744_, _08680_, \oc8051_golden_model_1.TCON [3]);
  and (_14745_, _08682_, \oc8051_golden_model_1.P1 [3]);
  or (_14746_, _14745_, _14744_);
  and (_14747_, _08668_, \oc8051_golden_model_1.SCON [3]);
  and (_14748_, _08677_, \oc8051_golden_model_1.SBUF [3]);
  or (_14749_, _14748_, _14747_);
  or (_14750_, _14749_, _14746_);
  and (_14751_, _08687_, \oc8051_golden_model_1.P2 [3]);
  and (_14752_, _08690_, \oc8051_golden_model_1.IP [3]);
  or (_14753_, _14752_, _14751_);
  and (_14754_, _08693_, \oc8051_golden_model_1.IE [3]);
  and (_14755_, _08695_, \oc8051_golden_model_1.P3 [3]);
  or (_14756_, _14755_, _14754_);
  or (_14757_, _14756_, _14753_);
  and (_14758_, _08675_, \oc8051_golden_model_1.TMOD [3]);
  and (_14759_, _08702_, \oc8051_golden_model_1.TL0 [3]);
  or (_14760_, _14759_, _14758_);
  or (_14761_, _14760_, _14757_);
  or (_14762_, _14761_, _14750_);
  or (_14763_, _14762_, _14743_);
  and (_14764_, _08728_, \oc8051_golden_model_1.DPL [3]);
  and (_14765_, _08732_, \oc8051_golden_model_1.PCON [3]);
  and (_14766_, _08716_, \oc8051_golden_model_1.TL1 [3]);
  or (_14767_, _14766_, _14765_);
  or (_14768_, _14767_, _14764_);
  and (_14769_, _08725_, \oc8051_golden_model_1.TH1 [3]);
  and (_14770_, _08712_, \oc8051_golden_model_1.TH0 [3]);
  or (_14771_, _14770_, _14769_);
  and (_14772_, _08723_, \oc8051_golden_model_1.DPH [3]);
  and (_14773_, _08719_, \oc8051_golden_model_1.SP [3]);
  or (_14774_, _14773_, _14772_);
  or (_14775_, _14774_, _14771_);
  or (_14776_, _14775_, _14768_);
  or (_14777_, _14776_, _14763_);
  or (_14778_, _14777_, _14736_);
  and (_14779_, _14778_, _07010_);
  or (_14780_, _14779_, _08743_);
  or (_14781_, _14780_, _14735_);
  and (_14782_, _08743_, _05983_);
  nor (_14783_, _14782_, _06021_);
  and (_14784_, _14783_, _14781_);
  and (_14785_, _08662_, _06021_);
  or (_14786_, _14785_, _05724_);
  or (_14787_, _14786_, _14784_);
  and (_14788_, _06148_, _05724_);
  nor (_14789_, _14788_, _08752_);
  and (_14790_, _14789_, _14787_);
  not (_14791_, _14677_);
  nand (_14792_, _08028_, _06215_);
  and (_14793_, _14792_, _14791_);
  and (_14794_, _14793_, _08752_);
  or (_14795_, _14794_, _08757_);
  or (_14796_, _14795_, _14790_);
  or (_14797_, _12299_, _08765_);
  and (_14798_, _14797_, _08764_);
  and (_14799_, _14798_, _14796_);
  or (_14800_, _14799_, _14678_);
  and (_14801_, _14800_, _08300_);
  and (_14802_, _10987_, _07031_);
  or (_14803_, _14802_, _05736_);
  or (_14804_, _14803_, _14801_);
  and (_14805_, _06148_, _05736_);
  nor (_14806_, _14805_, _08778_);
  and (_14807_, _14806_, _14804_);
  and (_14808_, _14792_, _08778_);
  or (_14809_, _14808_, _08783_);
  or (_14810_, _14809_, _14807_);
  nand (_14811_, _10988_, _08783_);
  and (_14812_, _14811_, _05734_);
  and (_14813_, _14812_, _14810_);
  nand (_14814_, _05853_, _05732_);
  nand (_14815_, _08286_, _14814_);
  or (_14816_, _14815_, _14813_);
  and (_14817_, _14816_, _14676_);
  or (_14818_, _14817_, _07210_);
  or (_14819_, _14675_, _07211_);
  and (_14820_, _14819_, _07052_);
  and (_14821_, _14820_, _14818_);
  nor (_14822_, _09122_, _08985_);
  or (_14823_, _14822_, _09123_);
  and (_14824_, _14823_, _07051_);
  or (_14825_, _14824_, _07050_);
  or (_14826_, _14825_, _14821_);
  and (_14827_, _14826_, _14673_);
  or (_14828_, _14827_, _06127_);
  nand (_14829_, _12079_, _06127_);
  and (_14830_, _14829_, _12766_);
  and (_14831_, _14830_, _14828_);
  and (_14832_, _05853_, _05752_);
  or (_14833_, _07058_, _14832_);
  or (_14834_, _14833_, _14831_);
  or (_14835_, _14681_, _07295_);
  and (_14836_, _14835_, _09154_);
  and (_14837_, _14836_, _14834_);
  nor (_14838_, _09163_, _09159_);
  nor (_14839_, _14838_, _09164_);
  and (_14840_, _14839_, _14235_);
  or (_14841_, _14840_, _14837_);
  and (_14842_, _14841_, _07069_);
  or (_14843_, _09184_, _09181_);
  nor (_14844_, _09185_, _07069_);
  and (_14845_, _14844_, _14843_);
  or (_14846_, _14845_, _07067_);
  or (_14847_, _14846_, _14842_);
  nor (_14848_, _08178_, _08029_);
  nor (_14849_, _14848_, _08179_);
  or (_14850_, _14849_, _07232_);
  and (_14851_, _14850_, _07304_);
  and (_14852_, _14851_, _14847_);
  or (_14853_, _14852_, _14254_);
  or (_14854_, _14080_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_14855_, _14854_, _14073_);
  and (_14856_, _14855_, _14853_);
  and (_14857_, _11891_, _09200_);
  and (_14858_, _12036_, _06127_);
  or (_14859_, _14858_, _14857_);
  and (_14860_, _14859_, _14460_);
  and (_14861_, _14860_, _01336_);
  and (_14862_, _14861_, _42882_);
  and (_14863_, _14862_, _14459_);
  or (_40795_, _14863_, _14856_);
  or (_14864_, _14080_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_14865_, _14864_, _14073_);
  nor (_14866_, _09185_, _09180_);
  nor (_14867_, _14866_, _09186_);
  or (_14868_, _14867_, _07069_);
  and (_14869_, _08292_, _08270_);
  nor (_14870_, _08292_, _08270_);
  or (_14871_, _14870_, _14869_);
  or (_14872_, _14871_, _08286_);
  nand (_14873_, _08581_, _08272_);
  nor (_14874_, _08581_, _08272_);
  not (_14875_, _14874_);
  and (_14876_, _14875_, _14873_);
  and (_14877_, _14876_, _08752_);
  nand (_14878_, _12718_, _12716_);
  nand (_14879_, _12717_, _10606_);
  and (_14880_, _14879_, _06991_);
  and (_14881_, _14880_, _14878_);
  nor (_14882_, _12717_, _12716_);
  or (_14883_, _14882_, _08378_);
  or (_14884_, _14878_, _08380_);
  and (_14885_, _08493_, _08272_);
  nor (_14886_, _08493_, _08272_);
  or (_14887_, _14886_, _14885_);
  or (_14888_, _14887_, _08381_);
  and (_14889_, _09180_, _06948_);
  or (_14890_, _14871_, _08383_);
  nor (_14891_, _06943_, _09880_);
  and (_14892_, _11921_, _06943_);
  or (_14893_, _14892_, _14891_);
  or (_14894_, _14893_, _08384_);
  and (_14895_, _14894_, _06949_);
  and (_14896_, _14895_, _14890_);
  or (_14897_, _14896_, _06955_);
  or (_14898_, _14897_, _14889_);
  and (_14899_, _14898_, _14888_);
  or (_14900_, _14899_, _06953_);
  and (_14901_, _14900_, _14884_);
  or (_14902_, _14901_, _07272_);
  nor (_14903_, _11921_, _05690_);
  nor (_14904_, _14903_, _06963_);
  and (_14905_, _14904_, _14902_);
  and (_14906_, _09158_, _06963_);
  or (_14907_, _14906_, _06975_);
  or (_14908_, _14907_, _14905_);
  and (_14909_, _14908_, _14883_);
  or (_14910_, _14909_, _06038_);
  nand (_14911_, _08272_, _06038_);
  and (_14912_, _14911_, _06036_);
  and (_14913_, _14912_, _14910_);
  not (_14914_, _12719_);
  and (_14915_, _14878_, _14914_);
  and (_14916_, _14915_, _06035_);
  or (_14917_, _14916_, _14913_);
  and (_14918_, _14917_, _05686_);
  or (_14919_, _11922_, _05686_);
  nand (_14920_, _14919_, _06233_);
  or (_14921_, _14920_, _14918_);
  nand (_14922_, _08272_, _06573_);
  and (_14923_, _14922_, _14921_);
  or (_14924_, _14923_, _06992_);
  and (_14925_, _09180_, _06053_);
  nand (_14926_, _08225_, _06992_);
  or (_14927_, _14926_, _14925_);
  and (_14928_, _14927_, _07308_);
  and (_14929_, _14928_, _14924_);
  or (_14930_, _14929_, _14881_);
  and (_14931_, _14930_, _05673_);
  or (_14932_, _11922_, _05673_);
  nand (_14933_, _14932_, _07009_);
  or (_14934_, _14933_, _14931_);
  nand (_14935_, _08270_, _08541_);
  and (_14936_, _14935_, _14934_);
  or (_14937_, _14936_, _07013_);
  or (_14938_, _09180_, _07231_);
  and (_14939_, _14938_, _08545_);
  and (_14940_, _14939_, _14937_);
  nor (_14941_, _08549_, _08270_);
  and (_14942_, _08650_, \oc8051_golden_model_1.B [4]);
  and (_14943_, _08654_, \oc8051_golden_model_1.ACC [4]);
  or (_14944_, _14943_, _14942_);
  and (_14945_, _08702_, \oc8051_golden_model_1.TL0 [4]);
  and (_14946_, _08704_, \oc8051_golden_model_1.PSW [4]);
  or (_14947_, _14946_, _14945_);
  or (_14948_, _14947_, _14944_);
  and (_14949_, _08680_, \oc8051_golden_model_1.TCON [4]);
  and (_14950_, _08668_, \oc8051_golden_model_1.SCON [4]);
  or (_14951_, _14950_, _14949_);
  and (_14952_, _08660_, \oc8051_golden_model_1.P0 [4]);
  and (_14953_, _08677_, \oc8051_golden_model_1.SBUF [4]);
  or (_14954_, _14953_, _14952_);
  or (_14955_, _14954_, _14951_);
  and (_14956_, _08687_, \oc8051_golden_model_1.P2 [4]);
  and (_14957_, _08690_, \oc8051_golden_model_1.IP [4]);
  or (_14958_, _14957_, _14956_);
  and (_14959_, _08693_, \oc8051_golden_model_1.IE [4]);
  and (_14960_, _08695_, \oc8051_golden_model_1.P3 [4]);
  or (_14961_, _14960_, _14959_);
  or (_14962_, _14961_, _14958_);
  and (_14963_, _08675_, \oc8051_golden_model_1.TMOD [4]);
  and (_14964_, _08682_, \oc8051_golden_model_1.P1 [4]);
  or (_14965_, _14964_, _14963_);
  or (_14966_, _14965_, _14962_);
  or (_14967_, _14966_, _14955_);
  or (_14968_, _14967_, _14948_);
  and (_14969_, _08728_, \oc8051_golden_model_1.DPL [4]);
  and (_14970_, _08719_, \oc8051_golden_model_1.SP [4]);
  and (_14971_, _08723_, \oc8051_golden_model_1.DPH [4]);
  or (_14972_, _14971_, _14970_);
  or (_14973_, _14972_, _14969_);
  and (_14974_, _08716_, \oc8051_golden_model_1.TL1 [4]);
  and (_14975_, _08725_, \oc8051_golden_model_1.TH1 [4]);
  or (_14976_, _14975_, _14974_);
  and (_14977_, _08732_, \oc8051_golden_model_1.PCON [4]);
  and (_14978_, _08712_, \oc8051_golden_model_1.TH0 [4]);
  or (_14979_, _14978_, _14977_);
  or (_14980_, _14979_, _14976_);
  or (_14981_, _14980_, _14973_);
  or (_14982_, _14981_, _14968_);
  or (_14983_, _14982_, _14941_);
  and (_14984_, _14983_, _07010_);
  or (_14985_, _14984_, _08743_);
  or (_14986_, _14985_, _14940_);
  and (_14987_, _08743_, _06758_);
  nor (_14988_, _14987_, _06021_);
  and (_14989_, _14988_, _14986_);
  and (_14990_, _08665_, _06021_);
  or (_14991_, _14990_, _05724_);
  or (_14992_, _14991_, _14989_);
  and (_14993_, _11922_, _05724_);
  nor (_14994_, _14993_, _08752_);
  and (_14995_, _14994_, _14992_);
  or (_14996_, _14995_, _14877_);
  and (_14997_, _14996_, _08765_);
  and (_14998_, _10986_, _08757_);
  or (_14999_, _14998_, _14997_);
  and (_15000_, _14999_, _08764_);
  and (_15001_, _14874_, _08301_);
  or (_15002_, _15001_, _15000_);
  and (_15003_, _15002_, _08300_);
  and (_15004_, _10983_, _07031_);
  or (_15005_, _15004_, _05736_);
  or (_15006_, _15005_, _15003_);
  and (_15007_, _11922_, _05736_);
  nor (_15008_, _15007_, _08778_);
  and (_15009_, _15008_, _15006_);
  and (_15010_, _14873_, _08778_);
  or (_15011_, _15010_, _08783_);
  or (_15012_, _15011_, _15009_);
  nand (_15013_, _10985_, _08783_);
  and (_15014_, _15013_, _05734_);
  and (_15015_, _15014_, _15012_);
  nand (_15016_, _11921_, _05732_);
  nand (_15017_, _15016_, _08286_);
  or (_15018_, _15017_, _15015_);
  and (_15019_, _15018_, _14872_);
  or (_15020_, _15019_, _07210_);
  and (_15021_, _10394_, _05495_);
  not (_15022_, _15021_);
  or (_15023_, _14871_, _07211_);
  and (_15024_, _15023_, _15022_);
  and (_15025_, _15024_, _15020_);
  nor (_15026_, _09123_, _08937_);
  or (_15027_, _15026_, _09124_);
  or (_15028_, _15027_, _06712_);
  and (_15029_, _15028_, _07051_);
  or (_15030_, _15029_, _15025_);
  not (_15031_, _06712_);
  or (_15032_, _15027_, _15031_);
  and (_15033_, _15032_, _08797_);
  and (_15034_, _15033_, _15030_);
  and (_15035_, _14887_, _07050_);
  or (_15036_, _15035_, _06127_);
  or (_15037_, _15036_, _15034_);
  nand (_15038_, _12075_, _06127_);
  and (_15039_, _15038_, _12766_);
  and (_15040_, _15039_, _15037_);
  and (_15041_, _11921_, _05752_);
  or (_15042_, _15041_, _07058_);
  or (_15043_, _15042_, _15040_);
  or (_15044_, _14882_, _07295_);
  and (_15045_, _15044_, _09154_);
  and (_15046_, _15045_, _15043_);
  nor (_15047_, _09164_, _09158_);
  nor (_15048_, _15047_, _09165_);
  and (_15049_, _15048_, _14235_);
  or (_15050_, _15049_, _07068_);
  or (_15051_, _15050_, _15046_);
  and (_15052_, _15051_, _14868_);
  or (_15053_, _15052_, _07067_);
  nor (_15054_, _08273_, _08179_);
  nor (_15055_, _15054_, _08274_);
  or (_15056_, _15055_, _07232_);
  and (_15057_, _15056_, _07304_);
  and (_15058_, _15057_, _15053_);
  or (_15059_, _15058_, _14254_);
  and (_15060_, _15059_, _14865_);
  and (_15061_, _12032_, _06127_);
  not (_15062_, _11884_);
  nor (_15063_, _15062_, _06127_);
  or (_15064_, _15063_, _15061_);
  and (_15065_, _15064_, _14460_);
  and (_15066_, _15065_, _01336_);
  and (_15067_, _15066_, _42882_);
  and (_15068_, _15067_, _14459_);
  or (_40797_, _15068_, _15060_);
  or (_15069_, _14080_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_15070_, _15069_, _14073_);
  nor (_15071_, _08612_, _07979_);
  and (_15072_, _15071_, _08301_);
  nand (_15073_, _12640_, _12638_);
  nand (_15074_, _12639_, _10606_);
  and (_15075_, _15074_, _06991_);
  and (_15076_, _15075_, _15073_);
  nor (_15077_, _12639_, _12638_);
  or (_15078_, _15077_, _08378_);
  or (_15079_, _15073_, _08380_);
  or (_15080_, _09179_, _06949_);
  nor (_15081_, _14869_, _07977_);
  or (_15082_, _15081_, _08293_);
  and (_15083_, _15082_, _08384_);
  nand (_15084_, _11917_, _06943_);
  or (_15085_, _06943_, \oc8051_golden_model_1.ACC [5]);
  and (_15086_, _15085_, _15084_);
  and (_15087_, _15086_, _08383_);
  or (_15088_, _15087_, _06948_);
  or (_15089_, _15088_, _15083_);
  and (_15090_, _15089_, _15080_);
  or (_15091_, _15090_, _06955_);
  nor (_15092_, _14885_, _07979_);
  or (_15093_, _15092_, _08494_);
  or (_15094_, _15093_, _08381_);
  and (_15095_, _15094_, _15091_);
  or (_15096_, _15095_, _06953_);
  and (_15097_, _15096_, _15079_);
  or (_15098_, _15097_, _07272_);
  nor (_15099_, _11916_, _05690_);
  nor (_15100_, _15099_, _06963_);
  and (_15101_, _15100_, _15098_);
  and (_15102_, _09157_, _06963_);
  or (_15103_, _15102_, _06975_);
  or (_15104_, _15103_, _15101_);
  and (_15105_, _15104_, _15078_);
  or (_15106_, _15105_, _06038_);
  nand (_15107_, _07979_, _06038_);
  and (_15108_, _15107_, _06036_);
  and (_15109_, _15108_, _15106_);
  not (_15110_, _12641_);
  and (_15111_, _15073_, _15110_);
  and (_15112_, _15111_, _06035_);
  or (_15113_, _15112_, _15109_);
  and (_15114_, _15113_, _05686_);
  or (_15115_, _11917_, _05686_);
  nand (_15116_, _15115_, _06233_);
  or (_15117_, _15116_, _15114_);
  nand (_15118_, _07979_, _06573_);
  and (_15119_, _15118_, _15117_);
  or (_15120_, _15119_, _06992_);
  and (_15121_, _09179_, _06053_);
  nand (_15122_, _07932_, _06992_);
  or (_15123_, _15122_, _15121_);
  and (_15124_, _15123_, _07308_);
  and (_15125_, _15124_, _15120_);
  or (_15126_, _15125_, _15076_);
  and (_15127_, _15126_, _05673_);
  or (_15128_, _11917_, _05673_);
  nand (_15129_, _15128_, _07009_);
  or (_15130_, _15129_, _15127_);
  nand (_15131_, _07977_, _08541_);
  and (_15132_, _15131_, _15130_);
  or (_15133_, _15132_, _07013_);
  or (_15134_, _09179_, _07231_);
  and (_15135_, _15134_, _08545_);
  and (_15136_, _15135_, _15133_);
  nor (_15137_, _08549_, _07977_);
  and (_15138_, _08675_, \oc8051_golden_model_1.TMOD [5]);
  and (_15139_, _08668_, \oc8051_golden_model_1.SCON [5]);
  or (_15140_, _15139_, _15138_);
  and (_15141_, _08702_, \oc8051_golden_model_1.TL0 [5]);
  and (_15142_, _08650_, \oc8051_golden_model_1.B [5]);
  or (_15143_, _15142_, _15141_);
  or (_15144_, _15143_, _15140_);
  and (_15145_, _08660_, \oc8051_golden_model_1.P0 [5]);
  and (_15146_, _08680_, \oc8051_golden_model_1.TCON [5]);
  or (_15147_, _15146_, _15145_);
  and (_15148_, _08682_, \oc8051_golden_model_1.P1 [5]);
  and (_15149_, _08704_, \oc8051_golden_model_1.PSW [5]);
  or (_15150_, _15149_, _15148_);
  or (_15151_, _15150_, _15147_);
  and (_15152_, _08693_, \oc8051_golden_model_1.IE [5]);
  and (_15153_, _08690_, \oc8051_golden_model_1.IP [5]);
  or (_15154_, _15153_, _15152_);
  and (_15155_, _08687_, \oc8051_golden_model_1.P2 [5]);
  and (_15156_, _08695_, \oc8051_golden_model_1.P3 [5]);
  or (_15157_, _15156_, _15155_);
  or (_15158_, _15157_, _15154_);
  and (_15159_, _08677_, \oc8051_golden_model_1.SBUF [5]);
  and (_15160_, _08654_, \oc8051_golden_model_1.ACC [5]);
  or (_15161_, _15160_, _15159_);
  or (_15162_, _15161_, _15158_);
  or (_15163_, _15162_, _15151_);
  or (_15164_, _15163_, _15144_);
  and (_15165_, _08712_, \oc8051_golden_model_1.TH0 [5]);
  and (_15166_, _08723_, \oc8051_golden_model_1.DPH [5]);
  and (_15167_, _08725_, \oc8051_golden_model_1.TH1 [5]);
  or (_15168_, _15167_, _15166_);
  or (_15169_, _15168_, _15165_);
  and (_15170_, _08732_, \oc8051_golden_model_1.PCON [5]);
  and (_15171_, _08716_, \oc8051_golden_model_1.TL1 [5]);
  or (_15172_, _15171_, _15170_);
  and (_15173_, _08728_, \oc8051_golden_model_1.DPL [5]);
  and (_15174_, _08719_, \oc8051_golden_model_1.SP [5]);
  or (_15175_, _15174_, _15173_);
  or (_15176_, _15175_, _15172_);
  or (_15177_, _15176_, _15169_);
  or (_15178_, _15177_, _15164_);
  or (_15179_, _15178_, _15137_);
  and (_15180_, _15179_, _07010_);
  or (_15181_, _15180_, _08743_);
  or (_15182_, _15181_, _15136_);
  and (_15183_, _08743_, _06359_);
  nor (_15184_, _15183_, _06021_);
  and (_15185_, _15184_, _15182_);
  and (_15186_, _08652_, _06021_);
  or (_15187_, _15186_, _05724_);
  or (_15188_, _15187_, _15185_);
  and (_15189_, _11917_, _05724_);
  nor (_15190_, _15189_, _08752_);
  and (_15191_, _15190_, _15188_);
  not (_15192_, _15071_);
  nand (_15194_, _08612_, _07979_);
  and (_15195_, _15194_, _15192_);
  and (_15196_, _15195_, _08752_);
  or (_15197_, _15196_, _08757_);
  or (_15198_, _15197_, _15191_);
  or (_15199_, _12306_, _08765_);
  and (_15200_, _15199_, _08764_);
  and (_15201_, _15200_, _15198_);
  or (_15202_, _15201_, _15072_);
  and (_15203_, _15202_, _08300_);
  and (_15204_, _10981_, _07031_);
  or (_15205_, _15204_, _05736_);
  or (_15206_, _15205_, _15203_);
  and (_15207_, _11917_, _05736_);
  nor (_15208_, _15207_, _08778_);
  and (_15209_, _15208_, _15206_);
  and (_15210_, _15194_, _08778_);
  or (_15211_, _15210_, _08783_);
  or (_15212_, _15211_, _15209_);
  nand (_15213_, _10982_, _08783_);
  and (_15214_, _15213_, _05734_);
  and (_15215_, _15214_, _15212_);
  nand (_15216_, _11916_, _05732_);
  nand (_15217_, _15216_, _08287_);
  or (_15218_, _15217_, _15215_);
  or (_15219_, _15082_, _08287_);
  and (_15220_, _15219_, _15022_);
  and (_15221_, _15220_, _15218_);
  nor (_15222_, _09124_, _08888_);
  or (_15223_, _15222_, _09125_);
  or (_15224_, _15223_, _06712_);
  and (_15225_, _15224_, _07051_);
  or (_15226_, _15225_, _15221_);
  or (_15227_, _15223_, _15031_);
  and (_15228_, _15227_, _08797_);
  and (_15229_, _15228_, _15226_);
  and (_15230_, _15093_, _07050_);
  or (_15231_, _15230_, _06127_);
  or (_15232_, _15231_, _15229_);
  nand (_15233_, _12070_, _06127_);
  and (_15234_, _15233_, _12766_);
  and (_15235_, _15234_, _15232_);
  and (_15236_, _11916_, _05752_);
  or (_15237_, _15236_, _07058_);
  or (_15238_, _15237_, _15235_);
  or (_15239_, _15077_, _07295_);
  and (_15240_, _15239_, _09154_);
  and (_15241_, _15240_, _15238_);
  or (_15242_, _09165_, _09157_);
  nor (_15243_, _09166_, _09154_);
  and (_15244_, _15243_, _15242_);
  or (_15245_, _15244_, _15241_);
  and (_15246_, _15245_, _07069_);
  or (_15247_, _09186_, _09179_);
  nor (_15248_, _09187_, _07069_);
  and (_15249_, _15248_, _15247_);
  or (_15250_, _15249_, _07067_);
  or (_15251_, _15250_, _15246_);
  nor (_15252_, _08274_, _07980_);
  nor (_15253_, _15252_, _08275_);
  or (_15254_, _15253_, _07232_);
  and (_15255_, _15254_, _07304_);
  and (_15256_, _15255_, _15251_);
  or (_15257_, _15256_, _14254_);
  and (_15258_, _15257_, _15070_);
  not (_15259_, _11880_);
  nor (_15260_, _15259_, _06127_);
  and (_15261_, _12027_, _06127_);
  or (_15262_, _15261_, _15260_);
  and (_15263_, _15262_, _14460_);
  and (_15264_, _15263_, _01336_);
  and (_15265_, _15264_, _42882_);
  and (_15266_, _15265_, _14459_);
  or (_40798_, _15266_, _15258_);
  or (_15267_, _14080_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_15268_, _15267_, _14073_);
  nor (_15269_, _09166_, _09156_);
  nor (_15270_, _15269_, _09167_);
  and (_15271_, _15270_, _14235_);
  nor (_15272_, _09125_, _08843_);
  or (_15273_, _15272_, _09126_);
  and (_15274_, _15273_, _07051_);
  nor (_15275_, _08293_, _07883_);
  or (_15276_, _15275_, _08294_);
  or (_15277_, _15276_, _08286_);
  nor (_15278_, _12691_, _12690_);
  or (_15279_, _15278_, _08378_);
  nand (_15280_, _12692_, _12690_);
  or (_15281_, _15280_, _08380_);
  or (_15282_, _09178_, _06949_);
  and (_15283_, _15276_, _08384_);
  nand (_15284_, _11909_, _06943_);
  or (_15285_, _06943_, \oc8051_golden_model_1.ACC [6]);
  and (_15286_, _15285_, _15284_);
  and (_15287_, _15286_, _08383_);
  or (_15288_, _15287_, _06948_);
  or (_15289_, _15288_, _15283_);
  and (_15290_, _15289_, _15282_);
  or (_15291_, _15290_, _06955_);
  nor (_15292_, _08494_, _07885_);
  or (_15293_, _15292_, _08495_);
  or (_15294_, _15293_, _08381_);
  and (_15295_, _15294_, _15291_);
  or (_15296_, _15295_, _06953_);
  and (_15297_, _15296_, _15281_);
  or (_15298_, _15297_, _07272_);
  nor (_15299_, _11908_, _05690_);
  nor (_15300_, _15299_, _06963_);
  and (_15301_, _15300_, _15298_);
  and (_15302_, _09156_, _06963_);
  or (_15303_, _15302_, _06975_);
  or (_15304_, _15303_, _15301_);
  and (_15305_, _15304_, _15279_);
  or (_15306_, _15305_, _06038_);
  nand (_15307_, _07885_, _06038_);
  and (_15308_, _15307_, _06036_);
  and (_15309_, _15308_, _15306_);
  not (_15310_, _12693_);
  and (_15311_, _15280_, _15310_);
  and (_15312_, _15311_, _06035_);
  or (_15313_, _15312_, _15309_);
  and (_15314_, _15313_, _05686_);
  or (_15315_, _11909_, _05686_);
  nand (_15316_, _15315_, _06233_);
  or (_15317_, _15316_, _15314_);
  nand (_15318_, _07885_, _06573_);
  and (_15319_, _15318_, _15317_);
  or (_15320_, _15319_, _06992_);
  and (_15321_, _09178_, _06053_);
  nand (_15322_, _07838_, _06992_);
  or (_15323_, _15322_, _15321_);
  and (_15324_, _15323_, _07308_);
  and (_15325_, _15324_, _15320_);
  nand (_15326_, _12691_, _10606_);
  and (_15327_, _15326_, _06991_);
  and (_15328_, _15327_, _15280_);
  or (_15329_, _15328_, _15325_);
  and (_15330_, _15329_, _05673_);
  or (_15331_, _11909_, _05673_);
  nand (_15332_, _15331_, _07009_);
  or (_15333_, _15332_, _15330_);
  nand (_15334_, _07883_, _08541_);
  and (_15335_, _15334_, _15333_);
  or (_15336_, _15335_, _07013_);
  or (_15337_, _09178_, _07231_);
  and (_15338_, _15337_, _08545_);
  and (_15339_, _15338_, _15336_);
  nor (_15340_, _08549_, _07883_);
  and (_15341_, _08654_, \oc8051_golden_model_1.ACC [6]);
  and (_15342_, _08650_, \oc8051_golden_model_1.B [6]);
  or (_15343_, _15342_, _15341_);
  and (_15344_, _08702_, \oc8051_golden_model_1.TL0 [6]);
  and (_15345_, _08677_, \oc8051_golden_model_1.SBUF [6]);
  or (_15346_, _15345_, _15344_);
  or (_15347_, _15346_, _15343_);
  and (_15348_, _08660_, \oc8051_golden_model_1.P0 [6]);
  and (_15349_, _08675_, \oc8051_golden_model_1.TMOD [6]);
  or (_15350_, _15349_, _15348_);
  and (_15351_, _08682_, \oc8051_golden_model_1.P1 [6]);
  and (_15352_, _08668_, \oc8051_golden_model_1.SCON [6]);
  or (_15353_, _15352_, _15351_);
  or (_15354_, _15353_, _15350_);
  and (_15355_, _08695_, \oc8051_golden_model_1.P3 [6]);
  and (_15356_, _08690_, \oc8051_golden_model_1.IP [6]);
  or (_15357_, _15356_, _15355_);
  and (_15358_, _08687_, \oc8051_golden_model_1.P2 [6]);
  and (_15359_, _08693_, \oc8051_golden_model_1.IE [6]);
  or (_15360_, _15359_, _15358_);
  or (_15361_, _15360_, _15357_);
  and (_15362_, _08680_, \oc8051_golden_model_1.TCON [6]);
  and (_15363_, _08704_, \oc8051_golden_model_1.PSW [6]);
  or (_15364_, _15363_, _15362_);
  or (_15365_, _15364_, _15361_);
  or (_15366_, _15365_, _15354_);
  or (_15367_, _15366_, _15347_);
  and (_15368_, _08716_, \oc8051_golden_model_1.TL1 [6]);
  and (_15369_, _08728_, \oc8051_golden_model_1.DPL [6]);
  and (_15370_, _08723_, \oc8051_golden_model_1.DPH [6]);
  or (_15371_, _15370_, _15369_);
  or (_15372_, _15371_, _15368_);
  and (_15373_, _08712_, \oc8051_golden_model_1.TH0 [6]);
  and (_15374_, _08725_, \oc8051_golden_model_1.TH1 [6]);
  or (_15375_, _15374_, _15373_);
  and (_15376_, _08732_, \oc8051_golden_model_1.PCON [6]);
  and (_15377_, _08719_, \oc8051_golden_model_1.SP [6]);
  or (_15378_, _15377_, _15376_);
  or (_15379_, _15378_, _15375_);
  or (_15380_, _15379_, _15372_);
  or (_15381_, _15380_, _15367_);
  or (_15382_, _15381_, _15340_);
  and (_15383_, _15382_, _07010_);
  or (_15384_, _15383_, _08743_);
  or (_15385_, _15384_, _15339_);
  and (_15386_, _08743_, _06084_);
  nor (_15387_, _15386_, _06021_);
  and (_15388_, _15387_, _15385_);
  not (_15389_, _08647_);
  and (_15390_, _15389_, _06021_);
  or (_15391_, _15390_, _05724_);
  or (_15392_, _15391_, _15388_);
  and (_15393_, _11909_, _05724_);
  nor (_15394_, _15393_, _08752_);
  and (_15395_, _15394_, _15392_);
  nand (_15396_, _08647_, _07885_);
  nor (_15397_, _08647_, _07885_);
  not (_15398_, _15397_);
  and (_15399_, _15398_, _15396_);
  and (_15400_, _15399_, _08752_);
  or (_15401_, _15400_, _15395_);
  and (_15402_, _15401_, _08765_);
  and (_15403_, _10980_, _08757_);
  or (_15404_, _15403_, _15402_);
  and (_15405_, _15404_, _08764_);
  and (_15406_, _15397_, _08301_);
  or (_15407_, _15406_, _15405_);
  and (_15408_, _15407_, _08300_);
  and (_15409_, _10977_, _07031_);
  or (_15410_, _15409_, _05736_);
  or (_15411_, _15410_, _15408_);
  and (_15412_, _11909_, _05736_);
  nor (_15413_, _15412_, _08778_);
  and (_15414_, _15413_, _15411_);
  and (_15415_, _15396_, _08778_);
  or (_15416_, _15415_, _08783_);
  or (_15417_, _15416_, _15414_);
  nand (_15418_, _10979_, _08783_);
  and (_15419_, _15418_, _05734_);
  and (_15420_, _15419_, _15417_);
  nand (_15421_, _11908_, _05732_);
  nand (_15422_, _15421_, _08286_);
  or (_15423_, _15422_, _15420_);
  and (_15424_, _15423_, _15277_);
  or (_15425_, _15424_, _07210_);
  or (_15426_, _15276_, _07211_);
  and (_15427_, _15426_, _07052_);
  and (_15428_, _15427_, _15425_);
  or (_15429_, _15428_, _15274_);
  and (_15430_, _15429_, _08797_);
  and (_15431_, _15293_, _07050_);
  or (_15432_, _15431_, _06127_);
  or (_15433_, _15432_, _15430_);
  nand (_15434_, _12063_, _06127_);
  and (_15435_, _15434_, _12766_);
  and (_15436_, _15435_, _15433_);
  and (_15437_, _11908_, _05752_);
  or (_15438_, _15437_, _07058_);
  or (_15439_, _15438_, _15436_);
  or (_15440_, _15278_, _07295_);
  and (_15441_, _15440_, _09154_);
  and (_15442_, _15441_, _15439_);
  or (_15443_, _15442_, _15271_);
  and (_15444_, _15443_, _07069_);
  or (_15445_, _09187_, _09178_);
  nor (_15446_, _09188_, _07069_);
  and (_15447_, _15446_, _15445_);
  or (_15448_, _15447_, _07067_);
  or (_15449_, _15448_, _15444_);
  nor (_15450_, _08275_, _07886_);
  nor (_15451_, _15450_, _08276_);
  or (_15452_, _15451_, _07232_);
  and (_15453_, _15452_, _07304_);
  and (_15454_, _15453_, _15449_);
  or (_15455_, _15454_, _14254_);
  and (_15456_, _15455_, _15268_);
  not (_15457_, _11875_);
  nor (_15458_, _15457_, _06127_);
  and (_15459_, _12020_, _06127_);
  or (_15460_, _15459_, _15458_);
  and (_15461_, _15460_, _14460_);
  and (_15462_, _15461_, _01336_);
  and (_15463_, _15462_, _42882_);
  and (_15464_, _15463_, _14459_);
  or (_40799_, _15464_, _15456_);
  nand (_15465_, _14080_, _09196_);
  or (_15466_, _14080_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_15467_, _15466_, _14073_);
  and (_15468_, _15467_, _15465_);
  and (_15469_, _14072_, _09229_);
  or (_40800_, _15469_, _15468_);
  nand (_15470_, _14071_, _07356_);
  or (_15471_, _15470_, _14068_);
  and (_15472_, _14077_, _07229_);
  and (_15473_, _15472_, _14076_);
  and (_15474_, _15473_, _14247_);
  or (_15475_, _15473_, _06880_);
  nand (_15476_, _15475_, _15470_);
  or (_15477_, _15476_, _15474_);
  and (_40801_, _15477_, _15471_);
  not (_15478_, _15473_);
  or (_15479_, _15478_, _14436_);
  or (_15480_, _15473_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_15481_, _15480_, _15470_);
  and (_15482_, _15481_, _15479_);
  and (_15483_, _14447_, _14443_);
  and (_15484_, _15483_, _14457_);
  and (_15485_, _15484_, _14467_);
  or (_40802_, _15485_, _15482_);
  or (_15486_, _15478_, _14660_);
  or (_15487_, _15473_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_15488_, _15487_, _15470_);
  and (_15489_, _15488_, _15486_);
  and (_15490_, _15484_, _14669_);
  or (_40803_, _15490_, _15489_);
  or (_15491_, _15478_, _14852_);
  or (_15492_, _15473_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_15493_, _15492_, _15470_);
  and (_15494_, _15493_, _15491_);
  and (_15495_, _15484_, _14862_);
  or (_40805_, _15495_, _15494_);
  or (_15496_, _15478_, _15058_);
  or (_15497_, _15473_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_15498_, _15497_, _15470_);
  and (_15499_, _15498_, _15496_);
  and (_15500_, _15484_, _15067_);
  or (_40806_, _15500_, _15499_);
  or (_15501_, _15478_, _15256_);
  or (_15502_, _15473_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_15503_, _15502_, _15470_);
  and (_15504_, _15503_, _15501_);
  and (_15505_, _15484_, _15265_);
  or (_40807_, _15505_, _15504_);
  or (_15506_, _15478_, _15454_);
  or (_15507_, _15473_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_15508_, _15507_, _15470_);
  and (_15509_, _15508_, _15506_);
  and (_15510_, _15484_, _15463_);
  or (_40808_, _15510_, _15509_);
  and (_15511_, _15473_, _09197_);
  or (_15512_, _15473_, _07740_);
  nand (_15513_, _15512_, _15470_);
  or (_15514_, _15513_, _15511_);
  or (_15515_, _15470_, _09229_);
  and (_40809_, _15515_, _15514_);
  and (_15516_, _14068_, _07628_);
  and (_15517_, _14071_, _08399_);
  not (_15518_, _15517_);
  or (_15519_, _15518_, _15516_);
  and (_15520_, _07306_, _07074_);
  and (_15521_, _15520_, _14076_);
  and (_15522_, _15521_, _14247_);
  nor (_15523_, _15521_, _06888_);
  or (_15524_, _15523_, _15517_);
  or (_15525_, _15524_, _15522_);
  and (_40813_, _15525_, _15519_);
  not (_15526_, _15521_);
  or (_15527_, _15526_, _14436_);
  or (_15528_, _15521_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_15529_, _15528_, _15518_);
  and (_15530_, _15529_, _15527_);
  and (_15531_, _14464_, _07628_);
  and (_15532_, _15531_, _15517_);
  or (_40814_, _15532_, _15530_);
  or (_15533_, _15526_, _14660_);
  or (_15534_, _15521_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_15535_, _15534_, _15518_);
  and (_15536_, _15535_, _15533_);
  and (_15537_, _14666_, _07628_);
  and (_15538_, _15537_, _15517_);
  or (_40815_, _15538_, _15536_);
  or (_15539_, _15526_, _14852_);
  or (_15540_, _15521_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_15541_, _15540_, _15518_);
  and (_15542_, _15541_, _15539_);
  and (_15543_, _14859_, _07628_);
  and (_15544_, _15543_, _15517_);
  or (_40816_, _15544_, _15542_);
  or (_15545_, _15526_, _15058_);
  or (_15546_, _15521_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_15547_, _15546_, _15518_);
  and (_15548_, _15547_, _15545_);
  and (_15549_, _15064_, _07628_);
  and (_15550_, _15549_, _15517_);
  or (_40818_, _15550_, _15548_);
  or (_15551_, _15526_, _15256_);
  or (_15552_, _15521_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_15553_, _15552_, _15518_);
  and (_15554_, _15553_, _15551_);
  and (_15555_, _15262_, _07628_);
  and (_15556_, _15555_, _15517_);
  or (_40819_, _15556_, _15554_);
  or (_15557_, _15526_, _15454_);
  or (_15558_, _15521_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_15559_, _15558_, _15518_);
  and (_15560_, _15559_, _15557_);
  and (_15561_, _15460_, _07628_);
  and (_15562_, _15561_, _15517_);
  or (_40820_, _15562_, _15560_);
  or (_15563_, _15526_, _09197_);
  or (_15564_, _15521_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_15565_, _15564_, _15518_);
  and (_15566_, _15565_, _15563_);
  and (_15567_, _15517_, _09230_);
  or (_40821_, _15567_, _15566_);
  and (_15568_, _14071_, _07080_);
  not (_15569_, _15568_);
  or (_15570_, _15569_, _15516_);
  and (_15571_, _14076_, _07307_);
  and (_15572_, _15571_, _14247_);
  nor (_15573_, _15571_, _06885_);
  or (_15574_, _15573_, _15568_);
  or (_15575_, _15574_, _15572_);
  and (_40823_, _15575_, _15570_);
  or (_15576_, _15571_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_15577_, _15576_, _15569_);
  not (_15578_, _15571_);
  or (_15579_, _15578_, _14436_);
  and (_15580_, _15579_, _15577_);
  and (_15581_, _15568_, _15531_);
  or (_40824_, _15581_, _15580_);
  or (_15582_, _15571_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_15583_, _15582_, _15569_);
  or (_15584_, _15578_, _14660_);
  and (_15585_, _15584_, _15583_);
  and (_15586_, _15568_, _15537_);
  or (_40825_, _15586_, _15585_);
  or (_15587_, _15571_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_15588_, _15587_, _15569_);
  or (_15589_, _15578_, _14852_);
  and (_15590_, _15589_, _15588_);
  and (_15591_, _15568_, _15543_);
  or (_40827_, _15591_, _15590_);
  or (_15592_, _15571_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_15593_, _15592_, _15569_);
  or (_15594_, _15578_, _15058_);
  and (_15595_, _15594_, _15593_);
  and (_15596_, _15568_, _15549_);
  or (_40828_, _15596_, _15595_);
  or (_15597_, _15571_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_15598_, _15597_, _15569_);
  or (_15599_, _15578_, _15256_);
  and (_15600_, _15599_, _15598_);
  and (_15601_, _15568_, _15555_);
  or (_40829_, _15601_, _15600_);
  or (_15602_, _15571_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_15603_, _15602_, _15569_);
  or (_15604_, _15578_, _15454_);
  and (_15605_, _15604_, _15603_);
  and (_15606_, _15568_, _15561_);
  or (_40830_, _15606_, _15605_);
  or (_15607_, _15571_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_15608_, _15607_, _15569_);
  or (_15609_, _15578_, _09197_);
  and (_15610_, _15609_, _15608_);
  and (_15611_, _15568_, _09230_);
  or (_40831_, _15611_, _15610_);
  and (_15612_, _07628_, _07622_);
  and (_15613_, _15612_, _14453_);
  and (_15614_, _15613_, _07081_);
  not (_15615_, _15614_);
  and (_15616_, _07615_, _07476_);
  and (_15617_, _15616_, _14078_);
  or (_15618_, _15617_, \oc8051_golden_model_1.IRAM[4] [0]);
  not (_15619_, _15617_);
  or (_15620_, _15619_, _14247_);
  and (_15621_, _15620_, _15618_);
  and (_15622_, _15621_, _15615_);
  and (_15623_, _15614_, _15516_);
  or (_40835_, _15623_, _15622_);
  or (_15624_, _15619_, _14436_);
  or (_15625_, _15617_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_15626_, _15625_, _15615_);
  and (_15627_, _15626_, _15624_);
  and (_15628_, _15614_, _15531_);
  or (_40836_, _15628_, _15627_);
  or (_15629_, _15619_, _14660_);
  or (_15630_, _15617_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_15631_, _15630_, _15615_);
  and (_15632_, _15631_, _15629_);
  and (_15633_, _15614_, _15537_);
  or (_40837_, _15633_, _15632_);
  or (_15634_, _15619_, _14852_);
  or (_15635_, _15617_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_15636_, _15635_, _15615_);
  and (_15637_, _15636_, _15634_);
  and (_15638_, _15614_, _15543_);
  or (_40838_, _15638_, _15637_);
  or (_15639_, _15619_, _15058_);
  or (_15640_, _15617_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_15641_, _15640_, _15615_);
  and (_15642_, _15641_, _15639_);
  and (_15643_, _15614_, _15549_);
  or (_40841_, _15643_, _15642_);
  or (_15644_, _15619_, _15256_);
  or (_15645_, _15617_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_15646_, _15645_, _15615_);
  and (_15647_, _15646_, _15644_);
  and (_15648_, _15614_, _15555_);
  or (_40842_, _15648_, _15647_);
  or (_15649_, _15619_, _15454_);
  or (_15650_, _15617_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_15651_, _15650_, _15615_);
  and (_15652_, _15651_, _15649_);
  and (_15653_, _15614_, _15561_);
  or (_40843_, _15653_, _15652_);
  or (_15654_, _15619_, _09197_);
  or (_15655_, _15617_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_15656_, _15655_, _15615_);
  and (_15657_, _15656_, _15654_);
  and (_15658_, _15614_, _09230_);
  or (_40844_, _15658_, _15657_);
  and (_15659_, _15616_, _15472_);
  not (_15660_, _15659_);
  or (_15661_, _15660_, _14247_);
  and (_15662_, _15613_, _07356_);
  not (_15663_, _15662_);
  or (_15664_, _15659_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_15665_, _15664_, _15663_);
  and (_15666_, _15665_, _15661_);
  and (_15667_, _15662_, _15516_);
  or (_40848_, _15667_, _15666_);
  or (_15668_, _15660_, _14436_);
  or (_15669_, _15659_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_15670_, _15669_, _15663_);
  and (_15671_, _15670_, _15668_);
  and (_15672_, _15662_, _15531_);
  or (_40849_, _15672_, _15671_);
  or (_15673_, _15660_, _14660_);
  or (_15674_, _15659_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_15675_, _15674_, _15663_);
  and (_15676_, _15675_, _15673_);
  and (_15677_, _15662_, _15537_);
  or (_40850_, _15677_, _15676_);
  or (_15678_, _15660_, _14852_);
  or (_15679_, _15659_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_15680_, _15679_, _15663_);
  and (_15681_, _15680_, _15678_);
  and (_15682_, _15662_, _15543_);
  or (_40851_, _15682_, _15681_);
  or (_15683_, _15660_, _15058_);
  or (_15684_, _15659_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_15685_, _15684_, _15663_);
  and (_15686_, _15685_, _15683_);
  and (_15687_, _15662_, _15549_);
  or (_40853_, _15687_, _15686_);
  or (_15688_, _15660_, _15256_);
  or (_15689_, _15659_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_15690_, _15689_, _15663_);
  and (_15691_, _15690_, _15688_);
  and (_15692_, _15662_, _15555_);
  or (_40854_, _15692_, _15691_);
  or (_15693_, _15660_, _15454_);
  or (_15694_, _15659_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_15695_, _15694_, _15663_);
  and (_15696_, _15695_, _15693_);
  and (_15697_, _15662_, _15561_);
  or (_40855_, _15697_, _15696_);
  or (_15698_, _15660_, _09197_);
  or (_15699_, _15659_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_15700_, _15699_, _15663_);
  and (_15701_, _15700_, _15698_);
  and (_15702_, _15662_, _09230_);
  or (_40856_, _15702_, _15701_);
  and (_15703_, _15613_, _08399_);
  not (_15704_, _15703_);
  and (_15705_, _15616_, _15520_);
  or (_15706_, _15705_, \oc8051_golden_model_1.IRAM[6] [0]);
  not (_15707_, _15705_);
  or (_15708_, _15707_, _14247_);
  and (_15709_, _15708_, _15706_);
  and (_15710_, _15709_, _15704_);
  and (_15711_, _15703_, _15516_);
  or (_40860_, _15711_, _15710_);
  or (_15712_, _15707_, _14436_);
  or (_15713_, _15705_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_15714_, _15713_, _15704_);
  and (_15715_, _15714_, _15712_);
  and (_15716_, _15703_, _15531_);
  or (_40861_, _15716_, _15715_);
  or (_15717_, _15707_, _14660_);
  or (_15718_, _15705_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_15719_, _15718_, _15704_);
  and (_15720_, _15719_, _15717_);
  and (_15721_, _15703_, _15537_);
  or (_40862_, _15721_, _15720_);
  or (_15722_, _15707_, _14852_);
  or (_15723_, _15705_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_15724_, _15723_, _15704_);
  and (_15725_, _15724_, _15722_);
  and (_15726_, _15703_, _15543_);
  or (_40863_, _15726_, _15725_);
  or (_15727_, _15707_, _15058_);
  or (_15728_, _15705_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_15729_, _15728_, _15704_);
  and (_15730_, _15729_, _15727_);
  and (_15731_, _15703_, _15549_);
  or (_40864_, _15731_, _15730_);
  or (_15732_, _15707_, _15256_);
  or (_15733_, _15705_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_15734_, _15733_, _15704_);
  and (_15735_, _15734_, _15732_);
  and (_15736_, _15703_, _15555_);
  or (_40865_, _15736_, _15735_);
  or (_15737_, _15707_, _15454_);
  or (_15738_, _15705_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_15739_, _15738_, _15704_);
  and (_15740_, _15739_, _15737_);
  and (_15741_, _15703_, _15561_);
  or (_40866_, _15741_, _15740_);
  and (_15742_, _15705_, _09197_);
  nor (_15743_, _15705_, _07751_);
  or (_15744_, _15743_, _15703_);
  or (_15745_, _15744_, _15742_);
  or (_15746_, _15704_, _09230_);
  and (_40867_, _15746_, _15745_);
  and (_15747_, _15613_, _07080_);
  not (_15748_, _15747_);
  or (_15749_, _15748_, _15516_);
  and (_15750_, _15616_, _07307_);
  and (_15751_, _15750_, _14247_);
  nor (_15752_, _15750_, _06895_);
  or (_15753_, _15752_, _15747_);
  or (_15754_, _15753_, _15751_);
  and (_40872_, _15754_, _15749_);
  or (_15755_, _15750_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_15756_, _15755_, _15748_);
  not (_15757_, _15750_);
  or (_15758_, _15757_, _14436_);
  and (_15759_, _15758_, _15756_);
  and (_15760_, _15747_, _15531_);
  or (_40873_, _15760_, _15759_);
  or (_15761_, _15750_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_15762_, _15761_, _15748_);
  or (_15763_, _15757_, _14660_);
  and (_15764_, _15763_, _15762_);
  and (_15765_, _15747_, _15537_);
  or (_40874_, _15765_, _15764_);
  or (_15766_, _15750_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_15767_, _15766_, _15748_);
  or (_15768_, _15757_, _14852_);
  and (_15769_, _15768_, _15767_);
  and (_15770_, _15747_, _15543_);
  or (_40876_, _15770_, _15769_);
  or (_15771_, _15750_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_15772_, _15771_, _15748_);
  or (_15773_, _15757_, _15058_);
  and (_15774_, _15773_, _15772_);
  and (_15775_, _15747_, _15549_);
  or (_40877_, _15775_, _15774_);
  or (_15776_, _15750_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_15777_, _15776_, _15748_);
  or (_15778_, _15757_, _15256_);
  and (_15779_, _15778_, _15777_);
  and (_15780_, _15747_, _15555_);
  or (_40878_, _15780_, _15779_);
  or (_15781_, _15750_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_15782_, _15781_, _15748_);
  or (_15783_, _15757_, _15454_);
  and (_15784_, _15783_, _15782_);
  and (_15785_, _15747_, _15561_);
  or (_40879_, _15785_, _15784_);
  or (_15786_, _15750_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_15787_, _15786_, _15748_);
  or (_15788_, _15757_, _09197_);
  and (_15789_, _15788_, _15787_);
  and (_15790_, _15747_, _09230_);
  or (_40880_, _15790_, _15789_);
  and (_15791_, _14075_, _07614_);
  and (_15792_, _15791_, _14078_);
  or (_15793_, _15792_, \oc8051_golden_model_1.IRAM[8] [0]);
  not (_15794_, _15792_);
  or (_15795_, _15794_, _14247_);
  and (_15796_, _15795_, _15793_);
  and (_15797_, _07629_, _14449_);
  and (_15798_, _15797_, _07081_);
  or (_15799_, _15798_, _15796_);
  not (_15800_, _15798_);
  or (_15801_, _15800_, _15516_);
  and (_40884_, _15801_, _15799_);
  or (_15802_, _15794_, _14436_);
  or (_15803_, _15792_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_15804_, _15803_, _15800_);
  and (_15805_, _15804_, _15802_);
  and (_15806_, _15798_, _15531_);
  or (_40885_, _15806_, _15805_);
  or (_15807_, _15794_, _14660_);
  or (_15808_, _15792_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_15809_, _15808_, _15800_);
  and (_15810_, _15809_, _15807_);
  and (_15811_, _15798_, _15537_);
  or (_40886_, _15811_, _15810_);
  or (_15812_, _15794_, _14852_);
  or (_15813_, _15792_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_15814_, _15813_, _15800_);
  and (_15815_, _15814_, _15812_);
  and (_15816_, _15798_, _15543_);
  or (_40887_, _15816_, _15815_);
  or (_15817_, _15794_, _15058_);
  or (_15818_, _15792_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_15819_, _15818_, _15800_);
  and (_15820_, _15819_, _15817_);
  and (_15821_, _15798_, _15549_);
  or (_40889_, _15821_, _15820_);
  or (_15822_, _15794_, _15256_);
  or (_15823_, _15792_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_15824_, _15823_, _15800_);
  and (_15825_, _15824_, _15822_);
  and (_15826_, _15798_, _15555_);
  or (_40890_, _15826_, _15825_);
  or (_15827_, _15794_, _15454_);
  or (_15828_, _15792_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_15829_, _15828_, _15800_);
  and (_15830_, _15829_, _15827_);
  and (_15831_, _15798_, _15561_);
  or (_40891_, _15831_, _15830_);
  or (_15832_, _15794_, _09197_);
  or (_15833_, _15792_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_15834_, _15833_, _15800_);
  and (_15835_, _15834_, _15832_);
  and (_15836_, _15798_, _09230_);
  or (_40892_, _15836_, _15835_);
  and (_15837_, _15791_, _15472_);
  or (_15838_, _15837_, \oc8051_golden_model_1.IRAM[9] [0]);
  not (_15839_, _15837_);
  or (_15840_, _15839_, _14247_);
  and (_15841_, _15840_, _15838_);
  and (_15842_, _15797_, _07356_);
  or (_15843_, _15842_, _15841_);
  not (_15844_, _15842_);
  or (_15845_, _15844_, _15516_);
  and (_40896_, _15845_, _15843_);
  or (_15846_, _15839_, _14436_);
  or (_15847_, _15837_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_15848_, _15847_, _15844_);
  and (_15849_, _15848_, _15846_);
  and (_15850_, _15842_, _15531_);
  or (_40897_, _15850_, _15849_);
  or (_15851_, _15839_, _14660_);
  or (_15852_, _15837_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_15853_, _15852_, _15844_);
  and (_15854_, _15853_, _15851_);
  and (_15855_, _15842_, _15537_);
  or (_40898_, _15855_, _15854_);
  or (_15856_, _15839_, _14852_);
  or (_15857_, _15837_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_15858_, _15857_, _15844_);
  and (_15859_, _15858_, _15856_);
  and (_15860_, _15842_, _15543_);
  or (_40899_, _15860_, _15859_);
  or (_15861_, _15839_, _15058_);
  or (_15862_, _15837_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_15863_, _15862_, _15844_);
  and (_15864_, _15863_, _15861_);
  and (_15865_, _15842_, _15549_);
  or (_40901_, _15865_, _15864_);
  or (_15866_, _15839_, _15256_);
  or (_15867_, _15837_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_15868_, _15867_, _15844_);
  and (_15869_, _15868_, _15866_);
  and (_15870_, _15842_, _15555_);
  or (_40902_, _15870_, _15869_);
  or (_15871_, _15839_, _15454_);
  or (_15872_, _15837_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_15873_, _15872_, _15844_);
  and (_15874_, _15873_, _15871_);
  and (_15875_, _15842_, _15561_);
  or (_40903_, _15875_, _15874_);
  nor (_15876_, _15839_, _09197_);
  nor (_15877_, _15837_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_15878_, _15877_, _15876_);
  nor (_15879_, _15878_, _15842_);
  and (_15880_, _15842_, _09230_);
  or (_40904_, _15880_, _15879_);
  and (_15881_, _15791_, _15520_);
  not (_15882_, _15881_);
  or (_15883_, _15882_, _14247_);
  and (_15884_, _15797_, _08399_);
  not (_15885_, _15884_);
  or (_15886_, _15881_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_15887_, _15886_, _15885_);
  and (_15888_, _15887_, _15883_);
  and (_15889_, _15884_, _15516_);
  or (_40908_, _15889_, _15888_);
  or (_15890_, _15882_, _14436_);
  or (_15891_, _15881_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_15892_, _15891_, _15885_);
  and (_15893_, _15892_, _15890_);
  and (_15894_, _15884_, _15531_);
  or (_40909_, _15894_, _15893_);
  or (_15895_, _15882_, _14660_);
  or (_15896_, _15881_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_15897_, _15896_, _15885_);
  and (_15898_, _15897_, _15895_);
  and (_15899_, _15884_, _15537_);
  or (_40910_, _15899_, _15898_);
  or (_15900_, _15882_, _14852_);
  or (_15901_, _15881_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_15902_, _15901_, _15885_);
  and (_15903_, _15902_, _15900_);
  and (_15904_, _15884_, _15543_);
  or (_40912_, _15904_, _15903_);
  or (_15905_, _15882_, _15058_);
  or (_15906_, _15881_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_15907_, _15906_, _15885_);
  and (_15908_, _15907_, _15905_);
  and (_15909_, _15884_, _15549_);
  or (_40913_, _15909_, _15908_);
  or (_15910_, _15882_, _15256_);
  or (_15911_, _15881_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_15912_, _15911_, _15885_);
  and (_15913_, _15912_, _15910_);
  and (_15914_, _15884_, _15555_);
  or (_40914_, _15914_, _15913_);
  or (_15915_, _15882_, _15454_);
  or (_15916_, _15881_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_15917_, _15916_, _15885_);
  and (_15918_, _15917_, _15915_);
  and (_15919_, _15884_, _15561_);
  or (_40915_, _15919_, _15918_);
  or (_15920_, _15882_, _09197_);
  or (_15921_, _15881_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_15922_, _15921_, _15885_);
  and (_15923_, _15922_, _15920_);
  and (_15924_, _15884_, _09230_);
  or (_40916_, _15924_, _15923_);
  not (_15925_, _07229_);
  and (_15926_, _14077_, _15925_);
  and (_15927_, _15791_, _15926_);
  nor (_15928_, _15927_, \oc8051_golden_model_1.IRAM[11] [0]);
  not (_15929_, _15927_);
  nor (_15930_, _15929_, _14247_);
  or (_15931_, _15930_, _15928_);
  and (_15932_, _15797_, _07080_);
  not (_15933_, _15932_);
  nand (_15934_, _15933_, _15931_);
  or (_15935_, _15933_, _15516_);
  and (_40919_, _15935_, _15934_);
  or (_15936_, _15927_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_15937_, _15936_, _15933_);
  or (_15938_, _15929_, _14436_);
  and (_15939_, _15938_, _15937_);
  and (_15940_, _15932_, _15531_);
  or (_40920_, _15940_, _15939_);
  or (_15941_, _15927_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_15942_, _15941_, _15933_);
  or (_15943_, _15929_, _14660_);
  and (_15944_, _15943_, _15942_);
  and (_15945_, _15932_, _15537_);
  or (_40921_, _15945_, _15944_);
  or (_15946_, _15927_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_15947_, _15946_, _15933_);
  or (_15948_, _15929_, _14852_);
  and (_15949_, _15948_, _15947_);
  and (_15950_, _15932_, _15543_);
  or (_40924_, _15950_, _15949_);
  or (_15951_, _15927_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_15952_, _15951_, _15933_);
  or (_15953_, _15929_, _15058_);
  and (_15954_, _15953_, _15952_);
  and (_15955_, _15932_, _15549_);
  or (_40925_, _15955_, _15954_);
  or (_15956_, _15927_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_15957_, _15956_, _15933_);
  or (_15958_, _15929_, _15256_);
  and (_15959_, _15958_, _15957_);
  and (_15960_, _15932_, _15555_);
  or (_40926_, _15960_, _15959_);
  or (_15961_, _15927_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_15962_, _15961_, _15933_);
  or (_15963_, _15929_, _15454_);
  and (_15964_, _15963_, _15962_);
  and (_15965_, _15932_, _15561_);
  or (_40927_, _15965_, _15964_);
  or (_15966_, _15927_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_15967_, _15966_, _15933_);
  or (_15968_, _15929_, _09197_);
  and (_15969_, _15968_, _15967_);
  and (_15970_, _15932_, _09230_);
  or (_40928_, _15970_, _15969_);
  not (_15971_, _07614_);
  and (_15972_, _14075_, _15971_);
  and (_15973_, _14078_, _15972_);
  not (_15974_, _15973_);
  or (_15975_, _15974_, _14247_);
  or (_15976_, _15973_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_15977_, _15976_, _15975_);
  and (_15978_, _07630_, _07081_);
  or (_15979_, _15978_, _15977_);
  not (_15980_, _15978_);
  or (_15981_, _15980_, _15516_);
  and (_40932_, _15981_, _15979_);
  and (_15982_, _14078_, _07617_);
  or (_15983_, _15982_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_15984_, _15983_, _15980_);
  not (_15985_, _15982_);
  or (_15986_, _15985_, _14436_);
  and (_15987_, _15986_, _15984_);
  and (_15988_, _15978_, _15531_);
  or (_40933_, _15988_, _15987_);
  or (_15989_, _15982_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_15990_, _15989_, _15980_);
  or (_15991_, _15985_, _14660_);
  and (_15992_, _15991_, _15990_);
  and (_15993_, _15978_, _15537_);
  or (_40934_, _15993_, _15992_);
  or (_15994_, _15982_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_15995_, _15994_, _15980_);
  or (_15996_, _15985_, _14852_);
  and (_15997_, _15996_, _15995_);
  and (_15998_, _15978_, _15543_);
  or (_40935_, _15998_, _15997_);
  or (_15999_, _15982_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_16000_, _15999_, _15980_);
  or (_16001_, _15985_, _15058_);
  and (_16002_, _16001_, _16000_);
  and (_16003_, _15978_, _15549_);
  or (_40936_, _16003_, _16002_);
  or (_16004_, _15982_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_16005_, _16004_, _15980_);
  or (_16006_, _15985_, _15256_);
  and (_16007_, _16006_, _16005_);
  and (_16008_, _15978_, _15555_);
  or (_40937_, _16008_, _16007_);
  or (_16009_, _15982_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_16010_, _16009_, _15980_);
  or (_16011_, _15985_, _15454_);
  and (_16012_, _16011_, _16010_);
  and (_16013_, _15978_, _15561_);
  or (_40939_, _16013_, _16012_);
  or (_16014_, _15982_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_16015_, _16014_, _15980_);
  or (_16016_, _15985_, _09197_);
  and (_16017_, _16016_, _16015_);
  and (_16018_, _15978_, _09230_);
  or (_40940_, _16018_, _16017_);
  and (_16019_, _15472_, _15972_);
  not (_16020_, _16019_);
  or (_16021_, _16020_, _14247_);
  and (_16022_, _07630_, _07356_);
  not (_16023_, _16022_);
  or (_16024_, _16019_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_16025_, _16024_, _16023_);
  and (_16026_, _16025_, _16021_);
  and (_16027_, _16022_, _15516_);
  or (_40943_, _16027_, _16026_);
  and (_16028_, _15472_, _07617_);
  or (_16029_, _16028_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_16030_, _16029_, _16023_);
  not (_16031_, _16028_);
  or (_16032_, _16031_, _14436_);
  and (_16033_, _16032_, _16030_);
  and (_16034_, _16022_, _15531_);
  or (_40945_, _16034_, _16033_);
  or (_16035_, _16028_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_16036_, _16035_, _16023_);
  or (_16037_, _16031_, _14660_);
  and (_16038_, _16037_, _16036_);
  and (_16039_, _16022_, _15537_);
  or (_40946_, _16039_, _16038_);
  or (_16040_, _16028_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_16041_, _16040_, _16023_);
  or (_16042_, _16031_, _14852_);
  and (_16043_, _16042_, _16041_);
  and (_16044_, _16022_, _15543_);
  or (_40947_, _16044_, _16043_);
  or (_16045_, _16028_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_16046_, _16045_, _16023_);
  or (_16047_, _16031_, _15058_);
  and (_16048_, _16047_, _16046_);
  and (_16049_, _16022_, _15549_);
  or (_40948_, _16049_, _16048_);
  or (_16050_, _16028_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_16051_, _16050_, _16023_);
  or (_16052_, _16031_, _15256_);
  and (_16053_, _16052_, _16051_);
  and (_16054_, _16022_, _15555_);
  or (_40949_, _16054_, _16053_);
  or (_16055_, _16028_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_16056_, _16055_, _16023_);
  or (_16057_, _16031_, _15454_);
  and (_16058_, _16057_, _16056_);
  and (_16059_, _16022_, _15561_);
  or (_40951_, _16059_, _16058_);
  nor (_16060_, _16019_, \oc8051_golden_model_1.IRAM[13] [7]);
  nor (_16061_, _16020_, _09197_);
  or (_16062_, _16061_, _16060_);
  nand (_16063_, _16062_, _16023_);
  or (_16064_, _16023_, _09230_);
  and (_40952_, _16064_, _16063_);
  and (_16065_, _15520_, _15972_);
  not (_16066_, _16065_);
  or (_16067_, _16066_, _14247_);
  and (_16068_, _08399_, _07630_);
  not (_16069_, _16068_);
  or (_16070_, _16065_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_16071_, _16070_, _16069_);
  and (_16072_, _16071_, _16067_);
  and (_16073_, _16068_, _15516_);
  or (_40956_, _16073_, _16072_);
  and (_16074_, _15520_, _07617_);
  or (_16075_, _16074_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_16076_, _16075_, _16069_);
  not (_16077_, _16074_);
  or (_16078_, _16077_, _14436_);
  and (_16079_, _16078_, _16076_);
  and (_16080_, _16068_, _15531_);
  or (_40957_, _16080_, _16079_);
  or (_16081_, _16074_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_16082_, _16081_, _16069_);
  or (_16083_, _16077_, _14660_);
  and (_16084_, _16083_, _16082_);
  and (_16085_, _16068_, _15537_);
  or (_40958_, _16085_, _16084_);
  or (_16086_, _16074_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_16087_, _16086_, _16069_);
  or (_16088_, _16077_, _14852_);
  and (_16089_, _16088_, _16087_);
  and (_16090_, _16068_, _15543_);
  or (_40959_, _16090_, _16089_);
  or (_16091_, _16074_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_16092_, _16091_, _16069_);
  or (_16093_, _16077_, _15058_);
  and (_16094_, _16093_, _16092_);
  and (_16095_, _16068_, _15549_);
  or (_40960_, _16095_, _16094_);
  or (_16096_, _16074_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_16097_, _16096_, _16069_);
  or (_16098_, _16077_, _15256_);
  and (_16099_, _16098_, _16097_);
  and (_16100_, _16068_, _15555_);
  or (_40962_, _16100_, _16099_);
  or (_16101_, _16074_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_16102_, _16101_, _16069_);
  or (_16103_, _16077_, _15454_);
  and (_16104_, _16103_, _16102_);
  and (_16105_, _16068_, _15561_);
  or (_40963_, _16105_, _16104_);
  or (_16106_, _16074_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_16107_, _16106_, _16069_);
  or (_16108_, _16077_, _09197_);
  and (_16109_, _16108_, _16107_);
  and (_16110_, _16068_, _09230_);
  or (_40964_, _16110_, _16109_);
  nand (_16111_, _15972_, _15926_);
  or (_16112_, _14247_, _16111_);
  or (_16113_, _07618_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_16114_, _16113_, _07632_);
  and (_16115_, _16114_, _16112_);
  and (_16116_, _15516_, _07631_);
  or (_40967_, _16116_, _16115_);
  or (_16117_, _07618_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_16118_, _16117_, _07632_);
  or (_16119_, _14436_, _07634_);
  and (_16120_, _16119_, _16118_);
  and (_16121_, _15531_, _07631_);
  or (_40968_, _16121_, _16120_);
  or (_16122_, _07618_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_16123_, _16122_, _07632_);
  or (_16124_, _14660_, _07634_);
  and (_16125_, _16124_, _16123_);
  and (_16126_, _15537_, _07631_);
  or (_40969_, _16126_, _16125_);
  or (_16127_, _07618_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_16128_, _16127_, _07632_);
  or (_16129_, _14852_, _07634_);
  and (_16130_, _16129_, _16128_);
  and (_16131_, _15543_, _07631_);
  or (_40970_, _16131_, _16130_);
  or (_16132_, _07618_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_16133_, _16132_, _07632_);
  or (_16134_, _15058_, _07634_);
  and (_16135_, _16134_, _16133_);
  and (_16136_, _15549_, _07631_);
  or (_40971_, _16136_, _16135_);
  or (_16137_, _15256_, _07634_);
  or (_16138_, _07618_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_16139_, _16138_, _07632_);
  and (_16140_, _16139_, _16137_);
  and (_16141_, _15555_, _07631_);
  or (_40972_, _16141_, _16140_);
  or (_16142_, _15454_, _07634_);
  or (_16143_, _07618_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_16144_, _16143_, _07632_);
  and (_16145_, _16144_, _16142_);
  and (_16146_, _15561_, _07631_);
  or (_40973_, _16146_, _16145_);
  nor (_16147_, _01336_, _09877_);
  nor (_16148_, _07698_, _09877_);
  and (_16149_, _07698_, _08672_);
  or (_16150_, _16149_, _16148_);
  or (_16151_, _16150_, _06020_);
  and (_16152_, _14186_, _07698_);
  or (_16153_, _16152_, _16148_);
  and (_16154_, _16153_, _09833_);
  nor (_16155_, _08127_, _09258_);
  or (_16156_, _16155_, _16148_);
  and (_16157_, _16156_, _06102_);
  nor (_16158_, _06938_, _09877_);
  and (_16159_, _07698_, \oc8051_golden_model_1.ACC [0]);
  or (_16160_, _16159_, _16148_);
  and (_16161_, _16160_, _06938_);
  or (_16162_, _16161_, _16158_);
  and (_16163_, _16162_, _06954_);
  or (_16164_, _16163_, _06043_);
  or (_16165_, _16164_, _16157_);
  and (_16166_, _14102_, _08361_);
  nor (_16167_, _08361_, _09877_);
  or (_16168_, _16167_, _06044_);
  or (_16169_, _16168_, _16166_);
  and (_16170_, _16169_, _16165_);
  or (_16171_, _16170_, _06239_);
  and (_16172_, _07698_, _06931_);
  or (_16173_, _16172_, _16148_);
  or (_16174_, _16173_, _06848_);
  and (_16175_, _16174_, _16171_);
  or (_16176_, _16175_, _06219_);
  or (_16177_, _16160_, _06220_);
  and (_16178_, _16177_, _06040_);
  and (_16179_, _16178_, _16176_);
  and (_16180_, _16148_, _06039_);
  or (_16181_, _16180_, _06032_);
  or (_16182_, _16181_, _16179_);
  or (_16183_, _16156_, _06033_);
  and (_16184_, _16183_, _16182_);
  or (_16185_, _16184_, _09269_);
  nor (_16186_, _09765_, _09763_);
  nor (_16187_, _16186_, _09766_);
  or (_16188_, _16187_, _09800_);
  and (_16189_, _16188_, _06027_);
  and (_16190_, _16189_, _16185_);
  and (_16191_, _14132_, _08361_);
  or (_16192_, _16191_, _16167_);
  and (_16193_, _16192_, _06026_);
  or (_16194_, _16193_, _09818_);
  or (_16195_, _16194_, _16190_);
  and (_16196_, _09120_, _07698_);
  or (_16197_, _16148_, _07012_);
  or (_16198_, _16197_, _16196_);
  or (_16199_, _16173_, _09827_);
  and (_16200_, _16199_, _05669_);
  and (_16201_, _16200_, _16198_);
  and (_16202_, _16201_, _16195_);
  or (_16203_, _16202_, _16154_);
  and (_16204_, _16203_, _09839_);
  nand (_16205_, _10184_, _05758_);
  or (_16206_, _10178_, _10133_);
  or (_16207_, _10184_, _16206_);
  and (_16208_, _16207_, _09832_);
  and (_16209_, _16208_, _16205_);
  or (_16210_, _16209_, _06019_);
  or (_16211_, _16210_, _16204_);
  and (_16212_, _16211_, _16151_);
  or (_16213_, _16212_, _06112_);
  and (_16214_, _14086_, _07698_);
  or (_16215_, _16148_, _08751_);
  or (_16216_, _16215_, _16214_);
  and (_16217_, _16216_, _08756_);
  and (_16218_, _16217_, _16213_);
  nor (_16219_, _12302_, _09258_);
  or (_16220_, _16219_, _16148_);
  nand (_16221_, _10995_, _07698_);
  and (_16222_, _16221_, _06284_);
  and (_16223_, _16222_, _16220_);
  or (_16224_, _16223_, _16218_);
  and (_16225_, _16224_, _07032_);
  nand (_16226_, _16150_, _06108_);
  nor (_16227_, _16226_, _16155_);
  or (_16228_, _16227_, _06277_);
  or (_16229_, _16228_, _16225_);
  nor (_16230_, _16148_, _06278_);
  nand (_16231_, _16230_, _16221_);
  and (_16232_, _16231_, _16229_);
  or (_16233_, _16232_, _06130_);
  and (_16234_, _14083_, _07698_);
  or (_16235_, _16148_, _08777_);
  or (_16236_, _16235_, _16234_);
  and (_16237_, _16236_, _08782_);
  and (_16238_, _16237_, _16233_);
  and (_16239_, _16220_, _06292_);
  or (_16240_, _16239_, _06316_);
  or (_16241_, _16240_, _16238_);
  or (_16242_, _16156_, _06718_);
  and (_16243_, _16242_, _16241_);
  or (_16244_, _16243_, _05652_);
  or (_16245_, _16148_, _05653_);
  and (_16246_, _16245_, _16244_);
  or (_16247_, _16246_, _06047_);
  or (_16248_, _16156_, _06048_);
  and (_16249_, _16248_, _01336_);
  and (_16250_, _16249_, _16247_);
  or (_16251_, _16250_, _16147_);
  and (_43324_, _16251_, _42882_);
  nor (_16252_, _01336_, _09842_);
  nor (_16253_, _07698_, _09842_);
  nor (_16254_, _10993_, _09258_);
  or (_16255_, _16254_, _16253_);
  or (_16256_, _16255_, _08782_);
  nor (_16257_, _08361_, _09842_);
  and (_16258_, _14273_, _08361_);
  or (_16259_, _16258_, _16257_);
  and (_16260_, _16259_, _06039_);
  nor (_16261_, _09258_, _07132_);
  or (_16262_, _16261_, _16253_);
  or (_16263_, _16262_, _06848_);
  or (_16264_, _07698_, \oc8051_golden_model_1.B [1]);
  and (_16265_, _14284_, _07698_);
  not (_16266_, _16265_);
  and (_16267_, _16266_, _16264_);
  or (_16268_, _16267_, _06954_);
  and (_16269_, _07698_, \oc8051_golden_model_1.ACC [1]);
  or (_16270_, _16269_, _16253_);
  and (_16271_, _16270_, _06938_);
  nor (_16272_, _06938_, _09842_);
  or (_16273_, _16272_, _06102_);
  or (_16274_, _16273_, _16271_);
  and (_16275_, _16274_, _06044_);
  and (_16276_, _16275_, _16268_);
  and (_16277_, _14266_, _08361_);
  or (_16278_, _16277_, _16257_);
  and (_16279_, _16278_, _06043_);
  or (_16280_, _16279_, _06239_);
  or (_16281_, _16280_, _16276_);
  and (_16282_, _16281_, _16263_);
  or (_16283_, _16282_, _06219_);
  or (_16284_, _16270_, _06220_);
  and (_16285_, _16284_, _06040_);
  and (_16286_, _16285_, _16283_);
  or (_16287_, _16286_, _16260_);
  and (_16288_, _16287_, _06033_);
  and (_16289_, _16277_, _14302_);
  or (_16290_, _16289_, _16257_);
  and (_16291_, _16290_, _06032_);
  or (_16292_, _16291_, _09269_);
  or (_16293_, _16292_, _16288_);
  nor (_16294_, _09768_, _09699_);
  nor (_16295_, _16294_, _09769_);
  or (_16296_, _16295_, _09800_);
  and (_16297_, _16296_, _06027_);
  and (_16298_, _16297_, _16293_);
  or (_16299_, _16257_, _14267_);
  and (_16300_, _16299_, _06026_);
  and (_16301_, _16300_, _16278_);
  or (_16302_, _16301_, _09818_);
  or (_16303_, _16302_, _16298_);
  and (_16304_, _09075_, _07698_);
  or (_16305_, _16253_, _07012_);
  or (_16306_, _16305_, _16304_);
  or (_16307_, _16262_, _09827_);
  and (_16308_, _16307_, _05669_);
  and (_16309_, _16308_, _16306_);
  and (_16310_, _16309_, _16303_);
  or (_16311_, _14367_, _09258_);
  and (_16312_, _16264_, _09833_);
  and (_16313_, _16312_, _16311_);
  or (_16314_, _16313_, _09832_);
  or (_16315_, _16314_, _16310_);
  nor (_16316_, _10179_, _10177_);
  or (_16317_, _16316_, _10180_);
  nor (_16318_, _16317_, _10184_);
  and (_16319_, _10184_, _10130_);
  or (_16320_, _16319_, _16318_);
  or (_16321_, _16320_, _09839_);
  and (_16322_, _16321_, _06020_);
  and (_16323_, _16322_, _16315_);
  nand (_16324_, _07698_, _06832_);
  and (_16325_, _16264_, _06019_);
  and (_16326_, _16325_, _16324_);
  or (_16327_, _16326_, _16323_);
  and (_16328_, _16327_, _08751_);
  or (_16329_, _14263_, _09258_);
  and (_16330_, _16264_, _06112_);
  and (_16331_, _16330_, _16329_);
  or (_16332_, _16331_, _06284_);
  or (_16333_, _16332_, _16328_);
  and (_16334_, _10994_, _07698_);
  or (_16335_, _16334_, _16253_);
  or (_16336_, _16335_, _08756_);
  and (_16337_, _16336_, _07032_);
  and (_16338_, _16337_, _16333_);
  or (_16339_, _14261_, _09258_);
  and (_16340_, _16264_, _06108_);
  and (_16341_, _16340_, _16339_);
  or (_16342_, _16341_, _06277_);
  or (_16343_, _16342_, _16338_);
  and (_16344_, _16269_, _08078_);
  or (_16345_, _16253_, _06278_);
  or (_16346_, _16345_, _16344_);
  and (_16347_, _16346_, _08777_);
  and (_16348_, _16347_, _16343_);
  or (_16349_, _16324_, _08078_);
  and (_16350_, _16264_, _06130_);
  and (_16351_, _16350_, _16349_);
  or (_16352_, _16351_, _06292_);
  or (_16353_, _16352_, _16348_);
  and (_16354_, _16353_, _16256_);
  or (_16355_, _16354_, _06316_);
  or (_16356_, _16267_, _06718_);
  and (_16357_, _16356_, _05653_);
  and (_16358_, _16357_, _16355_);
  and (_16359_, _16259_, _05652_);
  or (_16360_, _16359_, _06047_);
  or (_16361_, _16360_, _16358_);
  or (_16362_, _16253_, _06048_);
  or (_16363_, _16362_, _16265_);
  and (_16364_, _16363_, _01336_);
  and (_16365_, _16364_, _16361_);
  or (_16366_, _16365_, _16252_);
  and (_43325_, _16366_, _42882_);
  nor (_16367_, _01336_, _10002_);
  nor (_16368_, _07698_, _10002_);
  and (_16369_, _07698_, _08730_);
  or (_16370_, _16369_, _16368_);
  or (_16371_, _16370_, _06020_);
  and (_16372_, _14580_, _07698_);
  or (_16373_, _16372_, _16368_);
  and (_16374_, _16373_, _09833_);
  nor (_16375_, _08361_, _10002_);
  and (_16376_, _14479_, _08361_);
  or (_16377_, _16376_, _16375_);
  and (_16378_, _16377_, _06039_);
  and (_16379_, _14493_, _07698_);
  or (_16380_, _16379_, _16368_);
  and (_16381_, _16380_, _06102_);
  nor (_16382_, _06938_, _10002_);
  and (_16383_, _07698_, \oc8051_golden_model_1.ACC [2]);
  or (_16384_, _16383_, _16368_);
  and (_16385_, _16384_, _06938_);
  or (_16386_, _16385_, _16382_);
  and (_16387_, _16386_, _06954_);
  or (_16388_, _16387_, _06043_);
  or (_16389_, _16388_, _16381_);
  and (_16390_, _14497_, _08361_);
  or (_16391_, _16390_, _16375_);
  or (_16392_, _16391_, _06044_);
  and (_16393_, _16392_, _06848_);
  and (_16394_, _16393_, _16389_);
  nor (_16395_, _09258_, _07530_);
  or (_16396_, _16395_, _16368_);
  and (_16397_, _16396_, _06239_);
  or (_16398_, _16397_, _06219_);
  or (_16399_, _16398_, _16394_);
  or (_16400_, _16384_, _06220_);
  and (_16401_, _16400_, _06040_);
  and (_16402_, _16401_, _16399_);
  or (_16403_, _16402_, _16378_);
  and (_16404_, _16403_, _06033_);
  or (_16405_, _16375_, _14512_);
  and (_16406_, _16391_, _06032_);
  and (_16407_, _16406_, _16405_);
  or (_16408_, _16407_, _09269_);
  or (_16409_, _16408_, _16404_);
  or (_16410_, _09770_, _09652_);
  and (_16411_, _16410_, _09771_);
  or (_16412_, _16411_, _09800_);
  and (_16413_, _16412_, _06027_);
  and (_16414_, _16413_, _16409_);
  or (_16415_, _16375_, _14525_);
  and (_16416_, _16415_, _06026_);
  and (_16417_, _16416_, _16391_);
  or (_16418_, _16417_, _09818_);
  or (_16419_, _16418_, _16414_);
  and (_16420_, _09182_, _07698_);
  or (_16421_, _16368_, _07012_);
  or (_16422_, _16421_, _16420_);
  or (_16423_, _16396_, _09827_);
  and (_16424_, _16423_, _05669_);
  and (_16425_, _16424_, _16422_);
  and (_16426_, _16425_, _16419_);
  or (_16427_, _16426_, _16374_);
  and (_16428_, _16427_, _09839_);
  nor (_16429_, _10180_, _10131_);
  not (_16430_, _16429_);
  and (_16431_, _16430_, _10124_);
  nor (_16432_, _16430_, _10124_);
  nor (_16433_, _16432_, _16431_);
  or (_16434_, _16433_, _10184_);
  nand (_16435_, _10184_, _10121_);
  and (_16436_, _16435_, _09832_);
  and (_16437_, _16436_, _16434_);
  or (_16438_, _16437_, _06019_);
  or (_16439_, _16438_, _16428_);
  and (_16440_, _16439_, _16371_);
  or (_16441_, _16440_, _06112_);
  and (_16442_, _14596_, _07698_);
  or (_16443_, _16442_, _16368_);
  or (_16444_, _16443_, _08751_);
  and (_16445_, _16444_, _08756_);
  and (_16446_, _16445_, _16441_);
  and (_16447_, _10991_, _07698_);
  or (_16448_, _16447_, _16368_);
  and (_16449_, _16448_, _06284_);
  or (_16450_, _16449_, _16446_);
  and (_16451_, _16450_, _07032_);
  or (_16452_, _16368_, _08177_);
  and (_16453_, _16370_, _06108_);
  and (_16454_, _16453_, _16452_);
  or (_16455_, _16454_, _16451_);
  and (_16456_, _16455_, _06278_);
  and (_16457_, _16384_, _06277_);
  and (_16458_, _16457_, _16452_);
  or (_16459_, _16458_, _06130_);
  or (_16460_, _16459_, _16456_);
  and (_16461_, _14593_, _07698_);
  or (_16462_, _16368_, _08777_);
  or (_16463_, _16462_, _16461_);
  and (_16464_, _16463_, _08782_);
  and (_16465_, _16464_, _16460_);
  nor (_16466_, _10990_, _09258_);
  or (_16467_, _16466_, _16368_);
  and (_16468_, _16467_, _06292_);
  or (_16469_, _16468_, _06316_);
  or (_16470_, _16469_, _16465_);
  or (_16471_, _16380_, _06718_);
  and (_16472_, _16471_, _05653_);
  and (_16473_, _16472_, _16470_);
  and (_16474_, _16377_, _05652_);
  or (_16475_, _16474_, _06047_);
  or (_16476_, _16475_, _16473_);
  and (_16477_, _14657_, _07698_);
  or (_16478_, _16368_, _06048_);
  or (_16479_, _16478_, _16477_);
  and (_16480_, _16479_, _01336_);
  and (_16481_, _16480_, _16476_);
  or (_16482_, _16481_, _16367_);
  and (_43326_, _16482_, _42882_);
  nor (_16483_, _01336_, _09927_);
  nor (_16484_, _07698_, _09927_);
  and (_16485_, _07698_, _08662_);
  or (_16486_, _16485_, _16484_);
  or (_16487_, _16486_, _06020_);
  and (_16488_, _14778_, _07698_);
  or (_16489_, _16488_, _16484_);
  and (_16490_, _16489_, _09833_);
  nor (_16491_, _08361_, _09927_);
  and (_16492_, _14683_, _08361_);
  or (_16493_, _16492_, _16491_);
  or (_16494_, _16491_, _14708_);
  and (_16495_, _16494_, _16493_);
  or (_16496_, _16495_, _06033_);
  and (_16497_, _14672_, _07698_);
  or (_16498_, _16497_, _16484_);
  or (_16499_, _16498_, _06954_);
  and (_16500_, _07698_, \oc8051_golden_model_1.ACC [3]);
  or (_16501_, _16500_, _16484_);
  and (_16502_, _16501_, _06938_);
  nor (_16503_, _06938_, _09927_);
  or (_16504_, _16503_, _06102_);
  or (_16505_, _16504_, _16502_);
  and (_16506_, _16505_, _06044_);
  and (_16507_, _16506_, _16499_);
  and (_16508_, _16493_, _06043_);
  or (_16509_, _16508_, _06239_);
  or (_16510_, _16509_, _16507_);
  nor (_16511_, _09258_, _07353_);
  or (_16512_, _16511_, _16484_);
  or (_16513_, _16512_, _06848_);
  and (_16514_, _16513_, _16510_);
  or (_16515_, _16514_, _06219_);
  or (_16516_, _16501_, _06220_);
  and (_16517_, _16516_, _06040_);
  and (_16518_, _16517_, _16515_);
  and (_16519_, _14681_, _08361_);
  or (_16520_, _16519_, _16491_);
  and (_16521_, _16520_, _06039_);
  or (_16522_, _16521_, _06032_);
  or (_16523_, _16522_, _16518_);
  and (_16524_, _16523_, _16496_);
  or (_16525_, _16524_, _09269_);
  nor (_16526_, _09773_, _09594_);
  nor (_16527_, _16526_, _09774_);
  or (_16528_, _16527_, _09800_);
  and (_16529_, _16528_, _06027_);
  and (_16530_, _16529_, _16525_);
  and (_16531_, _14724_, _08361_);
  or (_16532_, _16531_, _16491_);
  and (_16533_, _16532_, _06026_);
  or (_16534_, _16533_, _09818_);
  or (_16535_, _16534_, _16530_);
  and (_16536_, _09181_, _07698_);
  or (_16537_, _16484_, _07012_);
  or (_16538_, _16537_, _16536_);
  or (_16539_, _16512_, _09827_);
  and (_16540_, _16539_, _05669_);
  and (_16541_, _16540_, _16538_);
  and (_16542_, _16541_, _16535_);
  or (_16543_, _16542_, _16490_);
  and (_16544_, _16543_, _09839_);
  nor (_16545_, _16431_, _10123_);
  nor (_16546_, _16545_, _10115_);
  and (_16547_, _16545_, _10115_);
  or (_16548_, _16547_, _16546_);
  or (_16549_, _16548_, _10184_);
  not (_16550_, _10112_);
  nand (_16551_, _10184_, _16550_);
  and (_16552_, _16551_, _09832_);
  and (_16553_, _16552_, _16549_);
  or (_16554_, _16553_, _06019_);
  or (_16555_, _16554_, _16544_);
  and (_16556_, _16555_, _16487_);
  or (_16557_, _16556_, _06112_);
  and (_16558_, _14793_, _07698_);
  or (_16559_, _16484_, _08751_);
  or (_16560_, _16559_, _16558_);
  and (_16561_, _16560_, _08756_);
  and (_16562_, _16561_, _16557_);
  and (_16563_, _12299_, _07698_);
  or (_16564_, _16563_, _16484_);
  and (_16565_, _16564_, _06284_);
  or (_16566_, _16565_, _16562_);
  and (_16567_, _16566_, _07032_);
  or (_16568_, _16484_, _08029_);
  and (_16569_, _16486_, _06108_);
  and (_16570_, _16569_, _16568_);
  or (_16571_, _16570_, _16567_);
  and (_16572_, _16571_, _06278_);
  and (_16573_, _16501_, _06277_);
  and (_16574_, _16573_, _16568_);
  or (_16575_, _16574_, _06130_);
  or (_16576_, _16575_, _16572_);
  and (_16577_, _14792_, _07698_);
  or (_16578_, _16484_, _08777_);
  or (_16579_, _16578_, _16577_);
  and (_16580_, _16579_, _08782_);
  and (_16581_, _16580_, _16576_);
  nor (_16582_, _10988_, _09258_);
  or (_16583_, _16582_, _16484_);
  and (_16584_, _16583_, _06292_);
  or (_16585_, _16584_, _06316_);
  or (_16586_, _16585_, _16581_);
  or (_16587_, _16498_, _06718_);
  and (_16588_, _16587_, _05653_);
  and (_16589_, _16588_, _16586_);
  and (_16590_, _16520_, _05652_);
  or (_16591_, _16590_, _06047_);
  or (_16592_, _16591_, _16589_);
  and (_16593_, _14849_, _07698_);
  or (_16594_, _16484_, _06048_);
  or (_16595_, _16594_, _16593_);
  and (_16596_, _16595_, _01336_);
  and (_16597_, _16596_, _16592_);
  or (_16598_, _16597_, _16483_);
  and (_43327_, _16598_, _42882_);
  nor (_16599_, _01336_, _09854_);
  nor (_16600_, _07698_, _09854_);
  and (_16601_, _08665_, _07698_);
  or (_16602_, _16601_, _16600_);
  or (_16603_, _16602_, _06020_);
  and (_16604_, _14983_, _07698_);
  or (_16605_, _16604_, _16600_);
  and (_16606_, _16605_, _09833_);
  nor (_16607_, _08361_, _09854_);
  and (_16608_, _14882_, _08361_);
  or (_16609_, _16608_, _16607_);
  and (_16610_, _16609_, _06039_);
  and (_16611_, _14887_, _07698_);
  or (_16612_, _16611_, _16600_);
  or (_16613_, _16612_, _06954_);
  and (_16614_, _07698_, \oc8051_golden_model_1.ACC [4]);
  or (_16615_, _16614_, _16600_);
  and (_16616_, _16615_, _06938_);
  nor (_16617_, _06938_, _09854_);
  or (_16618_, _16617_, _06102_);
  or (_16619_, _16618_, _16616_);
  and (_16620_, _16619_, _06044_);
  and (_16621_, _16620_, _16613_);
  and (_16622_, _14878_, _08361_);
  or (_16623_, _16622_, _16607_);
  and (_16624_, _16623_, _06043_);
  or (_16625_, _16624_, _06239_);
  or (_16626_, _16625_, _16621_);
  nor (_16627_, _08270_, _09258_);
  or (_16628_, _16627_, _16600_);
  or (_16629_, _16628_, _06848_);
  and (_16630_, _16629_, _16626_);
  or (_16631_, _16630_, _06219_);
  or (_16632_, _16615_, _06220_);
  and (_16633_, _16632_, _06040_);
  and (_16634_, _16633_, _16631_);
  or (_16635_, _16634_, _16610_);
  and (_16636_, _16635_, _06033_);
  or (_16637_, _16607_, _14914_);
  and (_16638_, _16623_, _06032_);
  and (_16639_, _16638_, _16637_);
  or (_16640_, _16639_, _09269_);
  or (_16641_, _16640_, _16636_);
  or (_16642_, _09777_, _09775_);
  and (_16643_, _16642_, _09778_);
  or (_16644_, _16643_, _09800_);
  and (_16645_, _16644_, _06027_);
  and (_16646_, _16645_, _16641_);
  or (_16647_, _16607_, _14879_);
  and (_16648_, _16647_, _06026_);
  and (_16649_, _16648_, _16623_);
  or (_16650_, _16649_, _09818_);
  or (_16651_, _16650_, _16646_);
  and (_16652_, _09180_, _07698_);
  or (_16653_, _16600_, _07012_);
  or (_16654_, _16653_, _16652_);
  or (_16655_, _16628_, _09827_);
  and (_16656_, _16655_, _05669_);
  and (_16657_, _16656_, _16654_);
  and (_16658_, _16657_, _16651_);
  or (_16659_, _16658_, _16606_);
  and (_16660_, _16659_, _09839_);
  nand (_16661_, _10184_, _10147_);
  nor (_16662_, _16545_, _10114_);
  or (_16663_, _16662_, _10113_);
  nand (_16664_, _16663_, _10150_);
  or (_16665_, _16663_, _10150_);
  and (_16666_, _16665_, _16664_);
  or (_16667_, _16666_, _10184_);
  and (_16668_, _16667_, _09832_);
  and (_16669_, _16668_, _16661_);
  or (_16670_, _16669_, _06019_);
  or (_16671_, _16670_, _16660_);
  and (_16672_, _16671_, _16603_);
  or (_16673_, _16672_, _06112_);
  and (_16674_, _14876_, _07698_);
  or (_16675_, _16600_, _08751_);
  or (_16676_, _16675_, _16674_);
  and (_16677_, _16676_, _08756_);
  and (_16678_, _16677_, _16673_);
  and (_16679_, _10986_, _07698_);
  or (_16680_, _16679_, _16600_);
  and (_16681_, _16680_, _06284_);
  or (_16682_, _16681_, _16678_);
  and (_16683_, _16682_, _07032_);
  or (_16684_, _16600_, _08273_);
  and (_16685_, _16602_, _06108_);
  and (_16686_, _16685_, _16684_);
  or (_16687_, _16686_, _16683_);
  and (_16688_, _16687_, _06278_);
  and (_16689_, _16615_, _06277_);
  and (_16690_, _16689_, _16684_);
  or (_16691_, _16690_, _06130_);
  or (_16692_, _16691_, _16688_);
  and (_16693_, _14873_, _07698_);
  or (_16694_, _16600_, _08777_);
  or (_16695_, _16694_, _16693_);
  and (_16696_, _16695_, _08782_);
  and (_16697_, _16696_, _16692_);
  nor (_16698_, _10985_, _09258_);
  or (_16699_, _16698_, _16600_);
  and (_16700_, _16699_, _06292_);
  or (_16701_, _16700_, _06316_);
  or (_16702_, _16701_, _16697_);
  or (_16703_, _16612_, _06718_);
  and (_16704_, _16703_, _05653_);
  and (_16705_, _16704_, _16702_);
  and (_16706_, _16609_, _05652_);
  or (_16707_, _16706_, _06047_);
  or (_16708_, _16707_, _16705_);
  and (_16709_, _15055_, _07698_);
  or (_16710_, _16600_, _06048_);
  or (_16711_, _16710_, _16709_);
  and (_16712_, _16711_, _01336_);
  and (_16713_, _16712_, _16708_);
  or (_16714_, _16713_, _16599_);
  and (_43328_, _16714_, _42882_);
  nor (_16715_, _01336_, _09855_);
  nor (_16716_, _07698_, _09855_);
  and (_16717_, _15179_, _07698_);
  or (_16718_, _16717_, _16716_);
  and (_16719_, _16718_, _09833_);
  nor (_16720_, _08361_, _09855_);
  and (_16721_, _15077_, _08361_);
  or (_16722_, _16721_, _16720_);
  and (_16723_, _16722_, _06039_);
  and (_16724_, _15093_, _07698_);
  or (_16725_, _16724_, _16716_);
  or (_16726_, _16725_, _06954_);
  and (_16727_, _07698_, \oc8051_golden_model_1.ACC [5]);
  or (_16728_, _16727_, _16716_);
  and (_16729_, _16728_, _06938_);
  nor (_16730_, _06938_, _09855_);
  or (_16731_, _16730_, _06102_);
  or (_16732_, _16731_, _16729_);
  and (_16733_, _16732_, _06044_);
  and (_16734_, _16733_, _16726_);
  and (_16735_, _15073_, _08361_);
  or (_16736_, _16735_, _16720_);
  and (_16737_, _16736_, _06043_);
  or (_16738_, _16737_, _06239_);
  or (_16739_, _16738_, _16734_);
  nor (_16740_, _07977_, _09258_);
  or (_16741_, _16740_, _16716_);
  or (_16742_, _16741_, _06848_);
  and (_16743_, _16742_, _16739_);
  or (_16744_, _16743_, _06219_);
  or (_16745_, _16728_, _06220_);
  and (_16746_, _16745_, _06040_);
  and (_16747_, _16746_, _16744_);
  or (_16748_, _16747_, _16723_);
  and (_16749_, _16748_, _06033_);
  or (_16750_, _16720_, _15110_);
  and (_16751_, _16736_, _06032_);
  and (_16752_, _16751_, _16750_);
  or (_16753_, _16752_, _09269_);
  or (_16754_, _16753_, _16749_);
  or (_16755_, _09465_, _09466_);
  and (_16756_, _16755_, _09779_);
  nor (_16757_, _16756_, _09780_);
  or (_16758_, _16757_, _09800_);
  and (_16759_, _16758_, _06027_);
  and (_16760_, _16759_, _16754_);
  or (_16761_, _16720_, _15074_);
  and (_16762_, _16761_, _06026_);
  and (_16763_, _16762_, _16736_);
  or (_16764_, _16763_, _09818_);
  or (_16765_, _16764_, _16760_);
  and (_16766_, _09179_, _07698_);
  or (_16767_, _16716_, _07012_);
  or (_16768_, _16767_, _16766_);
  or (_16769_, _16741_, _09827_);
  and (_16770_, _16769_, _05669_);
  and (_16771_, _16770_, _16768_);
  and (_16772_, _16771_, _16765_);
  or (_16773_, _16772_, _16719_);
  and (_16774_, _16773_, _09839_);
  and (_16775_, _10184_, _09832_);
  and (_16776_, _16775_, _10157_);
  not (_16777_, _10149_);
  and (_16778_, _16664_, _16777_);
  nor (_16779_, _16778_, _10160_);
  and (_16780_, _16778_, _10160_);
  or (_16781_, _16780_, _16779_);
  nor (_16782_, _10184_, _09839_);
  and (_16783_, _16782_, _16781_);
  or (_16784_, _16783_, _16776_);
  or (_16785_, _16784_, _16774_);
  and (_16786_, _16785_, _06020_);
  and (_16787_, _08652_, _07698_);
  or (_16788_, _16787_, _16716_);
  and (_16789_, _16788_, _06019_);
  or (_16790_, _16789_, _06112_);
  or (_16791_, _16790_, _16786_);
  and (_16792_, _15195_, _07698_);
  or (_16793_, _16716_, _08751_);
  or (_16794_, _16793_, _16792_);
  and (_16795_, _16794_, _08756_);
  and (_16796_, _16795_, _16791_);
  and (_16797_, _12306_, _07698_);
  or (_16798_, _16797_, _16716_);
  and (_16799_, _16798_, _06284_);
  or (_16800_, _16799_, _16796_);
  and (_16801_, _16800_, _07032_);
  or (_16802_, _16716_, _07980_);
  and (_16803_, _16788_, _06108_);
  and (_16804_, _16803_, _16802_);
  or (_16805_, _16804_, _16801_);
  and (_16806_, _16805_, _06278_);
  and (_16807_, _16728_, _06277_);
  and (_16808_, _16807_, _16802_);
  or (_16809_, _16808_, _06130_);
  or (_16810_, _16809_, _16806_);
  and (_16811_, _15194_, _07698_);
  or (_16812_, _16716_, _08777_);
  or (_16813_, _16812_, _16811_);
  and (_16814_, _16813_, _08782_);
  and (_16815_, _16814_, _16810_);
  nor (_16816_, _10982_, _09258_);
  or (_16817_, _16816_, _16716_);
  and (_16818_, _16817_, _06292_);
  or (_16819_, _16818_, _06316_);
  or (_16820_, _16819_, _16815_);
  or (_16821_, _16725_, _06718_);
  and (_16822_, _16821_, _05653_);
  and (_16823_, _16822_, _16820_);
  and (_16824_, _16722_, _05652_);
  or (_16825_, _16824_, _06047_);
  or (_16826_, _16825_, _16823_);
  and (_16827_, _15253_, _07698_);
  or (_16828_, _16716_, _06048_);
  or (_16829_, _16828_, _16827_);
  and (_16830_, _16829_, _01336_);
  and (_16831_, _16830_, _16826_);
  or (_16832_, _16831_, _16715_);
  and (_43329_, _16832_, _42882_);
  nor (_16833_, _01336_, _10089_);
  nor (_16834_, _07698_, _10089_);
  and (_16835_, _15389_, _07698_);
  or (_16836_, _16835_, _16834_);
  or (_16837_, _16836_, _06020_);
  and (_16838_, _15382_, _07698_);
  or (_16839_, _16838_, _16834_);
  and (_16840_, _16839_, _09833_);
  nor (_16841_, _08361_, _10089_);
  and (_16842_, _15278_, _08361_);
  or (_16843_, _16842_, _16841_);
  and (_16844_, _16843_, _06039_);
  and (_16845_, _15293_, _07698_);
  or (_16846_, _16845_, _16834_);
  or (_16847_, _16846_, _06954_);
  and (_16848_, _07698_, \oc8051_golden_model_1.ACC [6]);
  or (_16849_, _16848_, _16834_);
  and (_16850_, _16849_, _06938_);
  nor (_16851_, _06938_, _10089_);
  or (_16852_, _16851_, _06102_);
  or (_16853_, _16852_, _16850_);
  and (_16854_, _16853_, _06044_);
  and (_16855_, _16854_, _16847_);
  and (_16856_, _15280_, _08361_);
  or (_16857_, _16856_, _16841_);
  and (_16858_, _16857_, _06043_);
  or (_16859_, _16858_, _06239_);
  or (_16860_, _16859_, _16855_);
  nor (_16861_, _07883_, _09258_);
  or (_16862_, _16861_, _16834_);
  or (_16863_, _16862_, _06848_);
  and (_16864_, _16863_, _16860_);
  or (_16865_, _16864_, _06219_);
  or (_16866_, _16849_, _06220_);
  and (_16867_, _16866_, _06040_);
  and (_16868_, _16867_, _16865_);
  or (_16869_, _16868_, _16844_);
  and (_16870_, _16869_, _06033_);
  or (_16871_, _16841_, _15310_);
  and (_16872_, _16857_, _06032_);
  and (_16873_, _16872_, _16871_);
  or (_16874_, _16873_, _09269_);
  or (_16875_, _16874_, _16870_);
  not (_16876_, _09799_);
  or (_16877_, _09797_, _09781_);
  and (_16878_, _16877_, _16876_);
  or (_16879_, _16878_, _09800_);
  and (_16880_, _16879_, _06027_);
  and (_16881_, _16880_, _16875_);
  or (_16882_, _16841_, _15326_);
  and (_16883_, _16882_, _06026_);
  and (_16884_, _16883_, _16857_);
  or (_16885_, _16884_, _09818_);
  or (_16886_, _16885_, _16881_);
  and (_16887_, _09178_, _07698_);
  or (_16888_, _16834_, _07012_);
  or (_16889_, _16888_, _16887_);
  or (_16890_, _16862_, _09827_);
  and (_16891_, _16890_, _05669_);
  and (_16892_, _16891_, _16889_);
  and (_16893_, _16892_, _16886_);
  or (_16894_, _16893_, _16840_);
  and (_16895_, _16894_, _09839_);
  nor (_16896_, _16778_, _10158_);
  or (_16897_, _16896_, _10159_);
  nor (_16898_, _16897_, _10164_);
  and (_16899_, _16897_, _10164_);
  or (_16900_, _16899_, _16898_);
  or (_16901_, _16900_, _10184_);
  nor (_16902_, _10102_, _09839_);
  or (_16903_, _16902_, _16782_);
  and (_16904_, _16903_, _16901_);
  or (_16905_, _16904_, _06019_);
  or (_16906_, _16905_, _16895_);
  and (_16907_, _16906_, _16837_);
  or (_16908_, _16907_, _06112_);
  and (_16909_, _15399_, _07698_);
  or (_16910_, _16909_, _16834_);
  or (_16911_, _16910_, _08751_);
  and (_16912_, _16911_, _08756_);
  and (_16913_, _16912_, _16908_);
  and (_16914_, _10980_, _07698_);
  or (_16915_, _16914_, _16834_);
  and (_16916_, _16915_, _06284_);
  or (_16917_, _16916_, _16913_);
  and (_16918_, _16917_, _07032_);
  or (_16919_, _16834_, _07886_);
  and (_16920_, _16836_, _06108_);
  and (_16921_, _16920_, _16919_);
  or (_16922_, _16921_, _16918_);
  and (_16923_, _16922_, _06278_);
  and (_16924_, _16849_, _06277_);
  and (_16925_, _16924_, _16919_);
  or (_16926_, _16925_, _06130_);
  or (_16927_, _16926_, _16923_);
  and (_16928_, _15396_, _07698_);
  or (_16929_, _16834_, _08777_);
  or (_16930_, _16929_, _16928_);
  and (_16931_, _16930_, _08782_);
  and (_16932_, _16931_, _16927_);
  nor (_16933_, _10979_, _09258_);
  or (_16934_, _16933_, _16834_);
  and (_16935_, _16934_, _06292_);
  or (_16936_, _16935_, _06316_);
  or (_16937_, _16936_, _16932_);
  or (_16938_, _16846_, _06718_);
  and (_16939_, _16938_, _05653_);
  and (_16940_, _16939_, _16937_);
  and (_16941_, _16843_, _05652_);
  or (_16942_, _16941_, _06047_);
  or (_16943_, _16942_, _16940_);
  and (_16944_, _15451_, _07698_);
  or (_16945_, _16834_, _06048_);
  or (_16946_, _16945_, _16944_);
  and (_16947_, _16946_, _01336_);
  and (_16948_, _16947_, _16943_);
  or (_16949_, _16948_, _16833_);
  and (_43330_, _16949_, _42882_);
  nor (_16950_, _01336_, _05758_);
  nand (_16951_, _11015_, _08393_);
  nand (_16952_, _12303_, _06051_);
  and (_16953_, _16952_, _11050_);
  nor (_16954_, _06931_, \oc8051_golden_model_1.ACC [0]);
  nor (_16955_, _10913_, _16954_);
  not (_16956_, _10890_);
  and (_16957_, _16956_, _16955_);
  nor (_16958_, _10285_, _05758_);
  or (_16959_, _16958_, _10477_);
  or (_16960_, _10794_, _16959_);
  and (_16961_, _16960_, _12525_);
  nand (_16962_, _10781_, _12321_);
  and (_16963_, _14086_, _07701_);
  nor (_16964_, _07701_, _05758_);
  or (_16965_, _16964_, _08751_);
  or (_16966_, _16965_, _16963_);
  nor (_16967_, _09120_, \oc8051_golden_model_1.ACC [0]);
  nor (_16968_, _10955_, _16967_);
  or (_16969_, _10686_, _16968_);
  not (_16970_, _06650_);
  and (_16971_, _06133_, _05726_);
  not (_16972_, _16971_);
  and (_16973_, _10677_, _16955_);
  nor (_16974_, _12322_, _10606_);
  and (_16975_, _12322_, _10606_);
  or (_16976_, _16975_, _16974_);
  or (_16977_, _16976_, _10307_);
  not (_16978_, _10378_);
  or (_16979_, _16978_, _06931_);
  or (_16980_, _10400_, _06931_);
  nor (_16981_, _06530_, _05758_);
  and (_16982_, _06530_, _05758_);
  nor (_16983_, _16982_, _16981_);
  nand (_16984_, _16983_, _10400_);
  and (_16985_, _16984_, _10390_);
  and (_16986_, _16985_, _16980_);
  and (_16987_, _16986_, _06949_);
  or (_16988_, _16987_, _09120_);
  or (_16989_, _16986_, _10389_);
  and (_16990_, _16989_, _05698_);
  or (_16991_, _16990_, _06948_);
  and (_16992_, _16991_, _06954_);
  and (_16993_, _16992_, _16988_);
  nor (_16994_, _08127_, _10439_);
  or (_16995_, _16994_, _16964_);
  and (_16996_, _16995_, _06102_);
  or (_16997_, _16996_, _06043_);
  or (_16998_, _16997_, _16993_);
  and (_16999_, _14102_, _08359_);
  nor (_17000_, _08359_, _05758_);
  or (_17001_, _17000_, _06044_);
  or (_17002_, _17001_, _16999_);
  and (_17003_, _17002_, _06848_);
  and (_17004_, _17003_, _16998_);
  and (_17005_, _07701_, _06931_);
  or (_17006_, _17005_, _16964_);
  and (_17007_, _17006_, _06239_);
  or (_17008_, _17007_, _10378_);
  or (_17009_, _17008_, _17004_);
  and (_17010_, _17009_, _16979_);
  or (_17011_, _17010_, _06970_);
  or (_17012_, _09120_, _06971_);
  and (_17013_, _17012_, _06220_);
  and (_17014_, _17013_, _17011_);
  and (_17015_, _08127_, _06219_);
  or (_17016_, _17015_, _10376_);
  or (_17017_, _17016_, _17014_);
  nand (_17018_, _10376_, _09880_);
  and (_17019_, _17018_, _17017_);
  or (_17020_, _17019_, _06039_);
  or (_17021_, _16964_, _06040_);
  and (_17022_, _17021_, _06033_);
  and (_17023_, _17022_, _17020_);
  and (_17024_, _16995_, _06032_);
  or (_17025_, _17024_, _09269_);
  or (_17026_, _17025_, _17023_);
  nand (_17027_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nand (_17028_, _17027_, _09269_);
  and (_17029_, _17028_, _10469_);
  and (_17030_, _17029_, _17026_);
  and (_17031_, _16959_, _10468_);
  or (_17032_, _17031_, _12361_);
  or (_17033_, _17032_, _17030_);
  nor (_17034_, _10542_, _05758_);
  or (_17035_, _17034_, _10543_);
  or (_17036_, _17035_, _13935_);
  and (_17037_, _17036_, _06267_);
  and (_17038_, _17037_, _17033_);
  nor (_17039_, _10353_, _05758_);
  or (_17040_, _17039_, _10354_);
  or (_17041_, _17040_, _10306_);
  and (_17042_, _17041_, _12367_);
  or (_17043_, _17042_, _17038_);
  and (_17044_, _17043_, _16977_);
  or (_17045_, _17044_, _05676_);
  nand (_17046_, _06016_, _05676_);
  and (_17047_, _17046_, _06027_);
  and (_17048_, _17047_, _17045_);
  and (_17049_, _14132_, _08359_);
  or (_17050_, _17049_, _17000_);
  and (_17051_, _17050_, _06026_);
  or (_17052_, _17051_, _09818_);
  or (_17053_, _17052_, _17048_);
  and (_17054_, _09120_, _07701_);
  or (_17055_, _16964_, _07012_);
  or (_17056_, _17055_, _17054_);
  or (_17057_, _17006_, _09827_);
  and (_17058_, _17057_, _05669_);
  and (_17059_, _17058_, _17056_);
  and (_17060_, _17059_, _17053_);
  and (_17061_, _14186_, _07701_);
  or (_17062_, _17061_, _16964_);
  and (_17063_, _17062_, _09833_);
  or (_17064_, _17063_, _09832_);
  or (_17065_, _17064_, _17060_);
  nor (_17066_, _16775_, _05663_);
  and (_17067_, _17066_, _17065_);
  nor (_17068_, _06016_, _05664_);
  or (_17069_, _17068_, _06019_);
  or (_17070_, _17069_, _17067_);
  and (_17071_, _07701_, _08672_);
  or (_17072_, _17071_, _16964_);
  or (_17073_, _17072_, _06020_);
  and (_17074_, _17073_, _10662_);
  and (_17075_, _17074_, _17070_);
  nor (_17076_, _10662_, _06016_);
  or (_17077_, _17076_, _10669_);
  or (_17078_, _17077_, _17075_);
  or (_17079_, _10675_, _16955_);
  and (_17080_, _17079_, _10678_);
  and (_17081_, _17080_, _17078_);
  or (_17082_, _17081_, _16973_);
  and (_17083_, _17082_, _16972_);
  and (_17084_, _16971_, _16955_);
  or (_17085_, _17084_, _17083_);
  and (_17086_, _17085_, _16970_);
  and (_17087_, _16955_, _06650_);
  or (_17088_, _17087_, _10685_);
  or (_17089_, _17088_, _17086_);
  and (_17090_, _17089_, _16969_);
  or (_17091_, _17090_, _06282_);
  nand (_17092_, _12303_, _06282_);
  and (_17093_, _17092_, _10699_);
  and (_17094_, _17093_, _17091_);
  and (_17095_, _10698_, _12322_);
  or (_17096_, _17095_, _06112_);
  or (_17097_, _17096_, _17094_);
  and (_17098_, _17097_, _16966_);
  or (_17099_, _17098_, _06284_);
  or (_17100_, _16964_, _08756_);
  nand (_17101_, _05735_, _05567_);
  and (_17102_, _17101_, _17100_);
  and (_17103_, _17102_, _17099_);
  not (_17104_, _17101_);
  and (_17105_, _17104_, _10913_);
  or (_17106_, _17105_, _10731_);
  or (_17107_, _17106_, _17103_);
  or (_17108_, _10736_, _10955_);
  and (_17109_, _17108_, _10735_);
  and (_17110_, _17109_, _17107_);
  or (_17111_, _10741_, _10995_);
  and (_17112_, _17111_, _10743_);
  or (_17113_, _17112_, _17110_);
  or (_17114_, _10747_, _11036_);
  and (_17115_, _17114_, _07032_);
  and (_17116_, _17115_, _17113_);
  nand (_17117_, _17072_, _06108_);
  nor (_17118_, _17117_, _16994_);
  or (_17119_, _17118_, _10752_);
  or (_17120_, _17119_, _17116_);
  nand (_17121_, _16954_, _10752_);
  and (_17122_, _17121_, _10760_);
  and (_17123_, _17122_, _17120_);
  nor (_17124_, _10760_, _16954_);
  or (_17125_, _17124_, _10767_);
  or (_17126_, _17125_, _17123_);
  nand (_17127_, _10767_, _16954_);
  and (_17128_, _17127_, _06668_);
  and (_17129_, _17128_, _17126_);
  nor (_17130_, _16954_, _06668_);
  or (_17131_, _17130_, _10775_);
  or (_17132_, _17131_, _17129_);
  nand (_17133_, _10775_, _16967_);
  and (_17134_, _17133_, _06291_);
  and (_17135_, _17134_, _17132_);
  not (_17136_, _10781_);
  nand (_17137_, _17136_, _12302_);
  and (_17138_, _17137_, _11987_);
  or (_17139_, _17138_, _17135_);
  and (_17140_, _17139_, _16962_);
  or (_17141_, _17140_, _06130_);
  and (_17142_, _14083_, _07701_);
  or (_17143_, _16964_, _08777_);
  or (_17144_, _17143_, _17142_);
  and (_17145_, _17144_, _10304_);
  and (_17146_, _17145_, _17141_);
  or (_17147_, _17146_, _16961_);
  or (_17148_, _10796_, _17035_);
  and (_17149_, _17148_, _17147_);
  or (_17150_, _17149_, _06288_);
  or (_17151_, _17040_, _06289_);
  and (_17152_, _17151_, _10856_);
  and (_17153_, _17152_, _17150_);
  and (_17154_, _10824_, _16976_);
  or (_17155_, _17154_, _10854_);
  or (_17156_, _17155_, _17153_);
  nand (_17157_, _10854_, _10606_);
  and (_17158_, _17157_, _10890_);
  and (_17159_, _17158_, _17156_);
  or (_17160_, _17159_, _16957_);
  and (_17161_, _17160_, _10934_);
  and (_17162_, _10932_, _16968_);
  or (_17163_, _17162_, _06051_);
  or (_17164_, _17163_, _17161_);
  and (_17165_, _17164_, _16953_);
  and (_17166_, _10974_, _12322_);
  or (_17167_, _17166_, _11015_);
  or (_17168_, _17167_, _17165_);
  and (_17169_, _17168_, _16951_);
  or (_17170_, _17169_, _06316_);
  or (_17171_, _16995_, _06718_);
  and (_17172_, _17171_, _11060_);
  and (_17173_, _17172_, _17170_);
  nor (_17174_, _11064_, _05758_);
  nor (_17175_, _17174_, _12756_);
  or (_17176_, _17175_, _17173_);
  nand (_17177_, _11064_, _05784_);
  and (_17178_, _17177_, _05653_);
  and (_17179_, _17178_, _17176_);
  and (_17180_, _16964_, _05652_);
  or (_17181_, _17180_, _06047_);
  or (_17182_, _17181_, _17179_);
  or (_17183_, _16995_, _06048_);
  and (_17184_, _17183_, _11083_);
  and (_17185_, _17184_, _17182_);
  nor (_17186_, _11089_, _05758_);
  nor (_17187_, _17186_, _12779_);
  or (_17188_, _17187_, _17185_);
  nand (_17189_, _11089_, _05784_);
  and (_17190_, _17189_, _01336_);
  and (_17191_, _17190_, _17188_);
  or (_17192_, _17191_, _16950_);
  and (_43332_, _17192_, _42882_);
  nor (_17193_, _01336_, _05784_);
  nor (_17194_, _10835_, _10834_);
  nor (_17195_, _17194_, _10836_);
  or (_17196_, _17195_, _06289_);
  and (_17197_, _17196_, _10856_);
  and (_17198_, _07701_, _06832_);
  and (_17199_, _17198_, _08077_);
  nor (_17200_, _07701_, \oc8051_golden_model_1.ACC [1]);
  or (_17201_, _17200_, _08777_);
  or (_17202_, _17201_, _17199_);
  and (_17203_, _06460_, _05739_);
  nor (_17204_, _06834_, _17203_);
  not (_17205_, _10752_);
  or (_17206_, _10736_, _10951_);
  nor (_17207_, _10677_, _10669_);
  not (_17208_, _17207_);
  and (_17209_, _17208_, _10912_);
  or (_17210_, _10092_, _09839_);
  not (_17211_, _10954_);
  nor (_17212_, _10536_, _05758_);
  or (_17213_, _17212_, _10541_);
  nand (_17214_, _17213_, _17211_);
  or (_17215_, _17213_, _17211_);
  and (_17216_, _17215_, _12361_);
  and (_17217_, _17216_, _17214_);
  nand (_17218_, _10378_, _07132_);
  nor (_17219_, _10389_, _06948_);
  or (_17220_, _17219_, _09075_);
  nor (_17221_, _10400_, _07132_);
  nor (_17222_, _06530_, _05784_);
  and (_17223_, _06530_, _05784_);
  or (_17224_, _17223_, _17222_);
  and (_17225_, _17224_, _10400_);
  or (_17226_, _17225_, _10389_);
  or (_17227_, _17226_, _17221_);
  and (_17228_, _17227_, _05698_);
  or (_17229_, _17228_, _06948_);
  and (_17230_, _17229_, _06954_);
  and (_17231_, _17230_, _17220_);
  and (_17232_, _14284_, _07701_);
  nor (_17233_, _17232_, _17200_);
  and (_17234_, _17233_, _06102_);
  or (_17235_, _17234_, _10412_);
  or (_17236_, _17235_, _17231_);
  nor (_17237_, _10416_, \oc8051_golden_model_1.PSW [6]);
  nor (_17238_, _17237_, \oc8051_golden_model_1.ACC [1]);
  and (_17239_, _17237_, \oc8051_golden_model_1.ACC [1]);
  nor (_17240_, _17239_, _17238_);
  nand (_17241_, _17240_, _10412_);
  and (_17242_, _17241_, _06244_);
  and (_17243_, _17242_, _17236_);
  nor (_17244_, _08359_, _05784_);
  and (_17245_, _14266_, _08359_);
  nor (_17246_, _17245_, _17244_);
  nor (_17247_, _17246_, _06044_);
  nor (_17248_, _07701_, _05784_);
  nor (_17249_, _10439_, _07132_);
  or (_17250_, _17249_, _17248_);
  and (_17251_, _17250_, _06239_);
  or (_17252_, _17251_, _10378_);
  or (_17253_, _17252_, _17247_);
  or (_17254_, _17253_, _17243_);
  and (_17255_, _17254_, _17218_);
  or (_17256_, _17255_, _06970_);
  or (_17257_, _09075_, _06971_);
  and (_17258_, _17257_, _06220_);
  and (_17259_, _17258_, _17256_);
  nor (_17260_, _08077_, _06220_);
  or (_17261_, _17260_, _10376_);
  or (_17262_, _17261_, _17259_);
  nand (_17263_, _10376_, _09906_);
  and (_17264_, _17263_, _17262_);
  or (_17265_, _17264_, _06039_);
  and (_17266_, _14273_, _08359_);
  or (_17267_, _17266_, _17244_);
  or (_17268_, _17267_, _06040_);
  and (_17269_, _17268_, _06033_);
  nand (_17270_, _17269_, _17265_);
  nor (_17271_, _17244_, _14302_);
  or (_17272_, _17246_, _06033_);
  or (_17273_, _17272_, _17271_);
  and (_17274_, _17273_, _17270_);
  nor (_17275_, _17274_, _09269_);
  nor (_17276_, _09744_, _09743_);
  nor (_17277_, _17276_, _09745_);
  nand (_17278_, _17277_, _09269_);
  nand (_17279_, _17278_, _10469_);
  or (_17280_, _17279_, _17275_);
  nor (_17281_, _10234_, _05758_);
  or (_17282_, _17281_, _10284_);
  nor (_17283_, _17282_, _10912_);
  and (_17284_, _17282_, _10912_);
  or (_17285_, _17284_, _17283_);
  or (_17286_, _17285_, _10469_);
  and (_17287_, _17286_, _13935_);
  and (_17288_, _17287_, _17280_);
  or (_17289_, _17288_, _17217_);
  and (_17290_, _17289_, _06267_);
  nor (_17291_, _10308_, _05758_);
  or (_17292_, _17291_, _10352_);
  and (_17293_, _17292_, _10994_);
  nor (_17294_, _17292_, _10994_);
  or (_17295_, _17294_, _17293_);
  and (_17296_, _17295_, _06261_);
  or (_17297_, _17296_, _17290_);
  and (_17298_, _17297_, _10307_);
  nor (_17299_, _06016_, \oc8051_golden_model_1.ACC [0]);
  nor (_17300_, _17299_, _11035_);
  and (_17301_, _17299_, _11035_);
  or (_17302_, _17301_, _17300_);
  nor (_17303_, _16974_, _17302_);
  and (_17304_, _12323_, \oc8051_golden_model_1.PSW [7]);
  or (_17305_, _17304_, _17303_);
  and (_17306_, _17305_, _10306_);
  or (_17307_, _17306_, _05676_);
  or (_17308_, _17307_, _17298_);
  nand (_17309_, _06799_, _05676_);
  and (_17310_, _17309_, _06027_);
  and (_17311_, _17310_, _17308_);
  or (_17312_, _17244_, _14267_);
  nand (_17313_, _17312_, _06026_);
  nor (_17314_, _17313_, _17246_);
  or (_17315_, _17314_, _09818_);
  or (_17316_, _17315_, _17311_);
  and (_17317_, _09075_, _07701_);
  or (_17318_, _17248_, _07012_);
  or (_17319_, _17318_, _17317_);
  or (_17320_, _17250_, _09827_);
  and (_17321_, _17320_, _05669_);
  and (_17322_, _17321_, _17319_);
  and (_17323_, _17322_, _17316_);
  or (_17324_, _14367_, _10439_);
  nor (_17325_, _17200_, _05669_);
  and (_17326_, _17325_, _17324_);
  or (_17327_, _17326_, _09832_);
  or (_17328_, _17327_, _17323_);
  and (_17329_, _17328_, _17210_);
  or (_17330_, _17329_, _05663_);
  nand (_17331_, _06799_, _05663_);
  and (_17332_, _17331_, _06020_);
  and (_17333_, _17332_, _17330_);
  or (_17334_, _17198_, _06020_);
  nor (_17335_, _17334_, _17200_);
  or (_17336_, _17335_, _10661_);
  or (_17337_, _17336_, _17333_);
  nand (_17338_, _10661_, _06799_);
  and (_17339_, _17338_, _17207_);
  and (_17340_, _17339_, _17337_);
  or (_17341_, _17340_, _17209_);
  and (_17342_, _17341_, _16972_);
  and (_17343_, _16971_, _10912_);
  or (_17344_, _17343_, _17342_);
  and (_17345_, _17344_, _16970_);
  and (_17346_, _10912_, _06650_);
  or (_17347_, _17346_, _17345_);
  and (_17348_, _17347_, _10686_);
  and (_17349_, _10685_, _10954_);
  or (_17350_, _17349_, _06282_);
  or (_17351_, _17350_, _17348_);
  or (_17352_, _10994_, _06283_);
  and (_17353_, _17352_, _10699_);
  and (_17354_, _17353_, _17351_);
  and (_17355_, _10698_, _11035_);
  or (_17356_, _17355_, _17354_);
  and (_17357_, _17356_, _08751_);
  or (_17358_, _14263_, _10439_);
  nor (_17359_, _17200_, _08751_);
  and (_17360_, _17359_, _17358_);
  or (_17361_, _17360_, _06284_);
  or (_17362_, _17361_, _17357_);
  or (_17363_, _17248_, _08756_);
  and (_17364_, _17363_, _17101_);
  and (_17365_, _17364_, _17362_);
  and (_17366_, _17104_, _10910_);
  or (_17367_, _17366_, _10731_);
  or (_17368_, _17367_, _17365_);
  and (_17369_, _17368_, _17206_);
  or (_17370_, _17369_, _06279_);
  or (_17371_, _10992_, _10735_);
  and (_17372_, _17371_, _10747_);
  and (_17373_, _17372_, _17370_);
  and (_17375_, _10741_, _11033_);
  or (_17376_, _17375_, _17373_);
  and (_17377_, _17376_, _07032_);
  or (_17378_, _14261_, _10439_);
  nor (_17379_, _17200_, _07032_);
  and (_17380_, _17379_, _17378_);
  or (_17381_, _17380_, _17377_);
  and (_17382_, _17381_, _17205_);
  nor (_17383_, _10911_, _17205_);
  nor (_17384_, _17383_, _17382_);
  nand (_17386_, _17384_, _17204_);
  not (_17387_, _11991_);
  not (_17388_, _17204_);
  nand (_17389_, _17388_, _10911_);
  and (_17390_, _17389_, _17387_);
  and (_17391_, _17390_, _17386_);
  nor (_17392_, _17387_, _10911_);
  or (_17393_, _17392_, _10775_);
  or (_17394_, _17393_, _17391_);
  not (_17395_, _10775_);
  or (_17397_, _17395_, _10952_);
  and (_17398_, _17397_, _06291_);
  and (_17399_, _17398_, _17394_);
  nor (_17400_, _10993_, _06291_);
  or (_17401_, _17400_, _10781_);
  or (_17402_, _17401_, _17399_);
  nand (_17403_, _10781_, _11034_);
  and (_17404_, _17403_, _08777_);
  nand (_17405_, _17404_, _17402_);
  and (_17406_, _17405_, _17202_);
  or (_17408_, _17406_, _10303_);
  and (_17409_, _10794_, _06545_);
  not (_17410_, _17409_);
  and (_17411_, _10287_, _10283_);
  or (_17412_, _10304_, _10288_);
  or (_17413_, _17412_, _17411_);
  and (_17414_, _17413_, _17410_);
  and (_17415_, _17414_, _17408_);
  and (_17416_, _06513_, _05731_);
  and (_17417_, _10805_, _10803_);
  or (_17419_, _17417_, _10806_);
  and (_17420_, _17419_, _17409_);
  or (_17421_, _17420_, _17416_);
  nor (_17422_, _17421_, _17415_);
  not (_17423_, _17416_);
  or (_17424_, _17419_, _17423_);
  nand (_17425_, _17424_, _06289_);
  or (_17426_, _17425_, _17422_);
  and (_17427_, _17426_, _17197_);
  or (_17428_, _10865_, _10864_);
  nor (_17430_, _10866_, _10856_);
  and (_17431_, _17430_, _17428_);
  or (_17432_, _17431_, _10854_);
  or (_17433_, _17432_, _17427_);
  nand (_17434_, _10854_, _05758_);
  and (_17435_, _17434_, _10890_);
  and (_17436_, _17435_, _17433_);
  and (_17437_, _10394_, _05746_);
  or (_17438_, _10913_, _10912_);
  nor (_17439_, _10914_, _10890_);
  and (_17440_, _17439_, _17438_);
  or (_17441_, _17440_, _17437_);
  or (_17442_, _17441_, _17436_);
  not (_17443_, _06692_);
  nor (_17444_, _10955_, _10954_);
  nor (_17445_, _17444_, _10956_);
  and (_17446_, _17445_, _17443_);
  or (_17447_, _17446_, _10934_);
  and (_17448_, _17447_, _17442_);
  and (_17449_, _17445_, _06692_);
  or (_17450_, _17449_, _10976_);
  or (_17451_, _17450_, _17448_);
  nor (_17452_, _10995_, _10994_);
  nor (_17453_, _17452_, _10996_);
  or (_17454_, _17453_, _06052_);
  nor (_17455_, _11036_, _11035_);
  nor (_17456_, _17455_, _11037_);
  or (_17457_, _17456_, _11050_);
  and (_17458_, _17457_, _11016_);
  and (_17459_, _17458_, _17454_);
  and (_17460_, _17459_, _17451_);
  and (_17461_, _11015_, \oc8051_golden_model_1.ACC [0]);
  or (_17462_, _17461_, _06316_);
  or (_17463_, _17462_, _17460_);
  or (_17464_, _17233_, _06718_);
  and (_17465_, _17464_, _11060_);
  and (_17466_, _17465_, _17463_);
  nor (_17467_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  nor (_17468_, _11090_, _17467_);
  nor (_17469_, _17468_, _11060_);
  or (_17470_, _17469_, _11064_);
  or (_17471_, _17470_, _17466_);
  nand (_17472_, _11064_, _09956_);
  and (_17473_, _17472_, _05653_);
  and (_17474_, _17473_, _17471_);
  and (_17475_, _17267_, _05652_);
  or (_17476_, _17475_, _06047_);
  or (_17477_, _17476_, _17474_);
  or (_17478_, _17232_, _17248_);
  or (_17479_, _17478_, _06048_);
  and (_17480_, _17479_, _11083_);
  and (_17481_, _17480_, _17477_);
  and (_17482_, _17468_, _11082_);
  or (_17483_, _17482_, _11089_);
  or (_17484_, _17483_, _17481_);
  nand (_17485_, _11089_, _09956_);
  and (_17486_, _17485_, _01336_);
  and (_17487_, _17486_, _17484_);
  or (_17488_, _17487_, _17193_);
  and (_43333_, _17488_, _42882_);
  nor (_17489_, _01336_, _09956_);
  nand (_17490_, _11015_, _05784_);
  nor (_17491_, _10998_, _10991_);
  nor (_17492_, _17491_, _10999_);
  or (_17493_, _17492_, _06052_);
  and (_17494_, _17493_, _11050_);
  and (_17495_, _10837_, _10346_);
  nor (_17496_, _17495_, _10838_);
  or (_17497_, _17496_, _06289_);
  and (_17498_, _17497_, _10856_);
  and (_17499_, _14596_, _07701_);
  nor (_17500_, _07701_, _09956_);
  or (_17501_, _17500_, _08751_);
  or (_17502_, _17501_, _17499_);
  and (_17503_, _06227_, _05726_);
  and (_17504_, _10909_, _17503_);
  nand (_17505_, _10378_, _07530_);
  or (_17506_, _17219_, _09182_);
  nor (_17507_, _10400_, _07530_);
  nor (_17508_, _06530_, _09956_);
  and (_17509_, _06530_, _09956_);
  or (_17510_, _17509_, _17508_);
  and (_17511_, _17510_, _10400_);
  or (_17512_, _17511_, _10389_);
  or (_17513_, _17512_, _17507_);
  and (_17514_, _17513_, _05698_);
  or (_17515_, _17514_, _06948_);
  and (_17516_, _17515_, _06954_);
  and (_17517_, _17516_, _17506_);
  and (_17518_, _14493_, _07701_);
  or (_17519_, _17518_, _17500_);
  and (_17520_, _17519_, _06102_);
  or (_17521_, _17520_, _10412_);
  or (_17522_, _17521_, _17517_);
  nor (_17523_, _17238_, _09956_);
  and (_17524_, _10415_, \oc8051_golden_model_1.PSW [6]);
  nor (_17525_, _17524_, _17523_);
  nand (_17526_, _17525_, _10412_);
  and (_17527_, _17526_, _06244_);
  and (_17528_, _17527_, _17522_);
  nor (_17529_, _08359_, _09956_);
  and (_17530_, _14497_, _08359_);
  or (_17531_, _17530_, _17529_);
  and (_17532_, _17531_, _06043_);
  nor (_17533_, _10439_, _07530_);
  or (_17534_, _17533_, _17500_);
  and (_17535_, _17534_, _06239_);
  or (_17536_, _17535_, _10378_);
  or (_17537_, _17536_, _17532_);
  or (_17538_, _17537_, _17528_);
  and (_17539_, _17538_, _17505_);
  or (_17540_, _17539_, _06970_);
  or (_17541_, _09182_, _06971_);
  and (_17542_, _17541_, _06220_);
  and (_17543_, _17542_, _17540_);
  nor (_17544_, _08176_, _06220_);
  or (_17545_, _17544_, _10376_);
  or (_17546_, _17545_, _17543_);
  nand (_17547_, _10376_, _09861_);
  and (_17548_, _17547_, _17546_);
  or (_17549_, _17548_, _06039_);
  and (_17550_, _14479_, _08359_);
  or (_17551_, _17550_, _17529_);
  or (_17552_, _17551_, _06040_);
  and (_17553_, _17552_, _06033_);
  and (_17554_, _17553_, _17549_);
  or (_17555_, _17529_, _14512_);
  and (_17556_, _17531_, _06032_);
  and (_17557_, _17556_, _17555_);
  or (_17558_, _17557_, _09269_);
  or (_17559_, _17558_, _17554_);
  nor (_17560_, _09747_, _09745_);
  or (_17561_, _17560_, _09748_);
  nand (_17562_, _17561_, _09269_);
  and (_17563_, _17562_, _10469_);
  and (_17564_, _17563_, _17559_);
  and (_17565_, _07132_, \oc8051_golden_model_1.ACC [1]);
  and (_17566_, _06931_, _05758_);
  nor (_17567_, _17566_, _10912_);
  nor (_17568_, _17567_, _17565_);
  nor (_17569_, _10909_, _17568_);
  and (_17570_, _10909_, _17568_);
  nor (_17571_, _17570_, _17569_);
  nor (_17572_, _16955_, _10912_);
  and (_17573_, _17572_, \oc8051_golden_model_1.PSW [7]);
  or (_17574_, _17573_, _17571_);
  nand (_17575_, _17573_, _17571_);
  and (_17576_, _17575_, _10468_);
  and (_17577_, _17576_, _17574_);
  or (_17578_, _17577_, _12361_);
  or (_17579_, _17578_, _17564_);
  and (_17580_, _12150_, \oc8051_golden_model_1.ACC [1]);
  not (_17581_, _17580_);
  and (_17582_, _09120_, _05758_);
  or (_17583_, _17582_, _10954_);
  and (_17584_, _17583_, _17581_);
  nor (_17585_, _10949_, _17584_);
  and (_17586_, _10949_, _17584_);
  nor (_17587_, _17586_, _17585_);
  nor (_17588_, _16968_, _10954_);
  not (_17589_, _17588_);
  or (_17590_, _17589_, _17587_);
  and (_17591_, _17590_, \oc8051_golden_model_1.PSW [7]);
  nor (_17592_, _17587_, \oc8051_golden_model_1.PSW [7]);
  nor (_17593_, _17592_, _17591_);
  and (_17594_, _17589_, _17587_);
  or (_17595_, _17594_, _13935_);
  or (_17596_, _17595_, _17593_);
  and (_17597_, _17596_, _06267_);
  and (_17598_, _17597_, _17579_);
  and (_17599_, _08077_, \oc8051_golden_model_1.ACC [1]);
  and (_17600_, _08127_, _05758_);
  nor (_17601_, _17600_, _13785_);
  nor (_17602_, _17601_, _17599_);
  nor (_17603_, _10991_, _17602_);
  and (_17604_, _10991_, _17602_);
  nor (_17605_, _17604_, _17603_);
  and (_17606_, _12304_, \oc8051_golden_model_1.PSW [7]);
  not (_17607_, _17606_);
  and (_17608_, _17607_, _17605_);
  or (_17609_, _17607_, _17605_);
  nand (_17610_, _17609_, _10307_);
  or (_17611_, _17610_, _17608_);
  and (_17612_, _17611_, _12367_);
  or (_17613_, _17612_, _17598_);
  nor (_17614_, _17300_, _13874_);
  nor (_17615_, _12318_, _17614_);
  and (_17616_, _12318_, _17614_);
  nor (_17617_, _17616_, _17615_);
  not (_17618_, _17304_);
  or (_17619_, _17618_, _17617_);
  nand (_17620_, _17618_, _17617_);
  and (_17621_, _17620_, _10306_);
  nand (_17622_, _17621_, _17619_);
  and (_17623_, _17622_, _17613_);
  or (_17624_, _17623_, _05676_);
  nand (_17625_, _06403_, _05676_);
  and (_17626_, _17625_, _06027_);
  and (_17627_, _17626_, _17624_);
  or (_17628_, _17529_, _14525_);
  and (_17629_, _17628_, _06026_);
  and (_17630_, _17629_, _17531_);
  or (_17631_, _17630_, _09818_);
  or (_17632_, _17631_, _17627_);
  and (_17633_, _09182_, _07701_);
  or (_17634_, _17500_, _07012_);
  or (_17635_, _17634_, _17633_);
  or (_17636_, _17534_, _09827_);
  and (_17637_, _17636_, _05669_);
  and (_17638_, _17637_, _17635_);
  and (_17639_, _17638_, _17632_);
  and (_17640_, _14580_, _07701_);
  or (_17641_, _17640_, _17500_);
  and (_17642_, _17641_, _09833_);
  or (_17643_, _17642_, _09832_);
  or (_17644_, _17643_, _17639_);
  or (_17645_, _10028_, _09839_);
  and (_17646_, _17645_, _05664_);
  and (_17647_, _17646_, _17644_);
  nor (_17648_, _06403_, _05664_);
  or (_17649_, _17648_, _06019_);
  or (_17650_, _17649_, _17647_);
  and (_17651_, _07701_, _08730_);
  or (_17652_, _17651_, _17500_);
  or (_17653_, _17652_, _06020_);
  and (_17654_, _17653_, _10662_);
  and (_17655_, _17654_, _17650_);
  and (_17656_, _06094_, _05726_);
  nor (_17657_, _10662_, _06403_);
  or (_17658_, _17657_, _17656_);
  or (_17659_, _17658_, _17655_);
  not (_17660_, _17656_);
  or (_17661_, _10909_, _17660_);
  and (_17662_, _07266_, _05726_);
  not (_17663_, _17662_);
  and (_17664_, _17663_, _17661_);
  and (_17665_, _17664_, _17659_);
  and (_17666_, _06229_, _05726_);
  and (_17667_, _17662_, _10909_);
  or (_17668_, _17667_, _17666_);
  or (_17669_, _17668_, _17665_);
  not (_17670_, _17503_);
  not (_17671_, _17666_);
  or (_17672_, _10909_, _17671_);
  and (_17673_, _17672_, _17670_);
  and (_17674_, _17673_, _17669_);
  or (_17675_, _17674_, _17504_);
  and (_17676_, _17675_, _10687_);
  and (_17677_, _10681_, _10909_);
  or (_17678_, _17677_, _10685_);
  or (_17679_, _17678_, _17676_);
  or (_17680_, _10686_, _10949_);
  and (_17681_, _17680_, _17679_);
  or (_17682_, _17681_, _06282_);
  or (_17683_, _10991_, _06283_);
  and (_17684_, _17683_, _10699_);
  and (_17685_, _17684_, _17682_);
  nor (_17686_, _10699_, _11032_);
  or (_17687_, _17686_, _06112_);
  or (_17688_, _17687_, _17685_);
  and (_17689_, _17688_, _17502_);
  or (_17690_, _17689_, _06284_);
  or (_17691_, _17500_, _08756_);
  and (_17692_, _17691_, _17101_);
  and (_17693_, _17692_, _17690_);
  and (_17694_, _17104_, _10907_);
  or (_17695_, _17694_, _10731_);
  or (_17696_, _17695_, _17693_);
  or (_17697_, _10736_, _10947_);
  and (_17698_, _17697_, _10735_);
  and (_17699_, _17698_, _17696_);
  or (_17700_, _10741_, _10989_);
  and (_17701_, _17700_, _10743_);
  or (_17702_, _17701_, _17699_);
  or (_17703_, _10747_, _11030_);
  and (_17704_, _17703_, _07032_);
  and (_17705_, _17704_, _17702_);
  nand (_17706_, _17652_, _06108_);
  nor (_17707_, _17706_, _10990_);
  or (_17708_, _17707_, _10752_);
  or (_17709_, _17708_, _17705_);
  nand (_17710_, _10908_, _10752_);
  and (_17711_, _17710_, _10760_);
  and (_17712_, _17711_, _17709_);
  nor (_17713_, _10760_, _10908_);
  or (_17714_, _17713_, _10767_);
  or (_17715_, _17714_, _17712_);
  nand (_17716_, _10767_, _10908_);
  and (_17717_, _17716_, _06668_);
  and (_17718_, _17717_, _17715_);
  nor (_17719_, _10908_, _06668_);
  or (_17720_, _17719_, _10775_);
  or (_17721_, _17720_, _17718_);
  nand (_17722_, _10775_, _10948_);
  and (_17723_, _17722_, _06291_);
  and (_17724_, _17723_, _17721_);
  nand (_17725_, _17136_, _10990_);
  and (_17726_, _17725_, _11987_);
  or (_17727_, _17726_, _17724_);
  nand (_17728_, _10781_, _11031_);
  and (_17729_, _17728_, _17727_);
  or (_17730_, _17729_, _06130_);
  and (_17731_, _14593_, _07701_);
  or (_17732_, _17500_, _08777_);
  or (_17733_, _17732_, _17731_);
  and (_17734_, _17733_, _10304_);
  and (_17735_, _17734_, _17730_);
  nand (_17736_, _10289_, _10277_);
  nor (_17737_, _10304_, _10290_);
  and (_17738_, _17737_, _17736_);
  or (_17739_, _17738_, _17409_);
  or (_17740_, _17739_, _17735_);
  and (_17741_, _10807_, _10534_);
  nor (_17742_, _17741_, _10808_);
  or (_17743_, _17742_, _17410_);
  and (_17744_, _17743_, _17423_);
  and (_17745_, _17744_, _17740_);
  nand (_17746_, _17742_, _17416_);
  nand (_17747_, _17746_, _06289_);
  or (_17748_, _17747_, _17745_);
  and (_17749_, _17748_, _17498_);
  nand (_17750_, _10867_, _10604_);
  nor (_17751_, _10868_, _10856_);
  and (_17752_, _17751_, _17750_);
  or (_17753_, _17752_, _10854_);
  or (_17754_, _17753_, _17749_);
  nand (_17755_, _10854_, _05784_);
  and (_17756_, _17755_, _10890_);
  and (_17757_, _17756_, _17754_);
  nor (_17758_, _10916_, _10909_);
  nor (_17759_, _17758_, _10917_);
  and (_17760_, _17759_, _16956_);
  or (_17761_, _17760_, _17437_);
  or (_17762_, _17761_, _17757_);
  and (_17763_, _10957_, _10950_);
  nor (_17764_, _17763_, _10958_);
  and (_17765_, _17764_, _17443_);
  or (_17766_, _17765_, _10934_);
  and (_17767_, _17766_, _17762_);
  and (_17768_, _17764_, _06692_);
  or (_17769_, _17768_, _06051_);
  or (_17770_, _17769_, _17767_);
  and (_17771_, _17770_, _17494_);
  nand (_17772_, _11038_, _11032_);
  nor (_17773_, _11039_, _11050_);
  and (_17774_, _17773_, _17772_);
  or (_17775_, _17774_, _11015_);
  or (_17776_, _17775_, _17771_);
  and (_17777_, _17776_, _17490_);
  or (_17778_, _17777_, _06316_);
  or (_17779_, _17519_, _06718_);
  and (_17780_, _17779_, _11060_);
  and (_17781_, _17780_, _17778_);
  nor (_17782_, _17467_, _09956_);
  or (_17783_, _17782_, _11065_);
  nor (_17784_, _17783_, _11064_);
  nor (_17785_, _17784_, _12756_);
  or (_17786_, _17785_, _17781_);
  nand (_17787_, _11064_, _10010_);
  and (_17788_, _17787_, _05653_);
  and (_17789_, _17788_, _17786_);
  and (_17790_, _17551_, _05652_);
  or (_17791_, _17790_, _06047_);
  or (_17792_, _17791_, _17789_);
  and (_17793_, _14657_, _07701_);
  or (_17794_, _17793_, _17500_);
  or (_17795_, _17794_, _06048_);
  and (_17796_, _17795_, _11083_);
  and (_17797_, _17796_, _17792_);
  nor (_17798_, _11090_, \oc8051_golden_model_1.ACC [2]);
  nor (_17799_, _17798_, _11091_);
  and (_17800_, _17799_, _11082_);
  or (_17801_, _17800_, _11089_);
  or (_17802_, _17801_, _17797_);
  nand (_17803_, _11089_, _10010_);
  and (_17804_, _17803_, _01336_);
  and (_17805_, _17804_, _17802_);
  or (_17806_, _17805_, _17489_);
  and (_43334_, _17806_, _42882_);
  nor (_17807_, _01336_, _10010_);
  and (_17808_, _10291_, _10271_);
  nor (_17809_, _17808_, _10292_);
  or (_17810_, _17809_, _10304_);
  nor (_17811_, _17387_, _10906_);
  or (_17812_, _17811_, _10775_);
  nand (_17813_, _10906_, _06477_);
  or (_17814_, _10987_, _10735_);
  and (_17815_, _17814_, _10747_);
  and (_17816_, _14793_, _07701_);
  nor (_17817_, _07701_, _10010_);
  or (_17818_, _17817_, _08751_);
  or (_17819_, _17818_, _17816_);
  nor (_17820_, _10945_, _10946_);
  or (_17821_, _17820_, _06648_);
  nor (_17822_, _10662_, _05983_);
  nand (_17823_, _10378_, _07353_);
  nor (_17824_, _08359_, _10010_);
  and (_17825_, _14683_, _08359_);
  or (_17826_, _17825_, _17824_);
  or (_17827_, _17826_, _06044_);
  and (_17828_, _17827_, _06848_);
  and (_17829_, _14672_, _07701_);
  or (_17830_, _17829_, _17817_);
  and (_17831_, _17830_, _06102_);
  or (_17832_, _17219_, _09181_);
  nor (_17833_, _10400_, _07353_);
  nor (_17834_, _06530_, _10010_);
  and (_17835_, _06530_, _10010_);
  or (_17836_, _17835_, _17834_);
  and (_17837_, _17836_, _10400_);
  or (_17838_, _17837_, _10389_);
  or (_17839_, _17838_, _17833_);
  and (_17840_, _17839_, _05698_);
  or (_17841_, _17840_, _06948_);
  and (_17842_, _17841_, _06954_);
  and (_17843_, _17842_, _17832_);
  or (_17844_, _17843_, _17831_);
  and (_17845_, _17844_, _10413_);
  not (_17846_, \oc8051_golden_model_1.PSW [6]);
  nor (_17847_, _10415_, _17846_);
  nor (_17848_, _17847_, \oc8051_golden_model_1.ACC [3]);
  nor (_17849_, _17848_, _10416_);
  and (_17850_, _17849_, _10412_);
  or (_17851_, _17850_, _06043_);
  or (_17852_, _17851_, _17845_);
  and (_17853_, _17852_, _17828_);
  nor (_17854_, _10439_, _07353_);
  or (_17855_, _17854_, _17817_);
  and (_17856_, _17855_, _06239_);
  or (_17857_, _17856_, _10378_);
  or (_17858_, _17857_, _17853_);
  and (_17859_, _17858_, _17823_);
  or (_17860_, _17859_, _06970_);
  or (_17861_, _09181_, _06971_);
  and (_17862_, _17861_, _06220_);
  and (_17863_, _17862_, _17860_);
  nor (_17864_, _08028_, _06220_);
  or (_17865_, _17864_, _10376_);
  or (_17866_, _17865_, _17863_);
  nand (_17867_, _10376_, _08393_);
  and (_17868_, _17867_, _17866_);
  or (_17869_, _17868_, _06039_);
  and (_17870_, _14681_, _08359_);
  or (_17871_, _17870_, _17824_);
  or (_17872_, _17871_, _06040_);
  and (_17873_, _17872_, _06033_);
  and (_17874_, _17873_, _17869_);
  or (_17875_, _17824_, _14708_);
  and (_17876_, _17826_, _06032_);
  and (_17877_, _17876_, _17875_);
  or (_17878_, _17877_, _17874_);
  and (_17879_, _17878_, _09800_);
  or (_17880_, _09750_, _09748_);
  nor (_17881_, _09751_, _09800_);
  and (_17882_, _17881_, _17880_);
  or (_17883_, _17882_, _10468_);
  or (_17884_, _17883_, _17879_);
  and (_17885_, _07530_, \oc8051_golden_model_1.ACC [2]);
  nor (_17886_, _17569_, _17885_);
  nor (_17887_, _10905_, _10906_);
  and (_17888_, _17887_, _17886_);
  nor (_17889_, _17887_, _17886_);
  or (_17890_, _17889_, _17888_);
  nor (_17891_, _17890_, _10606_);
  and (_17892_, _17890_, _10606_);
  nor (_17893_, _17892_, _17891_);
  and (_17894_, _17571_, \oc8051_golden_model_1.PSW [7]);
  nor (_17895_, _17572_, _10606_);
  nor (_17896_, _17895_, _17894_);
  not (_17897_, _17896_);
  and (_17898_, _17897_, _17893_);
  nor (_17899_, _17897_, _17893_);
  nor (_17900_, _17899_, _17898_);
  or (_17901_, _17900_, _10469_);
  and (_17902_, _17901_, _17884_);
  or (_17903_, _17902_, _12361_);
  and (_17904_, _09030_, \oc8051_golden_model_1.ACC [2]);
  nor (_17905_, _17585_, _17904_);
  and (_17906_, _17820_, _17905_);
  nor (_17907_, _17820_, _17905_);
  or (_17908_, _17907_, _17906_);
  or (_17909_, _17908_, _10606_);
  nand (_17910_, _17908_, _10606_);
  and (_17911_, _17910_, _17909_);
  and (_17912_, _17911_, _17591_);
  nor (_17913_, _17911_, _17591_);
  nor (_17914_, _17913_, _17912_);
  or (_17915_, _17914_, _13935_);
  and (_17916_, _17915_, _06267_);
  and (_17917_, _17916_, _17903_);
  and (_17918_, _12305_, \oc8051_golden_model_1.PSW [7]);
  and (_17919_, _08176_, \oc8051_golden_model_1.ACC [2]);
  nor (_17920_, _17603_, _17919_);
  nor (_17921_, _12299_, _17920_);
  and (_17922_, _12299_, _17920_);
  nor (_17923_, _17922_, _17921_);
  and (_17924_, _17609_, _17923_);
  or (_17925_, _17924_, _10306_);
  or (_17926_, _17925_, _17918_);
  and (_17927_, _17926_, _12367_);
  or (_17928_, _17927_, _17917_);
  and (_17929_, _06403_, \oc8051_golden_model_1.ACC [2]);
  nor (_17930_, _17615_, _17929_);
  nor (_17931_, _12319_, _17930_);
  and (_17932_, _12319_, _17930_);
  nor (_17933_, _17932_, _17931_);
  and (_17934_, _17619_, _17933_);
  nor (_17935_, _17619_, _17933_);
  or (_17936_, _17935_, _10307_);
  or (_17937_, _17936_, _17934_);
  and (_17938_, _17937_, _17928_);
  or (_17939_, _17938_, _05676_);
  nand (_17940_, _05983_, _05676_);
  and (_17941_, _17940_, _06027_);
  and (_17942_, _17941_, _17939_);
  and (_17943_, _14724_, _08359_);
  or (_17944_, _17943_, _17824_);
  and (_17945_, _17944_, _06026_);
  or (_17946_, _17945_, _09818_);
  or (_17947_, _17946_, _17942_);
  and (_17948_, _09181_, _07701_);
  or (_17949_, _17817_, _07012_);
  or (_17950_, _17949_, _17948_);
  or (_17951_, _17855_, _09827_);
  and (_17952_, _17951_, _05669_);
  and (_17953_, _17952_, _17950_);
  and (_17954_, _17953_, _17947_);
  and (_17955_, _14778_, _07701_);
  or (_17956_, _17955_, _17817_);
  and (_17957_, _17956_, _09833_);
  or (_17958_, _17957_, _09832_);
  or (_17959_, _17958_, _17954_);
  or (_17960_, _09976_, _09839_);
  and (_17961_, _17960_, _05664_);
  and (_17962_, _17961_, _17959_);
  nor (_17963_, _05983_, _05664_);
  or (_17964_, _17963_, _06019_);
  or (_17965_, _17964_, _17962_);
  and (_17966_, _07701_, _08662_);
  or (_17967_, _17966_, _17817_);
  or (_17968_, _17967_, _06020_);
  and (_17969_, _17968_, _10662_);
  and (_17970_, _17969_, _17965_);
  or (_17971_, _17970_, _17822_);
  and (_17972_, _17971_, _17660_);
  and (_17973_, _17887_, _17656_);
  or (_17974_, _17973_, _17972_);
  and (_17975_, _17974_, _17663_);
  and (_17976_, _17662_, _17887_);
  or (_17977_, _17976_, _17975_);
  and (_17978_, _17977_, _17671_);
  and (_17979_, _17887_, _17666_);
  or (_17980_, _17979_, _17978_);
  and (_17981_, _17980_, _17670_);
  and (_17982_, _17887_, _17503_);
  or (_17983_, _17982_, _17981_);
  and (_17984_, _17983_, _16972_);
  and (_17985_, _16971_, _17887_);
  or (_17986_, _17985_, _06650_);
  or (_17987_, _17986_, _17984_);
  and (_17988_, _10394_, _05726_);
  nor (_17989_, _17887_, _16970_);
  nor (_17990_, _17989_, _17988_);
  and (_17991_, _17990_, _17987_);
  or (_17992_, _17820_, _06647_);
  and (_17993_, _17992_, _10685_);
  or (_17994_, _17993_, _17991_);
  and (_17995_, _17994_, _17821_);
  or (_17996_, _17995_, _06282_);
  or (_17997_, _12299_, _06283_);
  and (_17999_, _17997_, _10699_);
  and (_18000_, _17999_, _17996_);
  and (_18001_, _10698_, _12319_);
  or (_18002_, _18001_, _06112_);
  or (_18003_, _18002_, _18000_);
  nand (_18004_, _18003_, _17819_);
  and (_18005_, _18004_, _08756_);
  nor (_18006_, _17817_, _08756_);
  or (_18007_, _18006_, _11996_);
  or (_18008_, _18007_, _18005_);
  nor (_18009_, _11999_, _11998_);
  nand (_18010_, _11996_, _10905_);
  and (_18011_, _18010_, _18009_);
  and (_18012_, _18011_, _18008_);
  nor (_18013_, _18009_, _10905_);
  or (_18014_, _18013_, _18012_);
  and (_18015_, _18014_, _10736_);
  nor (_18016_, _10736_, _10945_);
  or (_18017_, _18016_, _18015_);
  nand (_18018_, _18017_, _10735_);
  and (_18019_, _18018_, _17815_);
  and (_18020_, _10741_, _11028_);
  or (_18021_, _18020_, _18019_);
  and (_18022_, _18021_, _07032_);
  nand (_18023_, _17967_, _06108_);
  nor (_18024_, _18023_, _10988_);
  or (_18025_, _18024_, _06477_);
  or (_18026_, _18025_, _18022_);
  and (_18027_, _18026_, _17813_);
  or (_18028_, _18027_, _06834_);
  nand (_18029_, _10906_, _06834_);
  and (_18030_, _18029_, _17387_);
  and (_18031_, _18030_, _18028_);
  or (_18032_, _18031_, _17812_);
  nand (_18033_, _10775_, _10946_);
  and (_18034_, _18033_, _06291_);
  and (_18035_, _18034_, _18032_);
  nor (_18036_, _10988_, _06291_);
  or (_18037_, _18036_, _10781_);
  or (_18038_, _18037_, _18035_);
  nand (_18039_, _10781_, _11029_);
  and (_18040_, _18039_, _08777_);
  and (_18041_, _18040_, _18038_);
  and (_18042_, _14792_, _07701_);
  or (_18043_, _18042_, _17817_);
  and (_18044_, _18043_, _06130_);
  or (_18045_, _18044_, _10303_);
  or (_18046_, _18045_, _18041_);
  and (_18047_, _18046_, _17810_);
  or (_18048_, _18047_, _10794_);
  and (_18049_, _10809_, _10528_);
  nor (_18050_, _18049_, _10810_);
  or (_18051_, _18050_, _10796_);
  and (_18052_, _18051_, _06289_);
  and (_18053_, _18052_, _18048_);
  and (_18054_, _10839_, _10341_);
  nor (_18055_, _18054_, _10840_);
  or (_18056_, _18055_, _10824_);
  and (_18057_, _18056_, _10826_);
  or (_18058_, _18057_, _18053_);
  and (_18059_, _10869_, _10598_);
  nor (_18060_, _18059_, _10870_);
  or (_18061_, _18060_, _10856_);
  and (_18062_, _18061_, _10855_);
  and (_18063_, _18062_, _18058_);
  nand (_18064_, _10854_, \oc8051_golden_model_1.ACC [2]);
  nand (_18065_, _18064_, _10889_);
  or (_18066_, _18065_, _18063_);
  nor (_18067_, _10918_, _17887_);
  and (_18068_, _10918_, _17887_);
  or (_18069_, _18068_, _18067_);
  or (_18070_, _18069_, _10889_);
  and (_18071_, _18070_, _10886_);
  and (_18072_, _18071_, _18066_);
  and (_18073_, _18069_, _10885_);
  or (_18074_, _18073_, _10932_);
  or (_18075_, _18074_, _18072_);
  and (_18076_, _10959_, _17820_);
  nor (_18077_, _10959_, _17820_);
  or (_18078_, _18077_, _18076_);
  or (_18079_, _18078_, _10934_);
  and (_18080_, _18079_, _06052_);
  and (_18081_, _18080_, _18075_);
  and (_18082_, _11000_, _12299_);
  nor (_18083_, _11000_, _12299_);
  or (_18084_, _18083_, _18082_);
  and (_18085_, _18084_, _06051_);
  or (_18086_, _18085_, _10974_);
  or (_18087_, _18086_, _18081_);
  and (_18088_, _11040_, _12319_);
  nor (_18089_, _11040_, _12319_);
  or (_18090_, _18089_, _18088_);
  or (_18091_, _18090_, _11050_);
  and (_18092_, _18091_, _11016_);
  and (_18093_, _18092_, _18087_);
  and (_18094_, _11015_, \oc8051_golden_model_1.ACC [2]);
  or (_18095_, _18094_, _06316_);
  or (_18096_, _18095_, _18093_);
  or (_18097_, _17830_, _06718_);
  and (_18098_, _18097_, _11060_);
  and (_18099_, _18098_, _18096_);
  nor (_18100_, _11065_, _10010_);
  or (_18101_, _18100_, _11066_);
  and (_18102_, _18101_, _11059_);
  or (_18103_, _18102_, _11064_);
  or (_18104_, _18103_, _18099_);
  nand (_18105_, _11064_, _09880_);
  and (_18106_, _18105_, _05653_);
  and (_18107_, _18106_, _18104_);
  and (_18108_, _17871_, _05652_);
  or (_18109_, _18108_, _06047_);
  or (_18110_, _18109_, _18107_);
  and (_18111_, _14849_, _07701_);
  or (_18112_, _17817_, _06048_);
  or (_18113_, _18112_, _18111_);
  and (_18114_, _18113_, _11083_);
  and (_18115_, _18114_, _18110_);
  nor (_18116_, _11091_, \oc8051_golden_model_1.ACC [3]);
  nor (_18117_, _18116_, _11092_);
  and (_18118_, _18117_, _11082_);
  or (_18119_, _18118_, _11089_);
  or (_18120_, _18119_, _18115_);
  nand (_18121_, _11089_, _09880_);
  and (_18122_, _18121_, _01336_);
  and (_18123_, _18122_, _18120_);
  or (_18124_, _18123_, _17807_);
  and (_43335_, _18124_, _42882_);
  nor (_18125_, _01336_, _09880_);
  not (_18126_, _17437_);
  or (_18127_, _10961_, _10944_);
  and (_18128_, _18127_, _10962_);
  or (_18129_, _18128_, _18126_);
  and (_18130_, _14876_, _07701_);
  nor (_18131_, _07701_, _09880_);
  or (_18132_, _18131_, _08751_);
  or (_18133_, _18132_, _18130_);
  or (_18134_, _10686_, _10944_);
  and (_18135_, _06095_, _05661_);
  and (_18136_, _18135_, _05726_);
  not (_18137_, _17909_);
  or (_18138_, _17912_, _18137_);
  and (_18139_, _09181_, _10010_);
  or (_18140_, _09181_, _10010_);
  and (_18141_, _18140_, _17905_);
  or (_18142_, _18141_, _18139_);
  nor (_18143_, _10944_, _18142_);
  and (_18144_, _10944_, _18142_);
  or (_18145_, _18144_, _18143_);
  or (_18146_, _18145_, _10606_);
  nand (_18147_, _18145_, _10606_);
  and (_18148_, _18147_, _18146_);
  and (_18149_, _18148_, _18138_);
  nor (_18150_, _18148_, _18138_);
  nor (_18151_, _18150_, _18149_);
  or (_18152_, _18151_, _13935_);
  nand (_18153_, _10378_, _08270_);
  nor (_18154_, _08359_, _09880_);
  and (_18155_, _14878_, _08359_);
  or (_18156_, _18155_, _18154_);
  or (_18157_, _18156_, _06044_);
  and (_18158_, _18157_, _06848_);
  and (_18159_, _14887_, _07701_);
  or (_18160_, _18159_, _18131_);
  and (_18161_, _18160_, _06102_);
  or (_18162_, _10390_, _09180_);
  nor (_18163_, _10400_, _08270_);
  or (_18164_, _06530_, \oc8051_golden_model_1.ACC [4]);
  nand (_18165_, _06530_, \oc8051_golden_model_1.ACC [4]);
  and (_18166_, _18165_, _18164_);
  and (_18167_, _18166_, _10400_);
  or (_18168_, _18167_, _10389_);
  or (_18169_, _18168_, _18163_);
  and (_18170_, _18169_, _10408_);
  and (_18171_, _18170_, _18162_);
  or (_18172_, _18171_, _18161_);
  and (_18173_, _18172_, _10413_);
  nor (_18174_, _10416_, \oc8051_golden_model_1.ACC [4]);
  nor (_18175_, _18174_, _10417_);
  and (_18176_, _18175_, _10412_);
  or (_18177_, _18176_, _06043_);
  or (_18178_, _18177_, _18173_);
  and (_18179_, _18178_, _18158_);
  nor (_18180_, _08270_, _10439_);
  or (_18181_, _18180_, _18131_);
  and (_18182_, _18181_, _06239_);
  or (_18183_, _18182_, _10378_);
  or (_18184_, _18183_, _18179_);
  and (_18185_, _18184_, _18153_);
  or (_18186_, _18185_, _06970_);
  or (_18187_, _09180_, _06971_);
  and (_18189_, _18187_, _06220_);
  and (_18190_, _18189_, _18186_);
  nor (_18191_, _08272_, _06220_);
  or (_18192_, _18191_, _10376_);
  or (_18193_, _18192_, _18190_);
  nand (_18194_, _10376_, _05758_);
  and (_18195_, _18194_, _18193_);
  or (_18196_, _18195_, _06039_);
  and (_18197_, _14882_, _08359_);
  or (_18198_, _18197_, _18154_);
  or (_18200_, _18198_, _06040_);
  and (_18201_, _18200_, _06033_);
  and (_18202_, _18201_, _18196_);
  or (_18203_, _18154_, _14914_);
  and (_18204_, _18156_, _06032_);
  and (_18205_, _18204_, _18203_);
  or (_18206_, _18205_, _09269_);
  or (_18207_, _18206_, _18202_);
  nor (_18208_, _09753_, _09751_);
  nor (_18209_, _18208_, _09754_);
  or (_18211_, _18209_, _09800_);
  and (_18212_, _18211_, _10469_);
  and (_18213_, _18212_, _18207_);
  or (_18214_, _17898_, _17891_);
  nor (_18215_, _07353_, \oc8051_golden_model_1.ACC [3]);
  nand (_18216_, _07353_, \oc8051_golden_model_1.ACC [3]);
  and (_18217_, _18216_, _17886_);
  or (_18218_, _18217_, _18215_);
  nor (_18219_, _10904_, _18218_);
  and (_18220_, _10904_, _18218_);
  nor (_18222_, _18220_, _18219_);
  and (_18223_, _18222_, \oc8051_golden_model_1.PSW [7]);
  nor (_18224_, _18222_, \oc8051_golden_model_1.PSW [7]);
  nor (_18225_, _18224_, _18223_);
  or (_18226_, _18225_, _18214_);
  and (_18227_, _18225_, _18214_);
  nor (_18228_, _18227_, _10469_);
  and (_18229_, _18228_, _18226_);
  or (_18230_, _18229_, _12361_);
  or (_18231_, _18230_, _18213_);
  and (_18233_, _18231_, _18152_);
  or (_18234_, _18233_, _06261_);
  nor (_18235_, _12305_, _10606_);
  or (_18236_, _17920_, _13781_);
  and (_18237_, _18236_, _13780_);
  nor (_18238_, _10986_, _18237_);
  and (_18239_, _10986_, _18237_);
  nor (_18240_, _18239_, _18238_);
  and (_18241_, _18240_, \oc8051_golden_model_1.PSW [7]);
  nor (_18242_, _18240_, \oc8051_golden_model_1.PSW [7]);
  nor (_18244_, _18242_, _18241_);
  and (_18245_, _18244_, _18235_);
  nor (_18246_, _18244_, _18235_);
  nor (_18247_, _18246_, _18245_);
  or (_18248_, _18247_, _06267_);
  and (_18249_, _18248_, _10307_);
  and (_18250_, _18249_, _18234_);
  nor (_18251_, _12324_, _10606_);
  or (_18252_, _17930_, _13880_);
  and (_18253_, _18252_, _13879_);
  nor (_18255_, _11027_, _18253_);
  and (_18256_, _11027_, _18253_);
  nor (_18257_, _18256_, _18255_);
  and (_18258_, _18257_, \oc8051_golden_model_1.PSW [7]);
  nor (_18259_, _18257_, \oc8051_golden_model_1.PSW [7]);
  nor (_18260_, _18259_, _18258_);
  or (_18261_, _18260_, _18251_);
  and (_18262_, _18260_, _18251_);
  nor (_18263_, _18262_, _10307_);
  and (_18264_, _18263_, _18261_);
  or (_18266_, _18264_, _05676_);
  or (_18267_, _18266_, _18250_);
  nand (_18268_, _06758_, _05676_);
  and (_18269_, _18268_, _06027_);
  and (_18270_, _18269_, _18267_);
  or (_18271_, _18154_, _14879_);
  and (_18272_, _18271_, _06026_);
  and (_18273_, _18272_, _18156_);
  or (_18274_, _18273_, _09818_);
  or (_18275_, _18274_, _18270_);
  and (_18277_, _09180_, _07701_);
  or (_18278_, _18131_, _07012_);
  or (_18279_, _18278_, _18277_);
  or (_18280_, _18181_, _09827_);
  and (_18281_, _18280_, _05669_);
  and (_18282_, _18281_, _18279_);
  and (_18283_, _18282_, _18275_);
  and (_18284_, _14983_, _07701_);
  or (_18285_, _18284_, _18131_);
  and (_18286_, _18285_, _09833_);
  or (_18288_, _18286_, _09832_);
  or (_18289_, _18288_, _18283_);
  or (_18290_, _09924_, _09839_);
  and (_18291_, _18290_, _05664_);
  and (_18292_, _18291_, _18289_);
  nor (_18293_, _06758_, _05664_);
  or (_18294_, _18293_, _06019_);
  or (_18295_, _18294_, _18292_);
  and (_18296_, _08665_, _07701_);
  or (_18297_, _18296_, _18131_);
  or (_18299_, _18297_, _06020_);
  and (_18300_, _18299_, _10662_);
  and (_18301_, _18300_, _18295_);
  nor (_18302_, _10662_, _06758_);
  or (_18303_, _18302_, _17656_);
  or (_18304_, _18303_, _18301_);
  not (_18305_, _06649_);
  or (_18306_, _10904_, _17660_);
  and (_18307_, _18306_, _18305_);
  and (_18308_, _18307_, _18304_);
  and (_18310_, _06098_, _05726_);
  and (_18311_, _10904_, _06649_);
  or (_18312_, _18311_, _18310_);
  or (_18313_, _18312_, _18308_);
  and (_18314_, _06136_, _05726_);
  not (_18315_, _18314_);
  not (_18316_, _18310_);
  or (_18317_, _10904_, _18316_);
  and (_18318_, _18317_, _18315_);
  and (_18319_, _18318_, _18313_);
  and (_18321_, _10904_, _18314_);
  or (_18322_, _18321_, _17666_);
  or (_18323_, _18322_, _18319_);
  or (_18324_, _10904_, _17671_);
  nand (_18325_, _18324_, _18323_);
  nor (_18326_, _18325_, _18136_);
  and (_18327_, _18136_, _10904_);
  or (_18328_, _18327_, _10685_);
  or (_18329_, _18328_, _18326_);
  and (_18330_, _18329_, _18134_);
  or (_18332_, _18330_, _06282_);
  or (_18333_, _10986_, _06283_);
  and (_18334_, _18333_, _10699_);
  and (_18335_, _18334_, _18332_);
  nor (_18336_, _10699_, _11026_);
  or (_18337_, _18336_, _06112_);
  or (_18338_, _18337_, _18335_);
  nand (_18339_, _18338_, _18133_);
  and (_18340_, _18339_, _08756_);
  nor (_18341_, _18131_, _08756_);
  or (_18343_, _18341_, _11996_);
  or (_18344_, _18343_, _18340_);
  and (_18345_, _18135_, _05735_);
  or (_18346_, _18345_, _10901_);
  nand (_18347_, _18346_, _17104_);
  and (_18348_, _18347_, _18344_);
  and (_18349_, _18345_, _10903_);
  or (_18350_, _18349_, _10731_);
  nor (_18351_, _18350_, _18348_);
  nor (_18352_, _10736_, _10942_);
  or (_18354_, _18352_, _06279_);
  or (_18355_, _18354_, _18351_);
  or (_18356_, _10983_, _10735_);
  and (_18357_, _18356_, _10747_);
  and (_18358_, _18357_, _18355_);
  and (_18359_, _10741_, _11023_);
  or (_18360_, _18359_, _18358_);
  and (_18361_, _18360_, _07032_);
  nand (_18362_, _18297_, _06108_);
  nor (_18363_, _18362_, _10985_);
  or (_18364_, _18363_, _10752_);
  or (_18365_, _18364_, _18361_);
  or (_18366_, _10902_, _17205_);
  and (_18367_, _18366_, _10760_);
  and (_18368_, _18367_, _18365_);
  and (_18369_, _10759_, _10902_);
  or (_18370_, _18369_, _10767_);
  or (_18371_, _18370_, _18368_);
  or (_18372_, _10766_, _10902_);
  and (_18373_, _18372_, _06668_);
  and (_18375_, _18373_, _18371_);
  and (_18376_, _10902_, _06667_);
  or (_18377_, _18376_, _10775_);
  or (_18378_, _18377_, _18375_);
  or (_18379_, _17395_, _10943_);
  and (_18380_, _18379_, _06291_);
  and (_18381_, _18380_, _18378_);
  nor (_18382_, _10985_, _06291_);
  or (_18383_, _18382_, _10781_);
  or (_18384_, _18383_, _18381_);
  nand (_18386_, _10781_, _11025_);
  and (_18387_, _18386_, _18384_);
  or (_18388_, _18387_, _06130_);
  and (_18389_, _14873_, _07701_);
  or (_18390_, _18131_, _08777_);
  or (_18391_, _18390_, _18389_);
  and (_18392_, _18391_, _10304_);
  and (_18393_, _18392_, _18388_);
  or (_18394_, _10293_, _10265_);
  and (_18395_, _10303_, _10294_);
  and (_18397_, _18395_, _18394_);
  or (_18398_, _18397_, _17409_);
  or (_18399_, _18398_, _18393_);
  or (_18400_, _10811_, _10521_);
  and (_18401_, _18400_, _10812_);
  or (_18402_, _18401_, _17410_);
  and (_18403_, _18402_, _17423_);
  and (_18404_, _18403_, _18399_);
  and (_18405_, _18401_, _17416_);
  or (_18406_, _18405_, _06288_);
  or (_18408_, _18406_, _18404_);
  or (_18409_, _10841_, _10335_);
  and (_18410_, _18409_, _10842_);
  or (_18411_, _18410_, _06289_);
  and (_18412_, _18411_, _10856_);
  and (_18413_, _18412_, _18408_);
  or (_18414_, _10871_, _10592_);
  and (_18415_, _18414_, _10872_);
  and (_18416_, _18415_, _10824_);
  or (_18417_, _18416_, _10854_);
  or (_18419_, _18417_, _18413_);
  nand (_18420_, _10854_, _10010_);
  and (_18421_, _18420_, _10890_);
  and (_18422_, _18421_, _18419_);
  or (_18423_, _10920_, _10904_);
  nor (_18424_, _10921_, _10890_);
  and (_18425_, _18424_, _18423_);
  or (_18426_, _18425_, _17437_);
  or (_18427_, _18426_, _18422_);
  and (_18428_, _18427_, _18129_);
  or (_18430_, _18428_, _06692_);
  or (_18431_, _18128_, _17443_);
  and (_18432_, _18431_, _10975_);
  and (_18433_, _18432_, _18430_);
  or (_18434_, _11002_, _10986_);
  and (_18435_, _11003_, _06051_);
  and (_18436_, _18435_, _18434_);
  or (_18437_, _11042_, _11027_);
  and (_18438_, _11043_, _10974_);
  and (_18439_, _18438_, _18437_);
  or (_18441_, _18439_, _11015_);
  or (_18442_, _18441_, _18436_);
  or (_18443_, _18442_, _18433_);
  nand (_18444_, _11015_, _10010_);
  and (_18445_, _18444_, _18443_);
  or (_18446_, _18445_, _06316_);
  or (_18447_, _18160_, _06718_);
  and (_18448_, _18447_, _11060_);
  and (_18449_, _18448_, _18446_);
  nor (_18450_, _11066_, _09880_);
  or (_18452_, _18450_, _11067_);
  and (_18453_, _18452_, _11059_);
  or (_18454_, _18453_, _11064_);
  or (_18455_, _18454_, _18449_);
  nand (_18456_, _11064_, _09906_);
  and (_18457_, _18456_, _05653_);
  and (_18458_, _18457_, _18455_);
  and (_18459_, _18198_, _05652_);
  or (_18460_, _18459_, _06047_);
  or (_18461_, _18460_, _18458_);
  and (_18463_, _15055_, _07701_);
  or (_18464_, _18131_, _06048_);
  or (_18465_, _18464_, _18463_);
  and (_18466_, _18465_, _11083_);
  and (_18467_, _18466_, _18461_);
  nor (_18468_, _11092_, \oc8051_golden_model_1.ACC [4]);
  nor (_18469_, _18468_, _11093_);
  and (_18470_, _18469_, _11082_);
  or (_18471_, _18470_, _11089_);
  or (_18472_, _18471_, _18467_);
  nand (_18474_, _11089_, _09906_);
  and (_18475_, _18474_, _01336_);
  and (_18476_, _18475_, _18472_);
  or (_18477_, _18476_, _18125_);
  and (_43336_, _18477_, _42882_);
  nor (_18478_, _01336_, _09906_);
  and (_18479_, _10295_, _10259_);
  nor (_18480_, _18479_, _10296_);
  or (_18481_, _18480_, _10304_);
  and (_18482_, _15195_, _07701_);
  nor (_18484_, _07701_, _09906_);
  or (_18485_, _18484_, _08751_);
  or (_18486_, _18485_, _18482_);
  and (_18487_, _10677_, _10899_);
  and (_18488_, _08937_, \oc8051_golden_model_1.ACC [4]);
  nor (_18489_, _18143_, _18488_);
  or (_18490_, _10941_, _18489_);
  nand (_18491_, _10941_, _18489_);
  and (_18492_, _18491_, _18490_);
  or (_18493_, _18492_, _10606_);
  nand (_18495_, _18492_, _10606_);
  and (_18496_, _18495_, _18493_);
  not (_18497_, _18146_);
  or (_18498_, _18149_, _18497_);
  nand (_18499_, _18498_, _18496_);
  or (_18500_, _18498_, _18496_);
  and (_18501_, _18500_, _18499_);
  or (_18502_, _18501_, _13935_);
  nand (_18503_, _10378_, _07977_);
  or (_18504_, _10390_, _09179_);
  nor (_18506_, _10400_, _07977_);
  or (_18507_, _06530_, \oc8051_golden_model_1.ACC [5]);
  nand (_18508_, _06530_, \oc8051_golden_model_1.ACC [5]);
  and (_18509_, _18508_, _18507_);
  and (_18510_, _18509_, _10400_);
  or (_18511_, _18510_, _10389_);
  or (_18512_, _18511_, _18506_);
  and (_18513_, _18512_, _10408_);
  and (_18514_, _18513_, _18504_);
  and (_18515_, _15093_, _07701_);
  or (_18517_, _18515_, _18484_);
  and (_18518_, _18517_, _06102_);
  or (_18519_, _18518_, _10412_);
  or (_18520_, _18519_, _18514_);
  nor (_18521_, _10431_, _10424_);
  nand (_18522_, _10431_, _10424_);
  nand (_18523_, _18522_, _10412_);
  or (_18524_, _18523_, _18521_);
  and (_18525_, _18524_, _06244_);
  and (_18526_, _18525_, _18520_);
  nor (_18528_, _08359_, _09906_);
  and (_18529_, _15073_, _08359_);
  or (_18530_, _18529_, _18528_);
  and (_18531_, _18530_, _06043_);
  nor (_18532_, _07977_, _10439_);
  or (_18533_, _18532_, _18484_);
  and (_18534_, _18533_, _06239_);
  or (_18535_, _18534_, _10378_);
  or (_18536_, _18535_, _18531_);
  or (_18537_, _18536_, _18526_);
  and (_18539_, _18537_, _18503_);
  or (_18540_, _18539_, _06970_);
  or (_18541_, _09179_, _06971_);
  and (_18542_, _18541_, _06220_);
  and (_18543_, _18542_, _18540_);
  nor (_18544_, _07979_, _06220_);
  or (_18545_, _18544_, _10376_);
  or (_18546_, _18545_, _18543_);
  nand (_18547_, _10376_, _05784_);
  and (_18548_, _18547_, _18546_);
  or (_18550_, _18548_, _06039_);
  and (_18551_, _15077_, _08359_);
  or (_18552_, _18551_, _18528_);
  or (_18553_, _18552_, _06040_);
  and (_18554_, _18553_, _06033_);
  and (_18555_, _18554_, _18550_);
  or (_18556_, _18528_, _15110_);
  and (_18557_, _18530_, _06032_);
  and (_18558_, _18557_, _18556_);
  or (_18559_, _18558_, _18555_);
  and (_18561_, _18559_, _09800_);
  or (_18562_, _09756_, _09754_);
  nor (_18563_, _09757_, _09800_);
  and (_18564_, _18563_, _18562_);
  or (_18565_, _18564_, _10468_);
  or (_18566_, _18565_, _18561_);
  and (_18567_, _08270_, \oc8051_golden_model_1.ACC [4]);
  nor (_18568_, _18219_, _18567_);
  and (_18569_, _10900_, _18568_);
  nor (_18570_, _10900_, _18568_);
  nor (_18572_, _18570_, _18569_);
  nor (_18573_, _18572_, _10606_);
  and (_18574_, _18572_, _10606_);
  nor (_18575_, _18574_, _18573_);
  nor (_18576_, _18227_, _18223_);
  not (_18577_, _18576_);
  and (_18578_, _18577_, _18575_);
  nor (_18579_, _18577_, _18575_);
  nor (_18580_, _18579_, _18578_);
  or (_18581_, _18580_, _10469_);
  and (_18583_, _18581_, _18566_);
  or (_18584_, _18583_, _12361_);
  and (_18585_, _18584_, _06267_);
  and (_18586_, _18585_, _18502_);
  and (_18587_, _08272_, \oc8051_golden_model_1.ACC [4]);
  nor (_18588_, _18238_, _18587_);
  nor (_18589_, _12306_, _18588_);
  and (_18590_, _12306_, _18588_);
  nor (_18591_, _18590_, _18589_);
  and (_18592_, _18591_, \oc8051_golden_model_1.PSW [7]);
  nor (_18594_, _18591_, \oc8051_golden_model_1.PSW [7]);
  nor (_18595_, _18594_, _18592_);
  nor (_18596_, _18245_, _18241_);
  not (_18597_, _18596_);
  or (_18598_, _18597_, _18595_);
  and (_18599_, _18597_, _18595_);
  nor (_18600_, _18599_, _06267_);
  and (_18601_, _18600_, _18598_);
  or (_18602_, _18601_, _18586_);
  and (_18603_, _18602_, _10307_);
  and (_18605_, _06758_, \oc8051_golden_model_1.ACC [4]);
  nor (_18606_, _18255_, _18605_);
  nor (_18607_, _12325_, _18606_);
  and (_18608_, _12325_, _18606_);
  nor (_18609_, _18608_, _18607_);
  and (_18610_, _18609_, \oc8051_golden_model_1.PSW [7]);
  nor (_18611_, _18609_, \oc8051_golden_model_1.PSW [7]);
  nor (_18612_, _18611_, _18610_);
  nor (_18613_, _18262_, _18258_);
  not (_18614_, _18613_);
  or (_18616_, _18614_, _18612_);
  and (_18617_, _18614_, _18612_);
  nor (_18618_, _18617_, _10307_);
  and (_18619_, _18618_, _18616_);
  or (_18620_, _18619_, _05676_);
  or (_18621_, _18620_, _18603_);
  nand (_18622_, _06359_, _05676_);
  and (_18623_, _18622_, _06027_);
  and (_18624_, _18623_, _18621_);
  or (_18625_, _18528_, _15074_);
  and (_18627_, _18625_, _06026_);
  and (_18628_, _18627_, _18530_);
  or (_18629_, _18628_, _09818_);
  or (_18630_, _18629_, _18624_);
  and (_18631_, _09179_, _07701_);
  or (_18632_, _18484_, _07012_);
  or (_18633_, _18632_, _18631_);
  or (_18634_, _18533_, _09827_);
  and (_18635_, _18634_, _05669_);
  and (_18636_, _18635_, _18633_);
  and (_18638_, _18636_, _18630_);
  and (_18639_, _15179_, _07701_);
  or (_18640_, _18639_, _18484_);
  and (_18641_, _18640_, _09833_);
  or (_18642_, _18641_, _09832_);
  or (_18643_, _18642_, _18638_);
  or (_18644_, _09894_, _09839_);
  and (_18645_, _18644_, _05664_);
  and (_18646_, _18645_, _18643_);
  nor (_18647_, _06359_, _05664_);
  or (_18649_, _18647_, _06019_);
  or (_18650_, _18649_, _18646_);
  and (_18651_, _08652_, _07701_);
  or (_18652_, _18651_, _18484_);
  or (_18653_, _18652_, _06020_);
  and (_18654_, _18653_, _10662_);
  and (_18655_, _18654_, _18650_);
  nor (_18656_, _10662_, _06359_);
  or (_18657_, _18656_, _17656_);
  or (_18658_, _18657_, _18655_);
  or (_18659_, _10899_, _17660_);
  and (_18660_, _18659_, _18658_);
  and (_18661_, _18660_, _18305_);
  and (_18662_, _10899_, _06649_);
  or (_18663_, _18662_, _18310_);
  or (_18664_, _18663_, _18661_);
  or (_18665_, _10899_, _18316_);
  and (_18666_, _18665_, _10678_);
  and (_18667_, _18666_, _18664_);
  or (_18668_, _18667_, _18487_);
  and (_18671_, _18668_, _16972_);
  and (_18672_, _16971_, _10899_);
  or (_18673_, _18672_, _18671_);
  and (_18674_, _18673_, _16970_);
  and (_18675_, _10899_, _06650_);
  or (_18676_, _18675_, _18674_);
  and (_18677_, _18676_, _10686_);
  nor (_18678_, _10686_, _10941_);
  or (_18679_, _18678_, _06282_);
  or (_18680_, _18679_, _18677_);
  or (_18682_, _12306_, _06283_);
  and (_18683_, _18682_, _10699_);
  and (_18684_, _18683_, _18680_);
  and (_18685_, _10698_, _12325_);
  or (_18686_, _18685_, _06112_);
  or (_18687_, _18686_, _18684_);
  and (_18688_, _18687_, _18486_);
  or (_18689_, _18688_, _06284_);
  or (_18690_, _18484_, _08756_);
  and (_18691_, _18690_, _11997_);
  and (_18692_, _18691_, _18689_);
  or (_18693_, _18345_, _10897_);
  and (_18694_, _18693_, _17104_);
  or (_18695_, _18694_, _18692_);
  or (_18696_, _18009_, _10897_);
  and (_18697_, _18696_, _18695_);
  or (_18698_, _18697_, _10731_);
  or (_18699_, _10736_, _10939_);
  and (_18700_, _18699_, _10735_);
  and (_18701_, _18700_, _18698_);
  or (_18704_, _10741_, _10981_);
  and (_18705_, _18704_, _10743_);
  or (_18706_, _18705_, _18701_);
  or (_18707_, _10747_, _11021_);
  and (_18708_, _18707_, _07032_);
  and (_18709_, _18708_, _18706_);
  nand (_18710_, _18652_, _06108_);
  nor (_18711_, _18710_, _10982_);
  or (_18712_, _18711_, _10752_);
  or (_18713_, _18712_, _18709_);
  and (_18715_, _10898_, _10752_);
  nor (_18716_, _18715_, _17203_);
  and (_18717_, _18716_, _18713_);
  not (_18718_, _10898_);
  nand (_18719_, _18718_, _17203_);
  nor (_18720_, _10765_, _06834_);
  nand (_18721_, _18720_, _18719_);
  or (_18722_, _18721_, _18717_);
  or (_18723_, _18720_, _18718_);
  and (_18724_, _18723_, _06668_);
  and (_18725_, _18724_, _18722_);
  nor (_18726_, _10898_, _06668_);
  or (_18727_, _18726_, _10775_);
  or (_18728_, _18727_, _18725_);
  nand (_18729_, _10775_, _09906_);
  or (_18730_, _18729_, _09179_);
  and (_18731_, _18730_, _06291_);
  and (_18732_, _18731_, _18728_);
  nand (_18733_, _17136_, _10982_);
  and (_18734_, _18733_, _11987_);
  or (_18737_, _18734_, _18732_);
  nand (_18738_, _10781_, _11022_);
  and (_18739_, _18738_, _08777_);
  and (_18740_, _18739_, _18737_);
  and (_18741_, _15194_, _07701_);
  or (_18742_, _18741_, _18484_);
  and (_18743_, _18742_, _06130_);
  or (_18744_, _18743_, _10303_);
  or (_18745_, _18744_, _18740_);
  and (_18746_, _18745_, _18481_);
  or (_18748_, _18746_, _10794_);
  and (_18749_, _10813_, _10518_);
  nor (_18750_, _18749_, _10814_);
  or (_18751_, _18750_, _10796_);
  and (_18752_, _18751_, _06289_);
  and (_18753_, _18752_, _18748_);
  and (_18754_, _10843_, _10329_);
  nor (_18755_, _18754_, _10844_);
  or (_18756_, _18755_, _10824_);
  and (_18757_, _18756_, _10826_);
  or (_18758_, _18757_, _18753_);
  and (_18759_, _10873_, _10589_);
  nor (_18760_, _18759_, _10874_);
  or (_18761_, _18760_, _10856_);
  and (_18762_, _18761_, _10855_);
  and (_18763_, _18762_, _18758_);
  and (_18764_, _10854_, \oc8051_golden_model_1.ACC [4]);
  or (_18765_, _18764_, _10887_);
  or (_18766_, _18765_, _18763_);
  nor (_18767_, _10885_, _06691_);
  not (_18770_, _18767_);
  nor (_18771_, _06136_, _06229_);
  nor (_18772_, _18771_, _06841_);
  or (_18773_, _18772_, _18770_);
  not (_18774_, _18773_);
  and (_18775_, _10922_, _10900_);
  nor (_18776_, _18775_, _10923_);
  and (_18777_, _18776_, _18774_);
  or (_18778_, _18777_, _10890_);
  and (_18779_, _18778_, _18766_);
  and (_18781_, _18776_, _18773_);
  or (_18782_, _18781_, _10932_);
  or (_18783_, _18782_, _18779_);
  and (_18784_, _10963_, _10941_);
  nor (_18785_, _18784_, _10964_);
  or (_18786_, _18785_, _10934_);
  and (_18787_, _18786_, _06052_);
  and (_18788_, _18787_, _18783_);
  and (_18789_, _11004_, _12306_);
  nor (_18790_, _11004_, _12306_);
  or (_18791_, _18790_, _18789_);
  and (_18792_, _18791_, _06051_);
  or (_18793_, _18792_, _10974_);
  or (_18794_, _18793_, _18788_);
  and (_18795_, _11044_, _12325_);
  nor (_18796_, _11044_, _12325_);
  or (_18797_, _18796_, _11050_);
  or (_18798_, _18797_, _18795_);
  and (_18799_, _18798_, _11016_);
  and (_18800_, _18799_, _18794_);
  and (_18803_, _11015_, \oc8051_golden_model_1.ACC [4]);
  or (_18804_, _18803_, _06316_);
  or (_18805_, _18804_, _18800_);
  or (_18806_, _18517_, _06718_);
  and (_18807_, _18806_, _11060_);
  and (_18808_, _18807_, _18805_);
  nor (_18809_, _11067_, _09906_);
  or (_18810_, _18809_, _11068_);
  nor (_18811_, _18810_, _11064_);
  nor (_18812_, _18811_, _12756_);
  or (_18814_, _18812_, _18808_);
  nand (_18815_, _11064_, _09861_);
  and (_18816_, _18815_, _05653_);
  and (_18817_, _18816_, _18814_);
  and (_18818_, _18552_, _05652_);
  or (_18819_, _18818_, _06047_);
  or (_18820_, _18819_, _18817_);
  and (_18821_, _15253_, _07701_);
  or (_18822_, _18484_, _06048_);
  or (_18823_, _18822_, _18821_);
  and (_18824_, _18823_, _11083_);
  and (_18825_, _18824_, _18820_);
  nor (_18826_, _11093_, \oc8051_golden_model_1.ACC [5]);
  nor (_18827_, _18826_, _11094_);
  and (_18828_, _18827_, _11082_);
  or (_18829_, _18828_, _11089_);
  or (_18830_, _18829_, _18825_);
  nand (_18831_, _11089_, _09861_);
  and (_18832_, _18831_, _01336_);
  and (_18833_, _18832_, _18830_);
  or (_18836_, _18833_, _18478_);
  and (_43338_, _18836_, _42882_);
  nor (_18837_, _01336_, _09861_);
  nand (_18838_, _11015_, _09906_);
  or (_18839_, _11006_, _10980_);
  and (_18840_, _18839_, _11007_);
  or (_18841_, _18840_, _06052_);
  and (_18842_, _18841_, _11050_);
  nor (_18843_, _10845_, _10368_);
  nor (_18844_, _18843_, _10846_);
  or (_18846_, _18844_, _06289_);
  and (_18847_, _18846_, _10856_);
  or (_18848_, _10893_, _10722_);
  and (_18849_, _15399_, _07701_);
  nor (_18850_, _07701_, _09861_);
  or (_18851_, _18850_, _08751_);
  or (_18852_, _18851_, _18849_);
  and (_18853_, _10669_, _10896_);
  and (_18854_, _15382_, _07701_);
  or (_18855_, _18854_, _18850_);
  and (_18856_, _18855_, _09833_);
  or (_18857_, _09179_, _09906_);
  and (_18858_, _09179_, _09906_);
  or (_18859_, _18489_, _18858_);
  and (_18860_, _18859_, _18857_);
  nor (_18861_, _18860_, _10938_);
  and (_18862_, _18860_, _10938_);
  nor (_18863_, _18862_, _18861_);
  and (_18864_, _18499_, _18493_);
  and (_18865_, _18864_, \oc8051_golden_model_1.PSW [7]);
  or (_18868_, _18865_, _18863_);
  nand (_18869_, _18865_, _18863_);
  and (_18870_, _18869_, _12361_);
  and (_18871_, _18870_, _18868_);
  nand (_18872_, _10378_, _07883_);
  or (_18873_, _10390_, _09178_);
  nor (_18874_, _10400_, _07883_);
  nor (_18875_, _06530_, _09861_);
  and (_18876_, _06530_, _09861_);
  or (_18877_, _18876_, _18875_);
  and (_18879_, _18877_, _10400_);
  or (_18880_, _18879_, _10389_);
  or (_18881_, _18880_, _18874_);
  and (_18882_, _18881_, _10408_);
  and (_18883_, _18882_, _18873_);
  and (_18884_, _15293_, _07701_);
  or (_18885_, _18884_, _18850_);
  and (_18886_, _18885_, _06102_);
  or (_18887_, _18886_, _10412_);
  or (_18888_, _18887_, _18883_);
  not (_18890_, _10426_);
  and (_18891_, _18521_, _18890_);
  or (_18892_, _18521_, _18890_);
  nand (_18893_, _18892_, _10412_);
  or (_18894_, _18893_, _18891_);
  and (_18895_, _18894_, _06244_);
  and (_18896_, _18895_, _18888_);
  nor (_18897_, _08359_, _09861_);
  and (_18898_, _15280_, _08359_);
  or (_18899_, _18898_, _18897_);
  and (_18901_, _18899_, _06043_);
  nor (_18902_, _07883_, _10439_);
  or (_18903_, _18902_, _18850_);
  and (_18904_, _18903_, _06239_);
  or (_18905_, _18904_, _10378_);
  or (_18906_, _18905_, _18901_);
  or (_18907_, _18906_, _18896_);
  and (_18908_, _18907_, _18872_);
  or (_18909_, _18908_, _06970_);
  or (_18910_, _09178_, _06971_);
  and (_18912_, _18910_, _06220_);
  and (_18913_, _18912_, _18909_);
  nor (_18914_, _07885_, _06220_);
  or (_18915_, _18914_, _10376_);
  or (_18916_, _18915_, _18913_);
  nand (_18917_, _10376_, _09956_);
  and (_18918_, _18917_, _18916_);
  or (_18919_, _18918_, _06039_);
  and (_18920_, _15278_, _08359_);
  or (_18921_, _18920_, _18897_);
  or (_18923_, _18921_, _06040_);
  and (_18924_, _18923_, _06033_);
  and (_18925_, _18924_, _18919_);
  or (_18926_, _18897_, _15310_);
  and (_18927_, _18899_, _06032_);
  and (_18928_, _18927_, _18926_);
  or (_18929_, _18928_, _09269_);
  or (_18930_, _18929_, _18925_);
  nor (_18931_, _09759_, _09757_);
  nor (_18932_, _18931_, _09760_);
  or (_18934_, _18932_, _09800_);
  and (_18935_, _18934_, _10469_);
  and (_18936_, _18935_, _18930_);
  nand (_18937_, _07977_, \oc8051_golden_model_1.ACC [5]);
  nor (_18938_, _07977_, \oc8051_golden_model_1.ACC [5]);
  or (_18939_, _18568_, _18938_);
  and (_18940_, _18939_, _18937_);
  nor (_18941_, _18940_, _10896_);
  and (_18942_, _18940_, _10896_);
  nor (_18943_, _18942_, _18941_);
  nor (_18945_, _18578_, _18573_);
  and (_18946_, _18945_, \oc8051_golden_model_1.PSW [7]);
  nand (_18947_, _18946_, _18943_);
  or (_18948_, _18946_, _18943_);
  and (_18949_, _18948_, _10468_);
  and (_18950_, _18949_, _18947_);
  or (_18951_, _18950_, _18936_);
  and (_18952_, _18951_, _13935_);
  or (_18953_, _18952_, _06261_);
  or (_18954_, _18953_, _18871_);
  or (_18956_, _18588_, _13769_);
  and (_18957_, _18956_, _13768_);
  nor (_18958_, _18957_, _10980_);
  and (_18959_, _18957_, _10980_);
  nor (_18960_, _18959_, _18958_);
  nor (_18961_, _18599_, _18592_);
  and (_18962_, _18961_, \oc8051_golden_model_1.PSW [7]);
  not (_18963_, _18962_);
  nor (_18964_, _18963_, _18960_);
  and (_18965_, _18963_, _18960_);
  or (_18967_, _18965_, _18964_);
  or (_18968_, _18967_, _06267_);
  and (_18969_, _18968_, _10307_);
  and (_18970_, _18969_, _18954_);
  or (_18971_, _18606_, _13887_);
  and (_18972_, _18971_, _13886_);
  nor (_18973_, _18972_, _11020_);
  and (_18974_, _18972_, _11020_);
  nor (_18975_, _18974_, _18973_);
  nor (_18976_, _18617_, _18610_);
  and (_18978_, _18976_, \oc8051_golden_model_1.PSW [7]);
  or (_18979_, _18978_, _18975_);
  nand (_18980_, _18978_, _18975_);
  and (_18981_, _18980_, _10306_);
  and (_18982_, _18981_, _18979_);
  or (_18983_, _18982_, _05676_);
  or (_18984_, _18983_, _18970_);
  nand (_18985_, _06084_, _05676_);
  and (_18986_, _18985_, _06027_);
  and (_18987_, _18986_, _18984_);
  or (_18989_, _18897_, _15326_);
  and (_18990_, _18989_, _06026_);
  and (_18991_, _18990_, _18899_);
  or (_18992_, _18991_, _09818_);
  or (_18993_, _18992_, _18987_);
  and (_18994_, _09178_, _07701_);
  or (_18995_, _18850_, _07012_);
  or (_18996_, _18995_, _18994_);
  or (_18997_, _18903_, _09827_);
  and (_18998_, _18997_, _05669_);
  and (_19000_, _18998_, _18996_);
  and (_19001_, _19000_, _18993_);
  or (_19002_, _19001_, _18856_);
  and (_19003_, _19002_, _12389_);
  nor (_19004_, _06084_, _05664_);
  not (_19005_, _09866_);
  nor (_19006_, _19005_, _09862_);
  and (_19007_, _19006_, _05662_);
  and (_19008_, _19007_, _09832_);
  or (_19009_, _19008_, _19004_);
  or (_19011_, _19009_, _19003_);
  and (_19012_, _19011_, _06020_);
  and (_19013_, _15389_, _07701_);
  or (_19014_, _19013_, _18850_);
  and (_19015_, _19014_, _06019_);
  or (_19016_, _19015_, _10661_);
  or (_19017_, _19016_, _19012_);
  nand (_19018_, _10661_, _06084_);
  and (_19019_, _19018_, _10675_);
  and (_19020_, _19019_, _19017_);
  or (_19022_, _19020_, _18853_);
  and (_19023_, _19022_, _18315_);
  and (_19024_, _10896_, _18314_);
  or (_19025_, _19024_, _19023_);
  and (_19026_, _19025_, _17671_);
  and (_19027_, _10896_, _17666_);
  or (_19028_, _19027_, _19026_);
  and (_19029_, _19028_, _17670_);
  and (_19030_, _10896_, _17503_);
  or (_19031_, _19030_, _19029_);
  and (_19033_, _19031_, _16972_);
  and (_19034_, _16971_, _10896_);
  or (_19035_, _19034_, _19033_);
  and (_19036_, _19035_, _16970_);
  and (_19037_, _10896_, _06650_);
  or (_19038_, _19037_, _19036_);
  and (_19039_, _19038_, _10686_);
  and (_19040_, _10685_, _10938_);
  or (_19041_, _19040_, _06282_);
  or (_19042_, _19041_, _19039_);
  or (_19044_, _10980_, _06283_);
  and (_19045_, _19044_, _10699_);
  and (_19046_, _19045_, _19042_);
  and (_19047_, _10698_, _11020_);
  or (_19048_, _19047_, _06112_);
  or (_19049_, _19048_, _19046_);
  and (_19050_, _19049_, _18852_);
  or (_19051_, _19050_, _06284_);
  or (_19052_, _18850_, _08756_);
  and (_19053_, _06093_, _05735_);
  not (_19055_, _19053_);
  and (_19056_, _19055_, _10725_);
  and (_19057_, _19056_, _19052_);
  and (_19058_, _19057_, _19051_);
  or (_19059_, _10893_, _10721_);
  and (_19060_, _19059_, _17104_);
  or (_19061_, _19060_, _19058_);
  and (_19062_, _19061_, _18848_);
  or (_19063_, _19062_, _10731_);
  or (_19064_, _10736_, _10935_);
  and (_19066_, _19064_, _10735_);
  and (_19067_, _19066_, _19063_);
  and (_19068_, _10977_, _06279_);
  or (_19069_, _19068_, _10741_);
  or (_19070_, _19069_, _19067_);
  or (_19071_, _10747_, _11017_);
  and (_19072_, _19071_, _07032_);
  and (_19073_, _19072_, _19070_);
  nand (_19074_, _19014_, _06108_);
  nor (_19075_, _19074_, _10979_);
  or (_19077_, _19075_, _10752_);
  or (_19078_, _19077_, _19073_);
  or (_19079_, _10895_, _17205_);
  and (_19080_, _19079_, _10760_);
  and (_19081_, _19080_, _19078_);
  and (_19082_, _10759_, _10895_);
  or (_19083_, _19082_, _10767_);
  or (_19084_, _19083_, _19081_);
  or (_19085_, _10766_, _10895_);
  and (_19086_, _19085_, _06668_);
  and (_19088_, _19086_, _19084_);
  and (_19089_, _10895_, _06667_);
  or (_19090_, _19089_, _10775_);
  or (_19091_, _19090_, _19088_);
  or (_19092_, _17395_, _10936_);
  and (_19093_, _19092_, _06291_);
  and (_19094_, _19093_, _19091_);
  nor (_19095_, _10979_, _06291_);
  or (_19096_, _19095_, _10781_);
  or (_19097_, _19096_, _19094_);
  nand (_19099_, _10781_, _11019_);
  and (_19100_, _19099_, _19097_);
  or (_19101_, _19100_, _06130_);
  and (_19102_, _15396_, _07701_);
  or (_19103_, _18850_, _08777_);
  or (_19104_, _19103_, _19102_);
  and (_19105_, _19104_, _10304_);
  and (_19106_, _19105_, _19101_);
  or (_19107_, _10297_, _10253_);
  nor (_19108_, _10304_, _10298_);
  and (_19110_, _19108_, _19107_);
  or (_19111_, _19110_, _17409_);
  or (_19112_, _19111_, _19106_);
  or (_19113_, _10815_, _10554_);
  and (_19114_, _19113_, _10816_);
  or (_19115_, _19114_, _17410_);
  and (_19116_, _19115_, _17423_);
  and (_19117_, _19116_, _19112_);
  nand (_19118_, _19114_, _17416_);
  nand (_19119_, _19118_, _06289_);
  or (_19121_, _19119_, _19117_);
  and (_19122_, _19121_, _18847_);
  or (_19123_, _10875_, _10626_);
  and (_19124_, _10876_, _10824_);
  and (_19125_, _19124_, _19123_);
  or (_19126_, _19125_, _10854_);
  or (_19127_, _19126_, _19122_);
  nand (_19128_, _10854_, _09906_);
  and (_19129_, _19128_, _10890_);
  and (_19130_, _19129_, _19127_);
  or (_19132_, _10924_, _10896_);
  and (_19133_, _19132_, _10925_);
  and (_19134_, _19133_, _16956_);
  or (_19135_, _19134_, _17437_);
  or (_19136_, _19135_, _19130_);
  nor (_19137_, _10965_, _10938_);
  nor (_19138_, _19137_, _10966_);
  and (_19139_, _19138_, _17443_);
  or (_19140_, _19139_, _10934_);
  and (_19141_, _19140_, _19136_);
  and (_19143_, _19138_, _06692_);
  or (_19144_, _19143_, _06051_);
  or (_19145_, _19144_, _19141_);
  and (_19146_, _19145_, _18842_);
  or (_19147_, _11046_, _11020_);
  and (_19148_, _11047_, _10974_);
  and (_19149_, _19148_, _19147_);
  or (_19150_, _19149_, _11015_);
  or (_19151_, _19150_, _19146_);
  and (_19152_, _19151_, _18838_);
  or (_19154_, _19152_, _06316_);
  or (_19155_, _18885_, _06718_);
  and (_19156_, _19155_, _11060_);
  and (_19157_, _19156_, _19154_);
  nor (_19158_, _11068_, _09861_);
  or (_19159_, _19158_, _11069_);
  and (_19160_, _19159_, _11059_);
  or (_19161_, _19160_, _11064_);
  or (_19162_, _19161_, _19157_);
  nand (_19163_, _11064_, _08393_);
  and (_19165_, _19163_, _05653_);
  and (_19166_, _19165_, _19162_);
  and (_19167_, _18921_, _05652_);
  or (_19168_, _19167_, _06047_);
  or (_19169_, _19168_, _19166_);
  and (_19170_, _15451_, _07701_);
  or (_19171_, _18850_, _06048_);
  or (_19172_, _19171_, _19170_);
  and (_19173_, _19172_, _11083_);
  and (_19174_, _19173_, _19169_);
  nor (_19176_, _11094_, \oc8051_golden_model_1.ACC [6]);
  nor (_19177_, _19176_, _11095_);
  and (_19178_, _19177_, _11082_);
  or (_19179_, _19178_, _11089_);
  or (_19180_, _19179_, _19174_);
  nand (_19181_, _11089_, _08393_);
  and (_19182_, _19181_, _01336_);
  and (_19183_, _19182_, _19180_);
  or (_19184_, _19183_, _18837_);
  and (_43339_, _19184_, _42882_);
  not (_19186_, \oc8051_golden_model_1.PCON [0]);
  nor (_19187_, _01336_, _19186_);
  nand (_19188_, _10995_, _07641_);
  nor (_19189_, _07641_, _19186_);
  nor (_19190_, _19189_, _06278_);
  nand (_19191_, _19190_, _19188_);
  and (_19192_, _09120_, _07641_);
  or (_19193_, _19189_, _07012_);
  or (_19194_, _19193_, _19192_);
  and (_19195_, _07641_, _06931_);
  nor (_19197_, _19195_, _19189_);
  nand (_19198_, _19197_, _09815_);
  nor (_19199_, _08127_, _11109_);
  or (_19200_, _19199_, _19189_);
  or (_19201_, _19200_, _06954_);
  and (_19202_, _07641_, \oc8051_golden_model_1.ACC [0]);
  nor (_19203_, _19202_, _19189_);
  nor (_19204_, _19203_, _06939_);
  nor (_19205_, _06938_, _19186_);
  or (_19206_, _19205_, _06102_);
  or (_19208_, _19206_, _19204_);
  and (_19209_, _19208_, _06848_);
  and (_19210_, _19209_, _19201_);
  nor (_19211_, _19197_, _06848_);
  or (_19212_, _19211_, _19210_);
  nand (_19213_, _19212_, _06220_);
  or (_19214_, _19203_, _06220_);
  and (_19215_, _19214_, _09817_);
  nand (_19216_, _19215_, _19213_);
  and (_19217_, _19216_, _19198_);
  and (_19219_, _19217_, _19194_);
  or (_19220_, _19219_, _09833_);
  and (_19221_, _14186_, _07641_);
  or (_19222_, _19221_, _19189_);
  or (_19223_, _19222_, _05669_);
  and (_19224_, _19223_, _06020_);
  and (_19225_, _19224_, _19220_);
  and (_19226_, _07641_, _08672_);
  or (_19227_, _19226_, _19189_);
  and (_19228_, _19227_, _06019_);
  or (_19230_, _19228_, _06112_);
  or (_19231_, _19230_, _19225_);
  and (_19232_, _14086_, _07641_);
  or (_19233_, _19189_, _08751_);
  or (_19234_, _19233_, _19232_);
  and (_19235_, _19234_, _08756_);
  and (_19236_, _19235_, _19231_);
  nor (_19237_, _12302_, _11109_);
  or (_19238_, _19237_, _19189_);
  and (_19239_, _19188_, _06284_);
  and (_19241_, _19239_, _19238_);
  or (_19242_, _19241_, _19236_);
  and (_19243_, _19242_, _07032_);
  nand (_19244_, _19227_, _06108_);
  nor (_19245_, _19244_, _19199_);
  or (_19246_, _19245_, _06277_);
  or (_19247_, _19246_, _19243_);
  and (_19248_, _19247_, _19191_);
  or (_19249_, _19248_, _06130_);
  and (_19250_, _14083_, _07641_);
  or (_19252_, _19189_, _08777_);
  or (_19253_, _19252_, _19250_);
  and (_19254_, _19253_, _08782_);
  and (_19255_, _19254_, _19249_);
  not (_19256_, _06408_);
  and (_19257_, _19238_, _06292_);
  or (_19258_, _19257_, _19256_);
  or (_19259_, _19258_, _19255_);
  or (_19260_, _19200_, _06408_);
  and (_19261_, _19260_, _01336_);
  and (_19263_, _19261_, _19259_);
  or (_19264_, _19263_, _19187_);
  and (_43340_, _19264_, _42882_);
  not (_19265_, \oc8051_golden_model_1.PCON [1]);
  nor (_19266_, _01336_, _19265_);
  and (_19267_, _09075_, _07641_);
  nor (_19268_, _07641_, _19265_);
  or (_19269_, _19268_, _07012_);
  or (_19270_, _19269_, _19267_);
  or (_19271_, _07641_, \oc8051_golden_model_1.PCON [1]);
  and (_19273_, _14284_, _07641_);
  not (_19274_, _19273_);
  and (_19275_, _19274_, _19271_);
  or (_19276_, _19275_, _06954_);
  and (_19277_, _07641_, \oc8051_golden_model_1.ACC [1]);
  or (_19278_, _19277_, _19268_);
  and (_19279_, _19278_, _06938_);
  nor (_19280_, _06938_, _19265_);
  or (_19281_, _19280_, _06102_);
  or (_19282_, _19281_, _19279_);
  and (_19284_, _19282_, _06848_);
  and (_19285_, _19284_, _19276_);
  nor (_19286_, _11109_, _07132_);
  or (_19287_, _19286_, _19268_);
  and (_19288_, _19287_, _06239_);
  or (_19289_, _19288_, _19285_);
  and (_19290_, _19289_, _06220_);
  and (_19291_, _19278_, _06219_);
  or (_19292_, _19291_, _09818_);
  or (_19293_, _19292_, _19290_);
  or (_19295_, _19287_, _09827_);
  and (_19296_, _19295_, _05669_);
  and (_19297_, _19296_, _19293_);
  and (_19298_, _19297_, _19270_);
  or (_19299_, _14367_, _11109_);
  and (_19300_, _19271_, _09833_);
  and (_19301_, _19300_, _19299_);
  or (_19302_, _19301_, _19298_);
  and (_19303_, _19302_, _06020_);
  nand (_19304_, _07641_, _06832_);
  and (_19306_, _19271_, _06019_);
  and (_19307_, _19306_, _19304_);
  or (_19308_, _19307_, _19303_);
  and (_19309_, _19308_, _08751_);
  or (_19310_, _14263_, _11109_);
  and (_19311_, _19271_, _06112_);
  and (_19312_, _19311_, _19310_);
  or (_19313_, _19312_, _06284_);
  or (_19314_, _19313_, _19309_);
  and (_19315_, _10994_, _07641_);
  or (_19317_, _19315_, _19268_);
  or (_19318_, _19317_, _08756_);
  and (_19319_, _19318_, _07032_);
  and (_19320_, _19319_, _19314_);
  or (_19321_, _14261_, _11109_);
  and (_19322_, _19271_, _06108_);
  and (_19323_, _19322_, _19321_);
  or (_19324_, _19323_, _06277_);
  or (_19325_, _19324_, _19320_);
  and (_19326_, _19277_, _08078_);
  or (_19328_, _19268_, _06278_);
  or (_19329_, _19328_, _19326_);
  and (_19330_, _19329_, _08777_);
  and (_19331_, _19330_, _19325_);
  or (_19332_, _19304_, _08078_);
  and (_19333_, _19271_, _06130_);
  and (_19334_, _19333_, _19332_);
  or (_19335_, _19334_, _06292_);
  or (_19336_, _19335_, _19331_);
  nor (_19337_, _10993_, _11109_);
  or (_19339_, _19337_, _19268_);
  or (_19340_, _19339_, _08782_);
  and (_19341_, _19340_, _06718_);
  and (_19342_, _19341_, _19336_);
  and (_19343_, _19275_, _06316_);
  or (_19344_, _19343_, _06047_);
  or (_19345_, _19344_, _19342_);
  or (_19346_, _19268_, _06048_);
  or (_19347_, _19346_, _19273_);
  and (_19348_, _19347_, _01336_);
  and (_19350_, _19348_, _19345_);
  or (_19351_, _19350_, _19266_);
  and (_43342_, _19351_, _42882_);
  not (_19352_, \oc8051_golden_model_1.PCON [2]);
  nor (_19353_, _01336_, _19352_);
  and (_19354_, _09182_, _07641_);
  nor (_19355_, _07641_, _19352_);
  or (_19356_, _19355_, _07012_);
  or (_19357_, _19356_, _19354_);
  nor (_19358_, _11109_, _07530_);
  nor (_19360_, _19358_, _19355_);
  nand (_19361_, _19360_, _09815_);
  and (_19362_, _14493_, _07641_);
  or (_19363_, _19362_, _19355_);
  or (_19364_, _19363_, _06954_);
  and (_19365_, _07641_, \oc8051_golden_model_1.ACC [2]);
  nor (_19366_, _19365_, _19355_);
  nor (_19367_, _19366_, _06939_);
  nor (_19368_, _06938_, _19352_);
  or (_19369_, _19368_, _06102_);
  or (_19371_, _19369_, _19367_);
  and (_19372_, _19371_, _06848_);
  and (_19373_, _19372_, _19364_);
  nor (_19374_, _19360_, _06848_);
  or (_19375_, _19374_, _19373_);
  nand (_19376_, _19375_, _06220_);
  or (_19377_, _19366_, _06220_);
  and (_19378_, _19377_, _09817_);
  nand (_19379_, _19378_, _19376_);
  and (_19380_, _19379_, _19361_);
  and (_19382_, _19380_, _19357_);
  or (_19383_, _19382_, _09833_);
  and (_19384_, _14580_, _07641_);
  or (_19385_, _19384_, _19355_);
  or (_19386_, _19385_, _05669_);
  and (_19387_, _19386_, _06020_);
  and (_19388_, _19387_, _19383_);
  and (_19389_, _07641_, _08730_);
  or (_19390_, _19389_, _19355_);
  and (_19391_, _19390_, _06019_);
  or (_19393_, _19391_, _06112_);
  or (_19394_, _19393_, _19388_);
  and (_19395_, _14596_, _07641_);
  or (_19396_, _19355_, _08751_);
  or (_19397_, _19396_, _19395_);
  and (_19398_, _19397_, _08756_);
  and (_19399_, _19398_, _19394_);
  and (_19400_, _10991_, _07641_);
  or (_19401_, _19400_, _19355_);
  and (_19402_, _19401_, _06284_);
  or (_19404_, _19402_, _19399_);
  and (_19405_, _19404_, _07032_);
  or (_19406_, _19355_, _08177_);
  and (_19407_, _19390_, _06108_);
  and (_19408_, _19407_, _19406_);
  or (_19409_, _19408_, _19405_);
  and (_19410_, _19409_, _06278_);
  nor (_19411_, _19366_, _06278_);
  and (_19412_, _19411_, _19406_);
  or (_19413_, _19412_, _06130_);
  or (_19415_, _19413_, _19410_);
  and (_19416_, _14593_, _07641_);
  or (_19417_, _19355_, _08777_);
  or (_19418_, _19417_, _19416_);
  and (_19419_, _19418_, _08782_);
  and (_19420_, _19419_, _19415_);
  nor (_19421_, _10990_, _11109_);
  or (_19422_, _19421_, _19355_);
  and (_19423_, _19422_, _06292_);
  or (_19424_, _19423_, _19420_);
  and (_19426_, _19424_, _06718_);
  and (_19427_, _19363_, _06316_);
  or (_19428_, _19427_, _06047_);
  or (_19429_, _19428_, _19426_);
  and (_19430_, _14657_, _07641_);
  or (_19431_, _19355_, _06048_);
  or (_19432_, _19431_, _19430_);
  and (_19433_, _19432_, _01336_);
  and (_19434_, _19433_, _19429_);
  or (_19435_, _19434_, _19353_);
  and (_43343_, _19435_, _42882_);
  not (_19437_, \oc8051_golden_model_1.PCON [3]);
  nor (_19438_, _01336_, _19437_);
  nor (_19439_, _07641_, _19437_);
  or (_19440_, _19439_, _08029_);
  and (_19441_, _07641_, _08662_);
  or (_19442_, _19441_, _19439_);
  and (_19443_, _19442_, _06108_);
  and (_19444_, _19443_, _19440_);
  and (_19445_, _09181_, _07641_);
  or (_19447_, _19439_, _07012_);
  or (_19448_, _19447_, _19445_);
  nor (_19449_, _11109_, _07353_);
  nor (_19450_, _19449_, _19439_);
  nand (_19451_, _19450_, _09815_);
  and (_19452_, _14672_, _07641_);
  or (_19453_, _19452_, _19439_);
  or (_19454_, _19453_, _06954_);
  and (_19455_, _07641_, \oc8051_golden_model_1.ACC [3]);
  nor (_19456_, _19455_, _19439_);
  nor (_19458_, _19456_, _06939_);
  nor (_19459_, _06938_, _19437_);
  or (_19460_, _19459_, _06102_);
  or (_19461_, _19460_, _19458_);
  and (_19462_, _19461_, _06848_);
  and (_19463_, _19462_, _19454_);
  nor (_19464_, _19450_, _06848_);
  or (_19465_, _19464_, _19463_);
  nand (_19466_, _19465_, _06220_);
  or (_19467_, _19456_, _06220_);
  and (_19469_, _19467_, _09817_);
  nand (_19470_, _19469_, _19466_);
  and (_19471_, _19470_, _19451_);
  and (_19472_, _19471_, _19448_);
  or (_19473_, _19472_, _09833_);
  and (_19474_, _14778_, _07641_);
  or (_19475_, _19474_, _19439_);
  or (_19476_, _19475_, _05669_);
  and (_19477_, _19476_, _06020_);
  and (_19478_, _19477_, _19473_);
  and (_19480_, _19442_, _06019_);
  or (_19481_, _19480_, _06112_);
  or (_19482_, _19481_, _19478_);
  and (_19483_, _14793_, _07641_);
  or (_19484_, _19483_, _19439_);
  or (_19485_, _19484_, _08751_);
  and (_19486_, _19485_, _08756_);
  and (_19487_, _19486_, _19482_);
  and (_19488_, _12299_, _07641_);
  or (_19489_, _19488_, _19439_);
  and (_19491_, _19489_, _06284_);
  or (_19492_, _19491_, _19487_);
  and (_19493_, _19492_, _07032_);
  or (_19494_, _19493_, _19444_);
  and (_19495_, _19494_, _06278_);
  nor (_19496_, _19456_, _06278_);
  and (_19497_, _19496_, _19440_);
  or (_19498_, _19497_, _06130_);
  or (_19499_, _19498_, _19495_);
  and (_19500_, _14792_, _07641_);
  or (_19502_, _19439_, _08777_);
  or (_19503_, _19502_, _19500_);
  and (_19504_, _19503_, _08782_);
  and (_19505_, _19504_, _19499_);
  nor (_19506_, _10988_, _11109_);
  or (_19507_, _19506_, _19439_);
  and (_19508_, _19507_, _06292_);
  or (_19509_, _19508_, _19505_);
  and (_19510_, _19509_, _06718_);
  and (_19511_, _19453_, _06316_);
  or (_19513_, _19511_, _06047_);
  or (_19514_, _19513_, _19510_);
  and (_19515_, _14849_, _07641_);
  or (_19516_, _19439_, _06048_);
  or (_19517_, _19516_, _19515_);
  and (_19518_, _19517_, _01336_);
  and (_19519_, _19518_, _19514_);
  or (_19520_, _19519_, _19438_);
  and (_43344_, _19520_, _42882_);
  not (_19521_, \oc8051_golden_model_1.PCON [4]);
  nor (_19523_, _01336_, _19521_);
  nor (_19524_, _07641_, _19521_);
  or (_19525_, _19524_, _08273_);
  and (_19526_, _08665_, _07641_);
  or (_19527_, _19526_, _19524_);
  and (_19528_, _19527_, _06108_);
  and (_19529_, _19528_, _19525_);
  or (_19530_, _19527_, _06020_);
  and (_19531_, _14887_, _07641_);
  or (_19532_, _19531_, _19524_);
  or (_19534_, _19532_, _06954_);
  and (_19535_, _07641_, \oc8051_golden_model_1.ACC [4]);
  or (_19536_, _19535_, _19524_);
  and (_19537_, _19536_, _06938_);
  nor (_19538_, _06938_, _19521_);
  or (_19539_, _19538_, _06102_);
  or (_19540_, _19539_, _19537_);
  and (_19541_, _19540_, _06848_);
  and (_19542_, _19541_, _19534_);
  nor (_19543_, _08270_, _11109_);
  or (_19545_, _19543_, _19524_);
  and (_19546_, _19545_, _06239_);
  or (_19547_, _19546_, _19542_);
  and (_19548_, _19547_, _06220_);
  and (_19549_, _19536_, _06219_);
  or (_19550_, _19549_, _09818_);
  or (_19551_, _19550_, _19548_);
  and (_19552_, _09180_, _07641_);
  or (_19553_, _19524_, _07012_);
  or (_19554_, _19553_, _19552_);
  or (_19556_, _19545_, _09827_);
  and (_19557_, _19556_, _05669_);
  and (_19558_, _19557_, _19554_);
  and (_19559_, _19558_, _19551_);
  and (_19560_, _14983_, _07641_);
  or (_19561_, _19560_, _19524_);
  and (_19562_, _19561_, _09833_);
  or (_19563_, _19562_, _06019_);
  or (_19564_, _19563_, _19559_);
  and (_19565_, _19564_, _19530_);
  or (_19567_, _19565_, _06112_);
  and (_19568_, _14876_, _07641_);
  or (_19569_, _19524_, _08751_);
  or (_19570_, _19569_, _19568_);
  and (_19571_, _19570_, _08756_);
  and (_19572_, _19571_, _19567_);
  and (_19573_, _10986_, _07641_);
  or (_19574_, _19573_, _19524_);
  and (_19575_, _19574_, _06284_);
  or (_19576_, _19575_, _19572_);
  and (_19578_, _19576_, _07032_);
  or (_19579_, _19578_, _19529_);
  and (_19580_, _19579_, _06278_);
  and (_19581_, _19536_, _06277_);
  and (_19582_, _19581_, _19525_);
  or (_19583_, _19582_, _06130_);
  or (_19584_, _19583_, _19580_);
  and (_19585_, _14873_, _07641_);
  or (_19586_, _19524_, _08777_);
  or (_19587_, _19586_, _19585_);
  and (_19589_, _19587_, _08782_);
  and (_19590_, _19589_, _19584_);
  nor (_19591_, _10985_, _11109_);
  or (_19592_, _19591_, _19524_);
  and (_19593_, _19592_, _06292_);
  or (_19594_, _19593_, _19590_);
  and (_19595_, _19594_, _06718_);
  and (_19596_, _19532_, _06316_);
  or (_19597_, _19596_, _06047_);
  or (_19598_, _19597_, _19595_);
  and (_19600_, _15055_, _07641_);
  or (_19601_, _19524_, _06048_);
  or (_19602_, _19601_, _19600_);
  and (_19603_, _19602_, _01336_);
  and (_19604_, _19603_, _19598_);
  or (_19605_, _19604_, _19523_);
  and (_43345_, _19605_, _42882_);
  not (_19606_, \oc8051_golden_model_1.PCON [5]);
  nor (_19607_, _01336_, _19606_);
  nor (_19608_, _07641_, _19606_);
  and (_19610_, _08652_, _07641_);
  or (_19611_, _19610_, _19608_);
  or (_19612_, _19611_, _06020_);
  and (_19613_, _15093_, _07641_);
  or (_19614_, _19613_, _19608_);
  or (_19615_, _19614_, _06954_);
  and (_19616_, _07641_, \oc8051_golden_model_1.ACC [5]);
  or (_19617_, _19616_, _19608_);
  and (_19618_, _19617_, _06938_);
  nor (_19619_, _06938_, _19606_);
  or (_19621_, _19619_, _06102_);
  or (_19622_, _19621_, _19618_);
  and (_19623_, _19622_, _06848_);
  and (_19624_, _19623_, _19615_);
  nor (_19625_, _07977_, _11109_);
  or (_19626_, _19625_, _19608_);
  and (_19627_, _19626_, _06239_);
  or (_19628_, _19627_, _19624_);
  and (_19629_, _19628_, _06220_);
  and (_19630_, _19617_, _06219_);
  or (_19632_, _19630_, _09818_);
  or (_19633_, _19632_, _19629_);
  and (_19634_, _09179_, _07641_);
  or (_19635_, _19608_, _07012_);
  or (_19636_, _19635_, _19634_);
  or (_19637_, _19626_, _09827_);
  and (_19638_, _19637_, _05669_);
  and (_19639_, _19638_, _19636_);
  and (_19640_, _19639_, _19633_);
  and (_19641_, _15179_, _07641_);
  or (_19643_, _19641_, _19608_);
  and (_19644_, _19643_, _09833_);
  or (_19645_, _19644_, _06019_);
  or (_19646_, _19645_, _19640_);
  and (_19647_, _19646_, _19612_);
  or (_19648_, _19647_, _06112_);
  and (_19649_, _15195_, _07641_);
  or (_19650_, _19649_, _19608_);
  or (_19651_, _19650_, _08751_);
  and (_19652_, _19651_, _08756_);
  and (_19654_, _19652_, _19648_);
  and (_19655_, _12306_, _07641_);
  or (_19656_, _19655_, _19608_);
  and (_19657_, _19656_, _06284_);
  or (_19658_, _19657_, _19654_);
  and (_19659_, _19658_, _07032_);
  or (_19660_, _19608_, _07980_);
  and (_19661_, _19611_, _06108_);
  and (_19662_, _19661_, _19660_);
  or (_19663_, _19662_, _19659_);
  and (_19665_, _19663_, _06278_);
  and (_19666_, _19617_, _06277_);
  and (_19667_, _19666_, _19660_);
  or (_19668_, _19667_, _06130_);
  or (_19669_, _19668_, _19665_);
  and (_19670_, _15194_, _07641_);
  or (_19671_, _19608_, _08777_);
  or (_19672_, _19671_, _19670_);
  and (_19673_, _19672_, _08782_);
  and (_19674_, _19673_, _19669_);
  nor (_19676_, _10982_, _11109_);
  or (_19677_, _19676_, _19608_);
  and (_19678_, _19677_, _06292_);
  or (_19679_, _19678_, _19674_);
  and (_19680_, _19679_, _06718_);
  and (_19681_, _19614_, _06316_);
  or (_19682_, _19681_, _06047_);
  or (_19683_, _19682_, _19680_);
  and (_19684_, _15253_, _07641_);
  or (_19685_, _19608_, _06048_);
  or (_19687_, _19685_, _19684_);
  and (_19688_, _19687_, _01336_);
  and (_19689_, _19688_, _19683_);
  or (_19690_, _19689_, _19607_);
  and (_43346_, _19690_, _42882_);
  not (_19691_, \oc8051_golden_model_1.PCON [6]);
  nor (_19692_, _01336_, _19691_);
  nor (_19693_, _07641_, _19691_);
  and (_19694_, _15389_, _07641_);
  or (_19695_, _19694_, _19693_);
  or (_19697_, _19695_, _06020_);
  and (_19698_, _15293_, _07641_);
  or (_19699_, _19698_, _19693_);
  or (_19700_, _19699_, _06954_);
  and (_19701_, _07641_, \oc8051_golden_model_1.ACC [6]);
  or (_19702_, _19701_, _19693_);
  and (_19703_, _19702_, _06938_);
  nor (_19704_, _06938_, _19691_);
  or (_19705_, _19704_, _06102_);
  or (_19706_, _19705_, _19703_);
  and (_19708_, _19706_, _06848_);
  and (_19709_, _19708_, _19700_);
  nor (_19710_, _07883_, _11109_);
  or (_19711_, _19710_, _19693_);
  and (_19712_, _19711_, _06239_);
  or (_19713_, _19712_, _19709_);
  and (_19714_, _19713_, _06220_);
  and (_19715_, _19702_, _06219_);
  or (_19716_, _19715_, _09818_);
  or (_19717_, _19716_, _19714_);
  and (_19719_, _09178_, _07641_);
  or (_19720_, _19693_, _07012_);
  or (_19721_, _19720_, _19719_);
  or (_19722_, _19711_, _09827_);
  and (_19723_, _19722_, _05669_);
  and (_19724_, _19723_, _19721_);
  and (_19725_, _19724_, _19717_);
  and (_19726_, _15382_, _07641_);
  or (_19727_, _19726_, _19693_);
  and (_19728_, _19727_, _09833_);
  or (_19730_, _19728_, _06019_);
  or (_19731_, _19730_, _19725_);
  and (_19732_, _19731_, _19697_);
  or (_19733_, _19732_, _06112_);
  and (_19734_, _15399_, _07641_);
  or (_19735_, _19734_, _19693_);
  or (_19736_, _19735_, _08751_);
  and (_19737_, _19736_, _08756_);
  and (_19738_, _19737_, _19733_);
  and (_19739_, _10980_, _07641_);
  or (_19741_, _19739_, _19693_);
  and (_19742_, _19741_, _06284_);
  or (_19743_, _19742_, _19738_);
  and (_19744_, _19743_, _07032_);
  or (_19745_, _19693_, _07886_);
  and (_19746_, _19695_, _06108_);
  and (_19747_, _19746_, _19745_);
  or (_19748_, _19747_, _19744_);
  and (_19749_, _19748_, _06278_);
  and (_19750_, _19702_, _06277_);
  and (_19752_, _19750_, _19745_);
  or (_19753_, _19752_, _06130_);
  or (_19754_, _19753_, _19749_);
  and (_19755_, _15396_, _07641_);
  or (_19756_, _19693_, _08777_);
  or (_19757_, _19756_, _19755_);
  and (_19758_, _19757_, _08782_);
  and (_19759_, _19758_, _19754_);
  nor (_19760_, _10979_, _11109_);
  or (_19761_, _19760_, _19693_);
  and (_19763_, _19761_, _06292_);
  or (_19764_, _19763_, _19759_);
  and (_19765_, _19764_, _06718_);
  and (_19766_, _19699_, _06316_);
  or (_19767_, _19766_, _06047_);
  or (_19768_, _19767_, _19765_);
  and (_19769_, _15451_, _07641_);
  or (_19770_, _19693_, _06048_);
  or (_19771_, _19770_, _19769_);
  and (_19772_, _19771_, _01336_);
  and (_19774_, _19772_, _19768_);
  or (_19775_, _19774_, _19692_);
  and (_43347_, _19775_, _42882_);
  not (_19776_, \oc8051_golden_model_1.TMOD [0]);
  nor (_19777_, _01336_, _19776_);
  nand (_19778_, _10995_, _07653_);
  nor (_19779_, _07653_, _19776_);
  nor (_19780_, _19779_, _06278_);
  nand (_19781_, _19780_, _19778_);
  and (_19782_, _09120_, _07653_);
  or (_19784_, _19779_, _07012_);
  or (_19785_, _19784_, _19782_);
  and (_19786_, _07653_, _06931_);
  nor (_19787_, _19786_, _19779_);
  nand (_19788_, _19787_, _09815_);
  nor (_19789_, _08127_, _11185_);
  or (_19790_, _19789_, _19779_);
  or (_19791_, _19790_, _06954_);
  and (_19792_, _07653_, \oc8051_golden_model_1.ACC [0]);
  nor (_19793_, _19792_, _19779_);
  nor (_19795_, _19793_, _06939_);
  nor (_19796_, _06938_, _19776_);
  or (_19797_, _19796_, _06102_);
  or (_19798_, _19797_, _19795_);
  and (_19799_, _19798_, _06848_);
  and (_19800_, _19799_, _19791_);
  nor (_19801_, _19787_, _06848_);
  or (_19802_, _19801_, _19800_);
  nand (_19803_, _19802_, _06220_);
  or (_19804_, _19793_, _06220_);
  and (_19806_, _19804_, _09817_);
  nand (_19807_, _19806_, _19803_);
  and (_19808_, _19807_, _19788_);
  and (_19809_, _19808_, _19785_);
  or (_19810_, _19809_, _09833_);
  and (_19811_, _14186_, _07653_);
  or (_19812_, _19811_, _19779_);
  or (_19813_, _19812_, _05669_);
  and (_19814_, _19813_, _06020_);
  and (_19815_, _19814_, _19810_);
  and (_19817_, _07653_, _08672_);
  or (_19818_, _19817_, _19779_);
  and (_19819_, _19818_, _06019_);
  or (_19820_, _19819_, _06112_);
  or (_19821_, _19820_, _19815_);
  and (_19822_, _14086_, _07653_);
  or (_19823_, _19779_, _08751_);
  or (_19824_, _19823_, _19822_);
  and (_19825_, _19824_, _08756_);
  and (_19826_, _19825_, _19821_);
  nor (_19828_, _12302_, _11185_);
  or (_19829_, _19828_, _19779_);
  and (_19830_, _19778_, _06284_);
  and (_19831_, _19830_, _19829_);
  or (_19832_, _19831_, _19826_);
  and (_19833_, _19832_, _07032_);
  nand (_19834_, _19818_, _06108_);
  nor (_19835_, _19834_, _19789_);
  or (_19836_, _19835_, _06277_);
  or (_19837_, _19836_, _19833_);
  and (_19839_, _19837_, _19781_);
  or (_19840_, _19839_, _06130_);
  and (_19841_, _14083_, _07653_);
  or (_19842_, _19779_, _08777_);
  or (_19843_, _19842_, _19841_);
  and (_19844_, _19843_, _08782_);
  and (_19845_, _19844_, _19840_);
  and (_19846_, _19829_, _06292_);
  or (_19847_, _19846_, _19256_);
  or (_19848_, _19847_, _19845_);
  or (_19850_, _19790_, _06408_);
  and (_19851_, _19850_, _01336_);
  and (_19852_, _19851_, _19848_);
  or (_19853_, _19852_, _19777_);
  and (_43349_, _19853_, _42882_);
  and (_19854_, _01340_, \oc8051_golden_model_1.TMOD [1]);
  or (_19855_, _14367_, _11185_);
  or (_19856_, _07653_, \oc8051_golden_model_1.TMOD [1]);
  and (_19857_, _19856_, _09833_);
  and (_19858_, _19857_, _19855_);
  and (_19861_, _09075_, _07653_);
  and (_19862_, _11185_, \oc8051_golden_model_1.TMOD [1]);
  or (_19863_, _19862_, _07012_);
  or (_19864_, _19863_, _19861_);
  and (_19865_, _14284_, _07653_);
  not (_19866_, _19865_);
  and (_19867_, _19866_, _19856_);
  or (_19868_, _19867_, _06954_);
  and (_19869_, _07653_, \oc8051_golden_model_1.ACC [1]);
  or (_19870_, _19869_, _19862_);
  and (_19873_, _19870_, _06938_);
  and (_19874_, _06939_, \oc8051_golden_model_1.TMOD [1]);
  or (_19875_, _19874_, _06102_);
  or (_19876_, _19875_, _19873_);
  and (_19877_, _19876_, _06848_);
  and (_19878_, _19877_, _19868_);
  nor (_19879_, _11185_, _07132_);
  or (_19880_, _19879_, _19862_);
  and (_19881_, _19880_, _06239_);
  or (_19882_, _19881_, _19878_);
  and (_19885_, _19882_, _06220_);
  and (_19886_, _19870_, _06219_);
  or (_19887_, _19886_, _09818_);
  or (_19888_, _19887_, _19885_);
  or (_19889_, _19880_, _09827_);
  and (_19890_, _19889_, _05669_);
  and (_19891_, _19890_, _19888_);
  and (_19892_, _19891_, _19864_);
  or (_19893_, _19892_, _19858_);
  and (_19894_, _19893_, _06020_);
  nand (_19897_, _07653_, _06832_);
  and (_19898_, _19856_, _06019_);
  and (_19899_, _19898_, _19897_);
  or (_19900_, _19899_, _19894_);
  and (_19901_, _19900_, _08751_);
  or (_19902_, _14263_, _11185_);
  and (_19903_, _19856_, _06112_);
  and (_19904_, _19903_, _19902_);
  or (_19905_, _19904_, _06284_);
  or (_19906_, _19905_, _19901_);
  and (_19909_, _10994_, _07653_);
  or (_19910_, _19909_, _19862_);
  or (_19911_, _19910_, _08756_);
  and (_19912_, _19911_, _07032_);
  and (_19913_, _19912_, _19906_);
  or (_19914_, _14261_, _11185_);
  and (_19915_, _19856_, _06108_);
  and (_19916_, _19915_, _19914_);
  or (_19917_, _19916_, _06277_);
  or (_19918_, _19917_, _19913_);
  and (_19921_, _19869_, _08078_);
  or (_19922_, _19862_, _06278_);
  or (_19923_, _19922_, _19921_);
  and (_19924_, _19923_, _08777_);
  and (_19925_, _19924_, _19918_);
  or (_19926_, _19897_, _08078_);
  and (_19927_, _19856_, _06130_);
  and (_19928_, _19927_, _19926_);
  or (_19929_, _19928_, _06292_);
  or (_19930_, _19929_, _19925_);
  nor (_19933_, _10993_, _11185_);
  or (_19934_, _19933_, _19862_);
  or (_19935_, _19934_, _08782_);
  and (_19936_, _19935_, _06718_);
  and (_19937_, _19936_, _19930_);
  and (_19938_, _19867_, _06316_);
  or (_19939_, _19938_, _06047_);
  or (_19940_, _19939_, _19937_);
  or (_19941_, _19862_, _06048_);
  or (_19942_, _19941_, _19865_);
  and (_19944_, _19942_, _01336_);
  and (_19945_, _19944_, _19940_);
  or (_19946_, _19945_, _19854_);
  and (_43350_, _19946_, _42882_);
  not (_19947_, \oc8051_golden_model_1.TMOD [2]);
  nor (_19948_, _01336_, _19947_);
  nor (_19949_, _07653_, _19947_);
  or (_19950_, _19949_, _08177_);
  and (_19951_, _07653_, _08730_);
  or (_19952_, _19951_, _19949_);
  and (_19954_, _19952_, _06108_);
  and (_19955_, _19954_, _19950_);
  and (_19956_, _09182_, _07653_);
  or (_19957_, _19949_, _07012_);
  or (_19958_, _19957_, _19956_);
  nor (_19959_, _11185_, _07530_);
  nor (_19960_, _19959_, _19949_);
  nand (_19961_, _19960_, _09815_);
  and (_19962_, _14493_, _07653_);
  or (_19963_, _19962_, _19949_);
  or (_19965_, _19963_, _06954_);
  and (_19966_, _07653_, \oc8051_golden_model_1.ACC [2]);
  nor (_19967_, _19966_, _19949_);
  nor (_19968_, _19967_, _06939_);
  nor (_19969_, _06938_, _19947_);
  or (_19970_, _19969_, _06102_);
  or (_19971_, _19970_, _19968_);
  and (_19972_, _19971_, _06848_);
  and (_19973_, _19972_, _19965_);
  nor (_19974_, _19960_, _06848_);
  or (_19976_, _19974_, _19973_);
  nand (_19977_, _19976_, _06220_);
  or (_19978_, _19967_, _06220_);
  and (_19979_, _19978_, _09817_);
  nand (_19980_, _19979_, _19977_);
  and (_19981_, _19980_, _19961_);
  and (_19982_, _19981_, _19958_);
  or (_19983_, _19982_, _09833_);
  and (_19984_, _14580_, _07653_);
  or (_19985_, _19984_, _19949_);
  or (_19987_, _19985_, _05669_);
  and (_19988_, _19987_, _06020_);
  and (_19989_, _19988_, _19983_);
  and (_19990_, _19952_, _06019_);
  or (_19991_, _19990_, _06112_);
  or (_19992_, _19991_, _19989_);
  and (_19993_, _14596_, _07653_);
  or (_19994_, _19993_, _19949_);
  or (_19995_, _19994_, _08751_);
  and (_19996_, _19995_, _08756_);
  and (_19998_, _19996_, _19992_);
  and (_19999_, _10991_, _07653_);
  or (_20000_, _19999_, _19949_);
  and (_20001_, _20000_, _06284_);
  or (_20002_, _20001_, _19998_);
  and (_20003_, _20002_, _07032_);
  or (_20004_, _20003_, _19955_);
  and (_20005_, _20004_, _06278_);
  nor (_20006_, _19967_, _06278_);
  and (_20007_, _20006_, _19950_);
  or (_20009_, _20007_, _06130_);
  or (_20010_, _20009_, _20005_);
  and (_20011_, _14593_, _07653_);
  or (_20012_, _19949_, _08777_);
  or (_20013_, _20012_, _20011_);
  and (_20014_, _20013_, _08782_);
  and (_20015_, _20014_, _20010_);
  nor (_20016_, _10990_, _11185_);
  or (_20017_, _20016_, _19949_);
  and (_20018_, _20017_, _06292_);
  or (_20020_, _20018_, _20015_);
  and (_20021_, _20020_, _06718_);
  and (_20022_, _19963_, _06316_);
  or (_20023_, _20022_, _06047_);
  or (_20024_, _20023_, _20021_);
  and (_20025_, _14657_, _07653_);
  or (_20026_, _19949_, _06048_);
  or (_20027_, _20026_, _20025_);
  and (_20028_, _20027_, _01336_);
  and (_20029_, _20028_, _20024_);
  or (_20031_, _20029_, _19948_);
  and (_43351_, _20031_, _42882_);
  and (_20032_, _01340_, \oc8051_golden_model_1.TMOD [3]);
  and (_20033_, _11185_, \oc8051_golden_model_1.TMOD [3]);
  or (_20034_, _20033_, _08029_);
  and (_20035_, _07653_, _08662_);
  or (_20036_, _20035_, _20033_);
  and (_20037_, _20036_, _06108_);
  and (_20038_, _20037_, _20034_);
  or (_20039_, _20036_, _06020_);
  and (_20041_, _09181_, _07653_);
  or (_20042_, _20033_, _07012_);
  or (_20043_, _20042_, _20041_);
  and (_20044_, _14672_, _07653_);
  or (_20045_, _20044_, _20033_);
  or (_20046_, _20045_, _06954_);
  and (_20047_, _07653_, \oc8051_golden_model_1.ACC [3]);
  or (_20048_, _20047_, _20033_);
  and (_20049_, _20048_, _06938_);
  and (_20050_, _06939_, \oc8051_golden_model_1.TMOD [3]);
  or (_20052_, _20050_, _06102_);
  or (_20053_, _20052_, _20049_);
  and (_20054_, _20053_, _06848_);
  and (_20055_, _20054_, _20046_);
  nor (_20056_, _11185_, _07353_);
  or (_20057_, _20056_, _20033_);
  and (_20058_, _20057_, _06239_);
  or (_20059_, _20058_, _20055_);
  and (_20060_, _20059_, _06220_);
  and (_20061_, _20048_, _06219_);
  or (_20063_, _20061_, _09818_);
  or (_20064_, _20063_, _20060_);
  or (_20065_, _20057_, _09827_);
  and (_20066_, _20065_, _05669_);
  and (_20067_, _20066_, _20064_);
  and (_20068_, _20067_, _20043_);
  and (_20069_, _14778_, _07653_);
  or (_20070_, _20069_, _20033_);
  and (_20071_, _20070_, _09833_);
  or (_20072_, _20071_, _06019_);
  or (_20074_, _20072_, _20068_);
  and (_20075_, _20074_, _20039_);
  or (_20076_, _20075_, _06112_);
  and (_20077_, _14793_, _07653_);
  or (_20078_, _20033_, _08751_);
  or (_20079_, _20078_, _20077_);
  and (_20080_, _20079_, _08756_);
  and (_20081_, _20080_, _20076_);
  and (_20082_, _12299_, _07653_);
  or (_20083_, _20082_, _20033_);
  and (_20085_, _20083_, _06284_);
  or (_20086_, _20085_, _20081_);
  and (_20087_, _20086_, _07032_);
  or (_20088_, _20087_, _20038_);
  and (_20089_, _20088_, _06278_);
  and (_20090_, _20048_, _06277_);
  and (_20091_, _20090_, _20034_);
  or (_20092_, _20091_, _06130_);
  or (_20093_, _20092_, _20089_);
  and (_20094_, _14792_, _07653_);
  or (_20096_, _20033_, _08777_);
  or (_20097_, _20096_, _20094_);
  and (_20098_, _20097_, _08782_);
  and (_20099_, _20098_, _20093_);
  nor (_20100_, _10988_, _11185_);
  or (_20101_, _20100_, _20033_);
  and (_20102_, _20101_, _06292_);
  or (_20103_, _20102_, _20099_);
  and (_20104_, _20103_, _06718_);
  and (_20105_, _20045_, _06316_);
  or (_20107_, _20105_, _06047_);
  or (_20108_, _20107_, _20104_);
  and (_20109_, _14849_, _07653_);
  or (_20110_, _20033_, _06048_);
  or (_20111_, _20110_, _20109_);
  and (_20112_, _20111_, _01336_);
  and (_20113_, _20112_, _20108_);
  or (_20114_, _20113_, _20032_);
  and (_43352_, _20114_, _42882_);
  and (_20115_, _01340_, \oc8051_golden_model_1.TMOD [4]);
  and (_20117_, _11185_, \oc8051_golden_model_1.TMOD [4]);
  and (_20118_, _08665_, _07653_);
  or (_20119_, _20118_, _20117_);
  or (_20120_, _20119_, _06020_);
  and (_20121_, _14887_, _07653_);
  or (_20122_, _20121_, _20117_);
  or (_20123_, _20122_, _06954_);
  and (_20124_, _07653_, \oc8051_golden_model_1.ACC [4]);
  or (_20125_, _20124_, _20117_);
  and (_20126_, _20125_, _06938_);
  and (_20128_, _06939_, \oc8051_golden_model_1.TMOD [4]);
  or (_20129_, _20128_, _06102_);
  or (_20130_, _20129_, _20126_);
  and (_20131_, _20130_, _06848_);
  and (_20132_, _20131_, _20123_);
  nor (_20133_, _08270_, _11185_);
  or (_20134_, _20133_, _20117_);
  and (_20135_, _20134_, _06239_);
  or (_20136_, _20135_, _20132_);
  and (_20137_, _20136_, _06220_);
  and (_20139_, _20125_, _06219_);
  or (_20140_, _20139_, _09818_);
  or (_20141_, _20140_, _20137_);
  and (_20142_, _09180_, _07653_);
  or (_20143_, _20117_, _07012_);
  or (_20144_, _20143_, _20142_);
  or (_20145_, _20134_, _09827_);
  and (_20146_, _20145_, _05669_);
  and (_20147_, _20146_, _20144_);
  and (_20148_, _20147_, _20141_);
  and (_20150_, _14983_, _07653_);
  or (_20151_, _20150_, _20117_);
  and (_20152_, _20151_, _09833_);
  or (_20153_, _20152_, _06019_);
  or (_20154_, _20153_, _20148_);
  and (_20155_, _20154_, _20120_);
  or (_20156_, _20155_, _06112_);
  and (_20157_, _14876_, _07653_);
  or (_20158_, _20117_, _08751_);
  or (_20159_, _20158_, _20157_);
  and (_20161_, _20159_, _08756_);
  and (_20162_, _20161_, _20156_);
  and (_20163_, _10986_, _07653_);
  or (_20164_, _20163_, _20117_);
  and (_20165_, _20164_, _06284_);
  or (_20166_, _20165_, _20162_);
  and (_20167_, _20166_, _07032_);
  or (_20168_, _20117_, _08273_);
  and (_20169_, _20119_, _06108_);
  and (_20170_, _20169_, _20168_);
  or (_20172_, _20170_, _20167_);
  and (_20173_, _20172_, _06278_);
  and (_20174_, _20125_, _06277_);
  and (_20175_, _20174_, _20168_);
  or (_20176_, _20175_, _06130_);
  or (_20177_, _20176_, _20173_);
  and (_20178_, _14873_, _07653_);
  or (_20179_, _20117_, _08777_);
  or (_20180_, _20179_, _20178_);
  and (_20181_, _20180_, _08782_);
  and (_20183_, _20181_, _20177_);
  nor (_20184_, _10985_, _11185_);
  or (_20185_, _20184_, _20117_);
  and (_20186_, _20185_, _06292_);
  or (_20187_, _20186_, _20183_);
  and (_20188_, _20187_, _06718_);
  and (_20189_, _20122_, _06316_);
  or (_20190_, _20189_, _06047_);
  or (_20191_, _20190_, _20188_);
  and (_20192_, _15055_, _07653_);
  or (_20194_, _20117_, _06048_);
  or (_20195_, _20194_, _20192_);
  and (_20196_, _20195_, _01336_);
  and (_20197_, _20196_, _20191_);
  or (_20198_, _20197_, _20115_);
  and (_43353_, _20198_, _42882_);
  and (_20199_, _01340_, \oc8051_golden_model_1.TMOD [5]);
  and (_20200_, _11185_, \oc8051_golden_model_1.TMOD [5]);
  or (_20201_, _20200_, _07980_);
  and (_20202_, _08652_, _07653_);
  or (_20204_, _20202_, _20200_);
  and (_20205_, _20204_, _06108_);
  and (_20206_, _20205_, _20201_);
  or (_20207_, _20204_, _06020_);
  and (_20208_, _15093_, _07653_);
  or (_20209_, _20208_, _20200_);
  or (_20210_, _20209_, _06954_);
  and (_20211_, _07653_, \oc8051_golden_model_1.ACC [5]);
  or (_20212_, _20211_, _20200_);
  and (_20213_, _20212_, _06938_);
  and (_20215_, _06939_, \oc8051_golden_model_1.TMOD [5]);
  or (_20216_, _20215_, _06102_);
  or (_20217_, _20216_, _20213_);
  and (_20218_, _20217_, _06848_);
  and (_20219_, _20218_, _20210_);
  nor (_20220_, _07977_, _11185_);
  or (_20221_, _20220_, _20200_);
  and (_20222_, _20221_, _06239_);
  or (_20223_, _20222_, _20219_);
  and (_20224_, _20223_, _06220_);
  and (_20226_, _20212_, _06219_);
  or (_20227_, _20226_, _09818_);
  or (_20228_, _20227_, _20224_);
  and (_20229_, _09179_, _07653_);
  or (_20230_, _20200_, _07012_);
  or (_20231_, _20230_, _20229_);
  or (_20232_, _20221_, _09827_);
  and (_20233_, _20232_, _05669_);
  and (_20234_, _20233_, _20231_);
  and (_20235_, _20234_, _20228_);
  and (_20237_, _15179_, _07653_);
  or (_20238_, _20237_, _20200_);
  and (_20239_, _20238_, _09833_);
  or (_20240_, _20239_, _06019_);
  or (_20241_, _20240_, _20235_);
  and (_20242_, _20241_, _20207_);
  or (_20243_, _20242_, _06112_);
  and (_20244_, _15195_, _07653_);
  or (_20245_, _20244_, _20200_);
  or (_20246_, _20245_, _08751_);
  and (_20248_, _20246_, _08756_);
  and (_20249_, _20248_, _20243_);
  and (_20250_, _12306_, _07653_);
  or (_20251_, _20250_, _20200_);
  and (_20252_, _20251_, _06284_);
  or (_20253_, _20252_, _20249_);
  and (_20254_, _20253_, _07032_);
  or (_20255_, _20254_, _20206_);
  and (_20256_, _20255_, _06278_);
  and (_20257_, _20212_, _06277_);
  and (_20259_, _20257_, _20201_);
  or (_20260_, _20259_, _06130_);
  or (_20261_, _20260_, _20256_);
  and (_20262_, _15194_, _07653_);
  or (_20263_, _20200_, _08777_);
  or (_20264_, _20263_, _20262_);
  and (_20265_, _20264_, _08782_);
  and (_20266_, _20265_, _20261_);
  nor (_20267_, _10982_, _11185_);
  or (_20268_, _20267_, _20200_);
  and (_20270_, _20268_, _06292_);
  or (_20271_, _20270_, _20266_);
  and (_20272_, _20271_, _06718_);
  and (_20273_, _20209_, _06316_);
  or (_20274_, _20273_, _06047_);
  or (_20275_, _20274_, _20272_);
  and (_20276_, _15253_, _07653_);
  or (_20277_, _20200_, _06048_);
  or (_20278_, _20277_, _20276_);
  and (_20279_, _20278_, _01336_);
  and (_20281_, _20279_, _20275_);
  or (_20282_, _20281_, _20199_);
  and (_43354_, _20282_, _42882_);
  and (_20283_, _01340_, \oc8051_golden_model_1.TMOD [6]);
  and (_20284_, _11185_, \oc8051_golden_model_1.TMOD [6]);
  or (_20285_, _20284_, _07886_);
  and (_20286_, _15389_, _07653_);
  or (_20287_, _20286_, _20284_);
  and (_20288_, _20287_, _06108_);
  and (_20289_, _20288_, _20285_);
  or (_20291_, _20287_, _06020_);
  and (_20292_, _15293_, _07653_);
  or (_20293_, _20292_, _20284_);
  or (_20294_, _20293_, _06954_);
  and (_20295_, _07653_, \oc8051_golden_model_1.ACC [6]);
  or (_20296_, _20295_, _20284_);
  and (_20297_, _20296_, _06938_);
  and (_20298_, _06939_, \oc8051_golden_model_1.TMOD [6]);
  or (_20299_, _20298_, _06102_);
  or (_20300_, _20299_, _20297_);
  and (_20302_, _20300_, _06848_);
  and (_20303_, _20302_, _20294_);
  nor (_20304_, _07883_, _11185_);
  or (_20305_, _20304_, _20284_);
  and (_20306_, _20305_, _06239_);
  or (_20307_, _20306_, _20303_);
  and (_20308_, _20307_, _06220_);
  and (_20309_, _20296_, _06219_);
  or (_20310_, _20309_, _09818_);
  or (_20311_, _20310_, _20308_);
  and (_20313_, _09178_, _07653_);
  or (_20314_, _20284_, _07012_);
  or (_20315_, _20314_, _20313_);
  or (_20316_, _20305_, _09827_);
  and (_20317_, _20316_, _05669_);
  and (_20318_, _20317_, _20315_);
  and (_20319_, _20318_, _20311_);
  and (_20320_, _15382_, _07653_);
  or (_20321_, _20320_, _20284_);
  and (_20322_, _20321_, _09833_);
  or (_20324_, _20322_, _06019_);
  or (_20325_, _20324_, _20319_);
  and (_20326_, _20325_, _20291_);
  or (_20327_, _20326_, _06112_);
  and (_20328_, _15399_, _07653_);
  or (_20329_, _20328_, _20284_);
  or (_20330_, _20329_, _08751_);
  and (_20331_, _20330_, _08756_);
  and (_20332_, _20331_, _20327_);
  and (_20333_, _10980_, _07653_);
  or (_20335_, _20333_, _20284_);
  and (_20336_, _20335_, _06284_);
  or (_20337_, _20336_, _20332_);
  and (_20338_, _20337_, _07032_);
  or (_20339_, _20338_, _20289_);
  and (_20340_, _20339_, _06278_);
  and (_20341_, _20296_, _06277_);
  and (_20342_, _20341_, _20285_);
  or (_20343_, _20342_, _06130_);
  or (_20344_, _20343_, _20340_);
  and (_20346_, _15396_, _07653_);
  or (_20347_, _20284_, _08777_);
  or (_20348_, _20347_, _20346_);
  and (_20349_, _20348_, _08782_);
  and (_20350_, _20349_, _20344_);
  nor (_20351_, _10979_, _11185_);
  or (_20352_, _20351_, _20284_);
  and (_20353_, _20352_, _06292_);
  or (_20354_, _20353_, _20350_);
  and (_20355_, _20354_, _06718_);
  and (_20357_, _20293_, _06316_);
  or (_20358_, _20357_, _06047_);
  or (_20359_, _20358_, _20355_);
  and (_20360_, _15451_, _07653_);
  or (_20361_, _20284_, _06048_);
  or (_20362_, _20361_, _20360_);
  and (_20363_, _20362_, _01336_);
  and (_20364_, _20363_, _20359_);
  or (_20365_, _20364_, _20283_);
  and (_43355_, _20365_, _42882_);
  not (_20367_, \oc8051_golden_model_1.DPL [0]);
  nor (_20368_, _01336_, _20367_);
  nand (_20369_, _10995_, _07733_);
  nor (_20370_, _07733_, _20367_);
  nor (_20371_, _20370_, _06278_);
  nand (_20372_, _20371_, _20369_);
  and (_20373_, _09120_, _07733_);
  or (_20374_, _20370_, _07012_);
  or (_20375_, _20374_, _20373_);
  and (_20376_, _07733_, _06931_);
  nor (_20378_, _20376_, _20370_);
  nand (_20379_, _20378_, _09815_);
  and (_20380_, _07733_, \oc8051_golden_model_1.ACC [0]);
  nor (_20381_, _20380_, _20370_);
  and (_20382_, _20381_, _06219_);
  nor (_20383_, _08127_, _11264_);
  or (_20384_, _20383_, _20370_);
  or (_20385_, _20384_, _06954_);
  nor (_20386_, _20381_, _06939_);
  nor (_20387_, _06938_, _20367_);
  or (_20389_, _20387_, _06102_);
  or (_20390_, _20389_, _20386_);
  and (_20391_, _20390_, _06848_);
  nand (_20392_, _20391_, _20385_);
  or (_20393_, _20378_, _06848_);
  and (_20394_, _20393_, _06220_);
  and (_20395_, _20394_, _20392_);
  or (_20396_, _20395_, _20382_);
  and (_20397_, _20396_, _11291_);
  and (_20398_, _11290_, \oc8051_golden_model_1.DPL [0]);
  or (_20400_, _20398_, _06110_);
  or (_20401_, _20400_, _20397_);
  or (_20402_, _06633_, _06111_);
  and (_20403_, _20402_, _09817_);
  nand (_20404_, _20403_, _20401_);
  and (_20405_, _20404_, _20379_);
  and (_20406_, _20405_, _20375_);
  or (_20407_, _20406_, _09833_);
  and (_20408_, _14186_, _07733_);
  or (_20409_, _20370_, _05669_);
  or (_20411_, _20409_, _20408_);
  and (_20412_, _20411_, _06020_);
  and (_20413_, _20412_, _20407_);
  and (_20414_, _07733_, _08672_);
  or (_20415_, _20414_, _20370_);
  and (_20416_, _20415_, _06019_);
  or (_20417_, _20416_, _06112_);
  or (_20418_, _20417_, _20413_);
  and (_20419_, _14086_, _07733_);
  or (_20420_, _20370_, _08751_);
  or (_20422_, _20420_, _20419_);
  and (_20423_, _20422_, _08756_);
  and (_20424_, _20423_, _20418_);
  nor (_20425_, _12302_, _11264_);
  or (_20426_, _20425_, _20370_);
  and (_20427_, _20369_, _06284_);
  and (_20428_, _20427_, _20426_);
  or (_20429_, _20428_, _20424_);
  and (_20430_, _20429_, _07032_);
  nand (_20431_, _20415_, _06108_);
  nor (_20433_, _20431_, _20383_);
  or (_20434_, _20433_, _06277_);
  or (_20435_, _20434_, _20430_);
  and (_20436_, _20435_, _20372_);
  or (_20437_, _20436_, _06130_);
  and (_20438_, _14083_, _07733_);
  or (_20439_, _20370_, _08777_);
  or (_20440_, _20439_, _20438_);
  and (_20441_, _20440_, _08782_);
  and (_20442_, _20441_, _20437_);
  and (_20444_, _20426_, _06292_);
  or (_20445_, _20444_, _19256_);
  or (_20446_, _20445_, _20442_);
  or (_20447_, _20384_, _06408_);
  and (_20448_, _20447_, _01336_);
  and (_20449_, _20448_, _20446_);
  or (_20450_, _20449_, _20368_);
  and (_43357_, _20450_, _42882_);
  not (_20451_, \oc8051_golden_model_1.DPL [1]);
  nor (_20452_, _01336_, _20451_);
  and (_20454_, _09075_, _07733_);
  nor (_20455_, _07733_, _20451_);
  or (_20456_, _20455_, _07012_);
  or (_20457_, _20456_, _20454_);
  or (_20458_, _07733_, \oc8051_golden_model_1.DPL [1]);
  and (_20459_, _14284_, _07733_);
  not (_20460_, _20459_);
  and (_20461_, _20460_, _20458_);
  or (_20462_, _20461_, _06954_);
  and (_20463_, _07733_, \oc8051_golden_model_1.ACC [1]);
  or (_20465_, _20463_, _20455_);
  and (_20466_, _20465_, _06938_);
  nor (_20467_, _06938_, _20451_);
  or (_20468_, _20467_, _06102_);
  or (_20469_, _20468_, _20466_);
  and (_20470_, _20469_, _06848_);
  and (_20471_, _20470_, _20462_);
  nor (_20472_, _11264_, _07132_);
  or (_20473_, _20472_, _20455_);
  and (_20474_, _20473_, _06239_);
  or (_20476_, _20474_, _06219_);
  or (_20477_, _20476_, _20471_);
  or (_20478_, _20465_, _06220_);
  and (_20479_, _20478_, _11291_);
  and (_20480_, _20479_, _20477_);
  nor (_20481_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_20482_, _20481_, _11295_);
  and (_20483_, _20482_, _11290_);
  or (_20484_, _20483_, _20480_);
  and (_20485_, _20484_, _06111_);
  nor (_20487_, _06832_, _06111_);
  or (_20488_, _20487_, _09818_);
  or (_20489_, _20488_, _20485_);
  or (_20490_, _20473_, _09827_);
  and (_20491_, _20490_, _05669_);
  and (_20492_, _20491_, _20489_);
  and (_20493_, _20492_, _20457_);
  or (_20494_, _14367_, _11264_);
  and (_20495_, _20458_, _09833_);
  and (_20496_, _20495_, _20494_);
  or (_20498_, _20496_, _20493_);
  and (_20499_, _20498_, _06020_);
  nand (_20500_, _07733_, _06832_);
  and (_20501_, _20458_, _06019_);
  and (_20502_, _20501_, _20500_);
  or (_20503_, _20502_, _20499_);
  and (_20504_, _20503_, _08751_);
  or (_20505_, _14263_, _11264_);
  and (_20506_, _20458_, _06112_);
  and (_20507_, _20506_, _20505_);
  or (_20509_, _20507_, _06284_);
  or (_20510_, _20509_, _20504_);
  nor (_20511_, _10993_, _11264_);
  or (_20512_, _20511_, _20455_);
  nand (_20513_, _10992_, _07733_);
  and (_20514_, _20513_, _20512_);
  or (_20515_, _20514_, _08756_);
  and (_20516_, _20515_, _07032_);
  and (_20517_, _20516_, _20510_);
  or (_20518_, _14261_, _11264_);
  and (_20520_, _20458_, _06108_);
  and (_20521_, _20520_, _20518_);
  or (_20522_, _20521_, _06277_);
  or (_20523_, _20522_, _20517_);
  nor (_20524_, _20455_, _06278_);
  nand (_20525_, _20524_, _20513_);
  and (_20526_, _20525_, _08777_);
  and (_20527_, _20526_, _20523_);
  or (_20528_, _20500_, _08078_);
  and (_20529_, _20458_, _06130_);
  and (_20531_, _20529_, _20528_);
  or (_20532_, _20531_, _06292_);
  or (_20533_, _20532_, _20527_);
  or (_20534_, _20512_, _08782_);
  and (_20535_, _20534_, _06718_);
  and (_20536_, _20535_, _20533_);
  and (_20537_, _20461_, _06316_);
  or (_20538_, _20537_, _06047_);
  or (_20539_, _20538_, _20536_);
  or (_20540_, _20455_, _06048_);
  or (_20542_, _20540_, _20459_);
  and (_20543_, _20542_, _01336_);
  and (_20544_, _20543_, _20539_);
  or (_20545_, _20544_, _20452_);
  and (_43358_, _20545_, _42882_);
  not (_20546_, \oc8051_golden_model_1.DPL [2]);
  nor (_20547_, _01336_, _20546_);
  nor (_20548_, _07733_, _20546_);
  or (_20549_, _20548_, _08177_);
  and (_20550_, _07733_, _08730_);
  or (_20552_, _20550_, _20548_);
  and (_20553_, _20552_, _06108_);
  and (_20554_, _20553_, _20549_);
  or (_20555_, _20552_, _06020_);
  and (_20556_, _14493_, _07733_);
  or (_20557_, _20556_, _20548_);
  or (_20558_, _20557_, _06954_);
  and (_20559_, _07733_, \oc8051_golden_model_1.ACC [2]);
  or (_20560_, _20559_, _20548_);
  and (_20561_, _20560_, _06938_);
  nor (_20563_, _06938_, _20546_);
  or (_20564_, _20563_, _06102_);
  or (_20565_, _20564_, _20561_);
  and (_20566_, _20565_, _06848_);
  and (_20567_, _20566_, _20558_);
  nor (_20568_, _11264_, _07530_);
  or (_20569_, _20568_, _20548_);
  and (_20570_, _20569_, _06239_);
  or (_20571_, _20570_, _06219_);
  or (_20572_, _20571_, _20567_);
  or (_20574_, _20560_, _06220_);
  and (_20575_, _20574_, _11291_);
  and (_20576_, _20575_, _20572_);
  nor (_20577_, _11295_, \oc8051_golden_model_1.DPL [2]);
  nor (_20578_, _20577_, _11296_);
  and (_20579_, _20578_, _11290_);
  or (_20580_, _20579_, _20576_);
  and (_20581_, _20580_, _06111_);
  nor (_20582_, _06445_, _06111_);
  or (_20583_, _20582_, _09818_);
  or (_20585_, _20583_, _20581_);
  and (_20586_, _09182_, _07733_);
  or (_20587_, _20548_, _07012_);
  or (_20588_, _20587_, _20586_);
  or (_20589_, _20569_, _09827_);
  and (_20590_, _20589_, _05669_);
  and (_20591_, _20590_, _20588_);
  and (_20592_, _20591_, _20585_);
  and (_20593_, _14580_, _07733_);
  or (_20594_, _20593_, _20548_);
  and (_20596_, _20594_, _09833_);
  or (_20597_, _20596_, _06019_);
  or (_20598_, _20597_, _20592_);
  and (_20599_, _20598_, _20555_);
  or (_20600_, _20599_, _06112_);
  and (_20601_, _14596_, _07733_);
  or (_20602_, _20601_, _20548_);
  or (_20603_, _20602_, _08751_);
  and (_20604_, _20603_, _08756_);
  and (_20605_, _20604_, _20600_);
  and (_20607_, _10991_, _07733_);
  or (_20608_, _20607_, _20548_);
  and (_20609_, _20608_, _06284_);
  or (_20610_, _20609_, _20605_);
  and (_20611_, _20610_, _07032_);
  or (_20612_, _20611_, _20554_);
  and (_20613_, _20612_, _06278_);
  and (_20614_, _20560_, _06277_);
  and (_20615_, _20614_, _20549_);
  or (_20616_, _20615_, _06130_);
  or (_20618_, _20616_, _20613_);
  and (_20619_, _14593_, _07733_);
  or (_20620_, _20548_, _08777_);
  or (_20621_, _20620_, _20619_);
  and (_20622_, _20621_, _08782_);
  and (_20623_, _20622_, _20618_);
  nor (_20624_, _10990_, _11264_);
  or (_20625_, _20624_, _20548_);
  and (_20626_, _20625_, _06292_);
  or (_20627_, _20626_, _20623_);
  and (_20629_, _20627_, _06718_);
  and (_20630_, _20557_, _06316_);
  or (_20631_, _20630_, _06047_);
  or (_20632_, _20631_, _20629_);
  and (_20633_, _14657_, _07733_);
  or (_20634_, _20548_, _06048_);
  or (_20635_, _20634_, _20633_);
  and (_20636_, _20635_, _01336_);
  and (_20637_, _20636_, _20632_);
  or (_20638_, _20637_, _20547_);
  and (_43359_, _20638_, _42882_);
  not (_20640_, \oc8051_golden_model_1.DPL [3]);
  nor (_20641_, _01336_, _20640_);
  nor (_20642_, _07733_, _20640_);
  or (_20643_, _20642_, _08029_);
  and (_20644_, _07733_, _08662_);
  or (_20645_, _20644_, _20642_);
  and (_20646_, _20645_, _06108_);
  and (_20647_, _20646_, _20643_);
  or (_20648_, _20645_, _06020_);
  and (_20650_, _14672_, _07733_);
  or (_20651_, _20650_, _20642_);
  or (_20652_, _20651_, _06954_);
  and (_20653_, _07733_, \oc8051_golden_model_1.ACC [3]);
  or (_20654_, _20653_, _20642_);
  and (_20655_, _20654_, _06938_);
  nor (_20656_, _06938_, _20640_);
  or (_20657_, _20656_, _06102_);
  or (_20658_, _20657_, _20655_);
  and (_20659_, _20658_, _06848_);
  and (_20661_, _20659_, _20652_);
  nor (_20662_, _11264_, _07353_);
  or (_20663_, _20662_, _20642_);
  and (_20664_, _20663_, _06239_);
  or (_20665_, _20664_, _06219_);
  or (_20666_, _20665_, _20661_);
  or (_20667_, _20654_, _06220_);
  and (_20668_, _20667_, _11291_);
  and (_20669_, _20668_, _20666_);
  nor (_20670_, _11296_, \oc8051_golden_model_1.DPL [3]);
  nor (_20672_, _20670_, _11297_);
  and (_20673_, _20672_, _11290_);
  or (_20674_, _20673_, _20669_);
  and (_20675_, _20674_, _06111_);
  nor (_20676_, _06215_, _06111_);
  or (_20677_, _20676_, _09818_);
  or (_20678_, _20677_, _20675_);
  and (_20679_, _09181_, _07733_);
  or (_20680_, _20642_, _07012_);
  or (_20681_, _20680_, _20679_);
  or (_20683_, _20663_, _09827_);
  and (_20684_, _20683_, _05669_);
  and (_20685_, _20684_, _20681_);
  and (_20686_, _20685_, _20678_);
  and (_20687_, _14778_, _07733_);
  or (_20688_, _20687_, _20642_);
  and (_20689_, _20688_, _09833_);
  or (_20690_, _20689_, _06019_);
  or (_20691_, _20690_, _20686_);
  and (_20692_, _20691_, _20648_);
  or (_20694_, _20692_, _06112_);
  and (_20695_, _14793_, _07733_);
  or (_20696_, _20642_, _08751_);
  or (_20697_, _20696_, _20695_);
  and (_20698_, _20697_, _08756_);
  and (_20699_, _20698_, _20694_);
  and (_20700_, _12299_, _07733_);
  or (_20701_, _20700_, _20642_);
  and (_20702_, _20701_, _06284_);
  or (_20703_, _20702_, _20699_);
  and (_20705_, _20703_, _07032_);
  or (_20706_, _20705_, _20647_);
  and (_20707_, _20706_, _06278_);
  and (_20708_, _20654_, _06277_);
  and (_20709_, _20708_, _20643_);
  or (_20710_, _20709_, _06130_);
  or (_20711_, _20710_, _20707_);
  and (_20712_, _14792_, _07733_);
  or (_20713_, _20642_, _08777_);
  or (_20714_, _20713_, _20712_);
  and (_20716_, _20714_, _08782_);
  and (_20717_, _20716_, _20711_);
  nor (_20718_, _10988_, _11264_);
  or (_20719_, _20718_, _20642_);
  and (_20720_, _20719_, _06292_);
  or (_20721_, _20720_, _20717_);
  and (_20722_, _20721_, _06718_);
  and (_20723_, _20651_, _06316_);
  or (_20724_, _20723_, _06047_);
  or (_20725_, _20724_, _20722_);
  and (_20727_, _14849_, _07733_);
  or (_20728_, _20642_, _06048_);
  or (_20729_, _20728_, _20727_);
  and (_20730_, _20729_, _01336_);
  and (_20731_, _20730_, _20725_);
  or (_20732_, _20731_, _20641_);
  and (_43361_, _20732_, _42882_);
  not (_20733_, \oc8051_golden_model_1.DPL [4]);
  nor (_20734_, _01336_, _20733_);
  nor (_20735_, _07733_, _20733_);
  or (_20737_, _20735_, _08273_);
  and (_20738_, _08665_, _07733_);
  or (_20739_, _20738_, _20735_);
  and (_20740_, _20739_, _06108_);
  and (_20741_, _20740_, _20737_);
  or (_20742_, _20739_, _06020_);
  and (_20743_, _14887_, _07733_);
  or (_20744_, _20743_, _20735_);
  or (_20745_, _20744_, _06954_);
  and (_20746_, _07733_, \oc8051_golden_model_1.ACC [4]);
  or (_20748_, _20746_, _20735_);
  and (_20749_, _20748_, _06938_);
  nor (_20750_, _06938_, _20733_);
  or (_20751_, _20750_, _06102_);
  or (_20752_, _20751_, _20749_);
  and (_20753_, _20752_, _06848_);
  and (_20754_, _20753_, _20745_);
  nor (_20755_, _08270_, _11264_);
  or (_20756_, _20755_, _20735_);
  and (_20757_, _20756_, _06239_);
  or (_20758_, _20757_, _06219_);
  or (_20759_, _20758_, _20754_);
  or (_20760_, _20748_, _06220_);
  and (_20761_, _20760_, _11291_);
  and (_20762_, _20761_, _20759_);
  nor (_20763_, _11297_, \oc8051_golden_model_1.DPL [4]);
  nor (_20764_, _20763_, _11298_);
  and (_20765_, _20764_, _11290_);
  or (_20766_, _20765_, _20762_);
  and (_20767_, _20766_, _06111_);
  nor (_20769_, _08581_, _06111_);
  or (_20770_, _20769_, _09818_);
  or (_20771_, _20770_, _20767_);
  and (_20772_, _09180_, _07733_);
  or (_20773_, _20735_, _07012_);
  or (_20774_, _20773_, _20772_);
  or (_20775_, _20756_, _09827_);
  and (_20776_, _20775_, _05669_);
  and (_20777_, _20776_, _20774_);
  and (_20778_, _20777_, _20771_);
  and (_20781_, _14983_, _07733_);
  or (_20782_, _20781_, _20735_);
  and (_20783_, _20782_, _09833_);
  or (_20784_, _20783_, _06019_);
  or (_20785_, _20784_, _20778_);
  and (_20786_, _20785_, _20742_);
  or (_20787_, _20786_, _06112_);
  and (_20788_, _14876_, _07733_);
  or (_20789_, _20788_, _20735_);
  or (_20790_, _20789_, _08751_);
  and (_20792_, _20790_, _08756_);
  and (_20793_, _20792_, _20787_);
  and (_20794_, _10986_, _07733_);
  or (_20795_, _20794_, _20735_);
  and (_20796_, _20795_, _06284_);
  or (_20797_, _20796_, _20793_);
  and (_20798_, _20797_, _07032_);
  or (_20799_, _20798_, _20741_);
  and (_20800_, _20799_, _06278_);
  and (_20801_, _20748_, _06277_);
  and (_20802_, _20801_, _20737_);
  or (_20803_, _20802_, _06130_);
  or (_20804_, _20803_, _20800_);
  and (_20805_, _14873_, _07733_);
  or (_20806_, _20735_, _08777_);
  or (_20807_, _20806_, _20805_);
  and (_20808_, _20807_, _08782_);
  and (_20809_, _20808_, _20804_);
  nor (_20810_, _10985_, _11264_);
  or (_20811_, _20810_, _20735_);
  and (_20813_, _20811_, _06292_);
  or (_20814_, _20813_, _20809_);
  and (_20815_, _20814_, _06718_);
  and (_20816_, _20744_, _06316_);
  or (_20817_, _20816_, _06047_);
  or (_20818_, _20817_, _20815_);
  and (_20819_, _15055_, _07733_);
  or (_20820_, _20735_, _06048_);
  or (_20821_, _20820_, _20819_);
  and (_20822_, _20821_, _01336_);
  and (_20825_, _20822_, _20818_);
  or (_20826_, _20825_, _20734_);
  and (_43362_, _20826_, _42882_);
  not (_20827_, \oc8051_golden_model_1.DPL [5]);
  nor (_20828_, _01336_, _20827_);
  nor (_20829_, _07733_, _20827_);
  and (_20830_, _08652_, _07733_);
  or (_20831_, _20830_, _20829_);
  or (_20832_, _20831_, _06020_);
  and (_20833_, _15093_, _07733_);
  or (_20834_, _20833_, _20829_);
  or (_20835_, _20834_, _06954_);
  and (_20836_, _07733_, \oc8051_golden_model_1.ACC [5]);
  or (_20837_, _20836_, _20829_);
  and (_20838_, _20837_, _06938_);
  nor (_20839_, _06938_, _20827_);
  or (_20840_, _20839_, _06102_);
  or (_20841_, _20840_, _20838_);
  and (_20842_, _20841_, _06848_);
  and (_20843_, _20842_, _20835_);
  nor (_20845_, _07977_, _11264_);
  or (_20846_, _20845_, _20829_);
  and (_20847_, _20846_, _06239_);
  or (_20848_, _20847_, _06219_);
  or (_20849_, _20848_, _20843_);
  or (_20850_, _20837_, _06220_);
  and (_20851_, _20850_, _11291_);
  and (_20852_, _20851_, _20849_);
  nor (_20853_, _11298_, \oc8051_golden_model_1.DPL [5]);
  nor (_20854_, _20853_, _11299_);
  and (_20857_, _20854_, _11290_);
  or (_20858_, _20857_, _20852_);
  and (_20859_, _20858_, _06111_);
  nor (_20860_, _08612_, _06111_);
  or (_20861_, _20860_, _09818_);
  or (_20862_, _20861_, _20859_);
  and (_20863_, _09179_, _07733_);
  or (_20864_, _20829_, _07012_);
  or (_20865_, _20864_, _20863_);
  or (_20866_, _20846_, _09827_);
  and (_20868_, _20866_, _05669_);
  and (_20869_, _20868_, _20865_);
  and (_20870_, _20869_, _20862_);
  and (_20871_, _15179_, _07733_);
  or (_20872_, _20871_, _20829_);
  and (_20873_, _20872_, _09833_);
  or (_20874_, _20873_, _06019_);
  or (_20875_, _20874_, _20870_);
  and (_20876_, _20875_, _20832_);
  or (_20877_, _20876_, _06112_);
  and (_20879_, _15195_, _07733_);
  or (_20880_, _20879_, _20829_);
  or (_20881_, _20880_, _08751_);
  and (_20882_, _20881_, _08756_);
  and (_20883_, _20882_, _20877_);
  and (_20884_, _12306_, _07733_);
  or (_20885_, _20884_, _20829_);
  and (_20886_, _20885_, _06284_);
  or (_20887_, _20886_, _20883_);
  and (_20888_, _20887_, _07032_);
  or (_20890_, _20829_, _07980_);
  and (_20891_, _20831_, _06108_);
  and (_20892_, _20891_, _20890_);
  or (_20893_, _20892_, _20888_);
  and (_20894_, _20893_, _06278_);
  and (_20895_, _20837_, _06277_);
  and (_20896_, _20895_, _20890_);
  or (_20897_, _20896_, _06130_);
  or (_20898_, _20897_, _20894_);
  and (_20899_, _15194_, _07733_);
  or (_20900_, _20829_, _08777_);
  or (_20901_, _20900_, _20899_);
  and (_20902_, _20901_, _08782_);
  and (_20903_, _20902_, _20898_);
  nor (_20904_, _10982_, _11264_);
  or (_20905_, _20904_, _20829_);
  and (_20906_, _20905_, _06292_);
  or (_20907_, _20906_, _20903_);
  and (_20908_, _20907_, _06718_);
  and (_20909_, _20834_, _06316_);
  or (_20912_, _20909_, _06047_);
  or (_20913_, _20912_, _20908_);
  and (_20914_, _15253_, _07733_);
  or (_20915_, _20829_, _06048_);
  or (_20916_, _20915_, _20914_);
  and (_20917_, _20916_, _01336_);
  and (_20918_, _20917_, _20913_);
  or (_20919_, _20918_, _20828_);
  and (_43363_, _20919_, _42882_);
  not (_20920_, \oc8051_golden_model_1.DPL [6]);
  nor (_20922_, _01336_, _20920_);
  nor (_20923_, _07733_, _20920_);
  and (_20924_, _15389_, _07733_);
  or (_20925_, _20924_, _20923_);
  or (_20926_, _20925_, _06020_);
  and (_20927_, _15293_, _07733_);
  or (_20928_, _20927_, _20923_);
  or (_20929_, _20928_, _06954_);
  and (_20930_, _07733_, \oc8051_golden_model_1.ACC [6]);
  or (_20931_, _20930_, _20923_);
  and (_20933_, _20931_, _06938_);
  nor (_20934_, _06938_, _20920_);
  or (_20935_, _20934_, _06102_);
  or (_20936_, _20935_, _20933_);
  and (_20937_, _20936_, _06848_);
  and (_20938_, _20937_, _20929_);
  nor (_20939_, _07883_, _11264_);
  or (_20940_, _20939_, _20923_);
  and (_20941_, _20940_, _06239_);
  or (_20942_, _20941_, _06219_);
  or (_20944_, _20942_, _20938_);
  or (_20945_, _20931_, _06220_);
  and (_20946_, _20945_, _11291_);
  and (_20947_, _20946_, _20944_);
  nor (_20948_, _11299_, \oc8051_golden_model_1.DPL [6]);
  nor (_20949_, _20948_, _11300_);
  and (_20950_, _20949_, _11290_);
  or (_20951_, _20950_, _20947_);
  and (_20952_, _20951_, _06111_);
  nor (_20953_, _08647_, _06111_);
  or (_20955_, _20953_, _09818_);
  or (_20956_, _20955_, _20952_);
  and (_20957_, _09178_, _07733_);
  or (_20958_, _20923_, _07012_);
  or (_20959_, _20958_, _20957_);
  or (_20960_, _20940_, _09827_);
  and (_20961_, _20960_, _05669_);
  and (_20962_, _20961_, _20959_);
  and (_20963_, _20962_, _20956_);
  and (_20964_, _15382_, _07733_);
  or (_20966_, _20964_, _20923_);
  and (_20967_, _20966_, _09833_);
  or (_20968_, _20967_, _06019_);
  or (_20969_, _20968_, _20963_);
  and (_20970_, _20969_, _20926_);
  or (_20971_, _20970_, _06112_);
  and (_20972_, _15399_, _07733_);
  or (_20973_, _20923_, _08751_);
  or (_20974_, _20973_, _20972_);
  and (_20975_, _20974_, _08756_);
  and (_20977_, _20975_, _20971_);
  and (_20978_, _10980_, _07733_);
  or (_20979_, _20978_, _20923_);
  and (_20980_, _20979_, _06284_);
  or (_20981_, _20980_, _20977_);
  and (_20982_, _20981_, _07032_);
  or (_20983_, _20923_, _07886_);
  and (_20984_, _20925_, _06108_);
  and (_20985_, _20984_, _20983_);
  or (_20986_, _20985_, _20982_);
  and (_20988_, _20986_, _06278_);
  and (_20989_, _20931_, _06277_);
  and (_20990_, _20989_, _20983_);
  or (_20991_, _20990_, _06130_);
  or (_20992_, _20991_, _20988_);
  and (_20993_, _15396_, _07733_);
  or (_20994_, _20923_, _08777_);
  or (_20995_, _20994_, _20993_);
  and (_20996_, _20995_, _08782_);
  and (_20997_, _20996_, _20992_);
  nor (_20999_, _10979_, _11264_);
  or (_21000_, _20999_, _20923_);
  and (_21001_, _21000_, _06292_);
  or (_21002_, _21001_, _20997_);
  and (_21003_, _21002_, _06718_);
  and (_21004_, _20928_, _06316_);
  or (_21005_, _21004_, _06047_);
  or (_21006_, _21005_, _21003_);
  and (_21007_, _15451_, _07733_);
  or (_21008_, _20923_, _06048_);
  or (_21010_, _21008_, _21007_);
  and (_21011_, _21010_, _01336_);
  and (_21012_, _21011_, _21006_);
  or (_21013_, _21012_, _20922_);
  and (_43364_, _21013_, _42882_);
  not (_21014_, \oc8051_golden_model_1.DPH [0]);
  nor (_21015_, _01336_, _21014_);
  nor (_21016_, _07802_, _21014_);
  and (_21017_, _07802_, \oc8051_golden_model_1.ACC [0]);
  and (_21018_, _21017_, _08127_);
  or (_21020_, _21018_, _21016_);
  or (_21021_, _21020_, _06278_);
  or (_21022_, _21016_, _07012_);
  and (_21023_, _09120_, _07802_);
  or (_21024_, _21023_, _21022_);
  and (_21025_, _07724_, _06931_);
  nor (_21026_, _21025_, _21016_);
  nand (_21027_, _21026_, _09815_);
  nor (_21028_, _08127_, _11359_);
  or (_21029_, _21028_, _21016_);
  or (_21030_, _21029_, _06954_);
  nor (_21031_, _21017_, _21016_);
  nor (_21032_, _21031_, _06939_);
  nor (_21033_, _06938_, _21014_);
  or (_21034_, _21033_, _06102_);
  or (_21035_, _21034_, _21032_);
  and (_21036_, _21035_, _06848_);
  nand (_21037_, _21036_, _21030_);
  or (_21038_, _21026_, _06848_);
  and (_21039_, _21038_, _06220_);
  and (_21042_, _21039_, _21037_);
  and (_21043_, _21031_, _06219_);
  or (_21044_, _21043_, _11290_);
  or (_21045_, _21044_, _21042_);
  nor (_21046_, _11302_, \oc8051_golden_model_1.DPH [0]);
  or (_21047_, _11388_, _11291_);
  or (_21048_, _21047_, _21046_);
  and (_21049_, _21048_, _21045_);
  or (_21050_, _21049_, _06110_);
  or (_21051_, _06111_, _06016_);
  and (_21053_, _21051_, _09817_);
  nand (_21054_, _21053_, _21050_);
  and (_21055_, _21054_, _21027_);
  and (_21056_, _21055_, _21024_);
  or (_21057_, _21056_, _09833_);
  and (_21058_, _14186_, _07724_);
  or (_21059_, _21016_, _05669_);
  or (_21060_, _21059_, _21058_);
  and (_21061_, _21060_, _06020_);
  and (_21062_, _21061_, _21057_);
  and (_21064_, _07802_, _08672_);
  or (_21065_, _21064_, _21016_);
  and (_21066_, _21065_, _06019_);
  or (_21067_, _21066_, _06112_);
  or (_21068_, _21067_, _21062_);
  and (_21069_, _14086_, _07724_);
  or (_21070_, _21016_, _08751_);
  or (_21071_, _21070_, _21069_);
  and (_21072_, _21071_, _08756_);
  and (_21073_, _21072_, _21068_);
  nor (_21075_, _12302_, _11359_);
  or (_21076_, _21075_, _21016_);
  nor (_21077_, _21018_, _08756_);
  and (_21078_, _21077_, _21076_);
  or (_21079_, _21078_, _21073_);
  and (_21080_, _21079_, _07032_);
  nand (_21081_, _21065_, _06108_);
  nor (_21082_, _21081_, _21028_);
  or (_21083_, _21082_, _06277_);
  or (_21084_, _21083_, _21080_);
  and (_21086_, _21084_, _21021_);
  or (_21087_, _21086_, _06130_);
  and (_21088_, _14083_, _07724_);
  or (_21089_, _21016_, _08777_);
  or (_21090_, _21089_, _21088_);
  and (_21091_, _21090_, _08782_);
  and (_21092_, _21091_, _21087_);
  and (_21093_, _21076_, _06292_);
  or (_21094_, _21093_, _19256_);
  or (_21095_, _21094_, _21092_);
  or (_21097_, _21029_, _06408_);
  and (_21098_, _21097_, _01336_);
  and (_21099_, _21098_, _21095_);
  or (_21100_, _21099_, _21015_);
  and (_43366_, _21100_, _42882_);
  not (_21101_, \oc8051_golden_model_1.DPH [1]);
  nor (_21102_, _01336_, _21101_);
  or (_21103_, _07802_, \oc8051_golden_model_1.DPH [1]);
  and (_21104_, _21103_, _09833_);
  or (_21105_, _14367_, _11359_);
  and (_21107_, _21105_, _21104_);
  nor (_21108_, _07802_, _21101_);
  nor (_21109_, _11359_, _07132_);
  or (_21110_, _21109_, _21108_);
  or (_21111_, _21110_, _06848_);
  and (_21112_, _14284_, _07724_);
  not (_21113_, _21112_);
  and (_21114_, _21113_, _21103_);
  and (_21115_, _21114_, _06102_);
  nor (_21116_, _06938_, _21101_);
  and (_21118_, _07802_, \oc8051_golden_model_1.ACC [1]);
  or (_21119_, _21118_, _21108_);
  and (_21120_, _21119_, _06938_);
  or (_21121_, _21120_, _21116_);
  and (_21122_, _21121_, _06954_);
  or (_21123_, _21122_, _06239_);
  or (_21124_, _21123_, _21115_);
  and (_21125_, _21124_, _21111_);
  or (_21126_, _21125_, _06219_);
  or (_21127_, _21119_, _06220_);
  and (_21129_, _21127_, _11291_);
  and (_21130_, _21129_, _21126_);
  or (_21131_, _11388_, \oc8051_golden_model_1.DPH [1]);
  nand (_21132_, _21131_, _11290_);
  nor (_21133_, _21132_, _11389_);
  or (_21134_, _21133_, _21130_);
  and (_21135_, _21134_, _06111_);
  nor (_21136_, _06799_, _06111_);
  or (_21137_, _21136_, _09818_);
  or (_21138_, _21137_, _21135_);
  or (_21140_, _21108_, _07012_);
  and (_21141_, _09075_, _07802_);
  or (_21142_, _21141_, _21140_);
  or (_21143_, _21110_, _09827_);
  and (_21144_, _21143_, _05669_);
  and (_21145_, _21144_, _21142_);
  and (_21146_, _21145_, _21138_);
  or (_21147_, _21146_, _21107_);
  and (_21148_, _21147_, _06020_);
  and (_21149_, _21103_, _06019_);
  nand (_21151_, _07724_, _06832_);
  and (_21152_, _21151_, _21149_);
  or (_21153_, _21152_, _21148_);
  and (_21154_, _21153_, _08751_);
  or (_21155_, _14263_, _11359_);
  and (_21156_, _21103_, _06112_);
  and (_21157_, _21156_, _21155_);
  or (_21158_, _21157_, _06284_);
  or (_21159_, _21158_, _21154_);
  nor (_21160_, _10993_, _11359_);
  or (_21162_, _21160_, _21108_);
  nand (_21163_, _10992_, _07724_);
  and (_21164_, _21163_, _21162_);
  or (_21165_, _21164_, _08756_);
  and (_21166_, _21165_, _07032_);
  and (_21167_, _21166_, _21159_);
  or (_21168_, _14261_, _11359_);
  and (_21169_, _21103_, _06108_);
  and (_21170_, _21169_, _21168_);
  or (_21171_, _21170_, _06277_);
  or (_21173_, _21171_, _21167_);
  nor (_21174_, _21108_, _06278_);
  nand (_21175_, _21174_, _21163_);
  and (_21176_, _21175_, _08777_);
  and (_21177_, _21176_, _21173_);
  or (_21178_, _21151_, _08078_);
  and (_21179_, _21103_, _06130_);
  and (_21180_, _21179_, _21178_);
  or (_21181_, _21180_, _06292_);
  or (_21182_, _21181_, _21177_);
  or (_21184_, _21162_, _08782_);
  and (_21185_, _21184_, _06718_);
  and (_21186_, _21185_, _21182_);
  and (_21187_, _21114_, _06316_);
  or (_21188_, _21187_, _06047_);
  or (_21189_, _21188_, _21186_);
  or (_21190_, _21108_, _06048_);
  or (_21191_, _21190_, _21112_);
  and (_21192_, _21191_, _01336_);
  and (_21193_, _21192_, _21189_);
  or (_21195_, _21193_, _21102_);
  and (_43367_, _21195_, _42882_);
  and (_21196_, _01340_, \oc8051_golden_model_1.DPH [2]);
  and (_21197_, _11359_, \oc8051_golden_model_1.DPH [2]);
  and (_21198_, _07802_, _08730_);
  or (_21199_, _21198_, _21197_);
  or (_21200_, _21199_, _06020_);
  and (_21201_, _14493_, _07724_);
  or (_21202_, _21201_, _21197_);
  or (_21203_, _21202_, _06954_);
  and (_21204_, _07802_, \oc8051_golden_model_1.ACC [2]);
  or (_21205_, _21204_, _21197_);
  and (_21206_, _21205_, _06938_);
  and (_21207_, _06939_, \oc8051_golden_model_1.DPH [2]);
  or (_21208_, _21207_, _06102_);
  or (_21209_, _21208_, _21206_);
  and (_21210_, _21209_, _06848_);
  and (_21211_, _21210_, _21203_);
  nor (_21212_, _11359_, _07530_);
  or (_21213_, _21212_, _21197_);
  and (_21216_, _21213_, _06239_);
  or (_21217_, _21216_, _06219_);
  or (_21218_, _21217_, _21211_);
  or (_21219_, _21205_, _06220_);
  and (_21220_, _21219_, _11291_);
  and (_21221_, _21220_, _21218_);
  or (_21222_, _11389_, \oc8051_golden_model_1.DPH [2]);
  nor (_21223_, _11390_, _11291_);
  and (_21224_, _21223_, _21222_);
  or (_21225_, _21224_, _21221_);
  and (_21227_, _21225_, _06111_);
  nor (_21228_, _06403_, _06111_);
  or (_21229_, _21228_, _09818_);
  or (_21230_, _21229_, _21227_);
  or (_21231_, _21197_, _07012_);
  and (_21232_, _09182_, _07802_);
  or (_21233_, _21232_, _21231_);
  or (_21234_, _21213_, _09827_);
  and (_21235_, _21234_, _05669_);
  and (_21236_, _21235_, _21233_);
  and (_21238_, _21236_, _21230_);
  and (_21239_, _14580_, _07724_);
  or (_21240_, _21239_, _21197_);
  and (_21241_, _21240_, _09833_);
  or (_21242_, _21241_, _06019_);
  or (_21243_, _21242_, _21238_);
  and (_21244_, _21243_, _21200_);
  or (_21245_, _21244_, _06112_);
  and (_21246_, _14596_, _07724_);
  or (_21247_, _21197_, _08751_);
  or (_21249_, _21247_, _21246_);
  and (_21250_, _21249_, _08756_);
  and (_21251_, _21250_, _21245_);
  and (_21252_, _10991_, _07802_);
  or (_21253_, _21252_, _21197_);
  and (_21254_, _21253_, _06284_);
  or (_21255_, _21254_, _21251_);
  and (_21256_, _21255_, _07032_);
  or (_21257_, _21197_, _08177_);
  and (_21258_, _21199_, _06108_);
  and (_21260_, _21258_, _21257_);
  or (_21261_, _21260_, _21256_);
  and (_21262_, _21261_, _06278_);
  and (_21263_, _21205_, _06277_);
  and (_21264_, _21263_, _21257_);
  or (_21265_, _21264_, _06130_);
  or (_21266_, _21265_, _21262_);
  and (_21267_, _14593_, _07724_);
  or (_21268_, _21197_, _08777_);
  or (_21269_, _21268_, _21267_);
  and (_21271_, _21269_, _08782_);
  and (_21272_, _21271_, _21266_);
  nor (_21273_, _10990_, _11359_);
  or (_21274_, _21273_, _21197_);
  and (_21275_, _21274_, _06292_);
  or (_21276_, _21275_, _21272_);
  and (_21277_, _21276_, _06718_);
  and (_21278_, _21202_, _06316_);
  or (_21279_, _21278_, _06047_);
  or (_21280_, _21279_, _21277_);
  and (_21282_, _14657_, _07724_);
  or (_21283_, _21197_, _06048_);
  or (_21284_, _21283_, _21282_);
  and (_21285_, _21284_, _01336_);
  and (_21286_, _21285_, _21280_);
  or (_21287_, _21286_, _21196_);
  and (_43368_, _21287_, _42882_);
  and (_21288_, _01340_, \oc8051_golden_model_1.DPH [3]);
  and (_21289_, _11359_, \oc8051_golden_model_1.DPH [3]);
  or (_21290_, _21289_, _08029_);
  and (_21292_, _07802_, _08662_);
  or (_21293_, _21292_, _21289_);
  and (_21294_, _21293_, _06108_);
  and (_21295_, _21294_, _21290_);
  or (_21296_, _21293_, _06020_);
  and (_21297_, _14672_, _07724_);
  or (_21298_, _21297_, _21289_);
  or (_21299_, _21298_, _06954_);
  and (_21300_, _07802_, \oc8051_golden_model_1.ACC [3]);
  or (_21301_, _21300_, _21289_);
  and (_21303_, _21301_, _06938_);
  and (_21304_, _06939_, \oc8051_golden_model_1.DPH [3]);
  or (_21305_, _21304_, _06102_);
  or (_21306_, _21305_, _21303_);
  and (_21307_, _21306_, _06848_);
  and (_21308_, _21307_, _21299_);
  nor (_21309_, _11359_, _07353_);
  or (_21310_, _21309_, _21289_);
  and (_21311_, _21310_, _06239_);
  or (_21312_, _21311_, _06219_);
  or (_21314_, _21312_, _21308_);
  or (_21315_, _21301_, _06220_);
  and (_21316_, _21315_, _11291_);
  and (_21317_, _21316_, _21314_);
  or (_21318_, _11390_, \oc8051_golden_model_1.DPH [3]);
  nor (_21319_, _11391_, _11291_);
  and (_21320_, _21319_, _21318_);
  or (_21321_, _21320_, _21317_);
  and (_21322_, _21321_, _06111_);
  nor (_21323_, _06111_, _05983_);
  or (_21325_, _21323_, _09818_);
  or (_21326_, _21325_, _21322_);
  or (_21327_, _21289_, _07012_);
  and (_21328_, _09181_, _07802_);
  or (_21329_, _21328_, _21327_);
  or (_21330_, _21310_, _09827_);
  and (_21331_, _21330_, _05669_);
  and (_21332_, _21331_, _21329_);
  and (_21333_, _21332_, _21326_);
  and (_21334_, _14778_, _07724_);
  or (_21336_, _21334_, _21289_);
  and (_21337_, _21336_, _09833_);
  or (_21338_, _21337_, _06019_);
  or (_21339_, _21338_, _21333_);
  and (_21340_, _21339_, _21296_);
  or (_21341_, _21340_, _06112_);
  and (_21342_, _14793_, _07802_);
  or (_21343_, _21342_, _21289_);
  or (_21344_, _21343_, _08751_);
  and (_21345_, _21344_, _08756_);
  and (_21347_, _21345_, _21341_);
  and (_21348_, _12299_, _07802_);
  or (_21349_, _21348_, _21289_);
  and (_21350_, _21349_, _06284_);
  or (_21351_, _21350_, _21347_);
  and (_21352_, _21351_, _07032_);
  or (_21353_, _21352_, _21295_);
  and (_21354_, _21353_, _06278_);
  and (_21355_, _21301_, _06277_);
  and (_21356_, _21355_, _21290_);
  or (_21358_, _21356_, _06130_);
  or (_21359_, _21358_, _21354_);
  and (_21360_, _14792_, _07724_);
  or (_21361_, _21289_, _08777_);
  or (_21362_, _21361_, _21360_);
  and (_21363_, _21362_, _08782_);
  and (_21364_, _21363_, _21359_);
  nor (_21365_, _10988_, _11359_);
  or (_21366_, _21365_, _21289_);
  and (_21367_, _21366_, _06292_);
  or (_21369_, _21367_, _21364_);
  and (_21370_, _21369_, _06718_);
  and (_21371_, _21298_, _06316_);
  or (_21372_, _21371_, _06047_);
  or (_21373_, _21372_, _21370_);
  and (_21374_, _14849_, _07724_);
  or (_21375_, _21289_, _06048_);
  or (_21376_, _21375_, _21374_);
  and (_21377_, _21376_, _01336_);
  and (_21378_, _21377_, _21373_);
  or (_21380_, _21378_, _21288_);
  and (_43369_, _21380_, _42882_);
  not (_21381_, \oc8051_golden_model_1.DPH [4]);
  nor (_21382_, _01336_, _21381_);
  nor (_21383_, _07802_, _21381_);
  or (_21384_, _21383_, _08273_);
  and (_21385_, _08665_, _07802_);
  or (_21386_, _21385_, _21383_);
  and (_21387_, _21386_, _06108_);
  and (_21388_, _21387_, _21384_);
  or (_21390_, _21386_, _06020_);
  and (_21391_, _14887_, _07724_);
  or (_21392_, _21391_, _21383_);
  or (_21393_, _21392_, _06954_);
  and (_21394_, _07802_, \oc8051_golden_model_1.ACC [4]);
  or (_21395_, _21394_, _21383_);
  and (_21396_, _21395_, _06938_);
  nor (_21397_, _06938_, _21381_);
  or (_21398_, _21397_, _06102_);
  or (_21399_, _21398_, _21396_);
  and (_21400_, _21399_, _06848_);
  and (_21401_, _21400_, _21393_);
  nor (_21402_, _08270_, _11359_);
  or (_21403_, _21402_, _21383_);
  and (_21404_, _21403_, _06239_);
  or (_21405_, _21404_, _06219_);
  or (_21406_, _21405_, _21401_);
  or (_21407_, _21395_, _06220_);
  and (_21408_, _21407_, _11291_);
  and (_21409_, _21408_, _21406_);
  or (_21412_, _11391_, \oc8051_golden_model_1.DPH [4]);
  nor (_21413_, _11392_, _11291_);
  and (_21414_, _21413_, _21412_);
  or (_21415_, _21414_, _21409_);
  and (_21416_, _21415_, _06111_);
  nor (_21417_, _06758_, _06111_);
  or (_21418_, _21417_, _09818_);
  or (_21419_, _21418_, _21416_);
  or (_21420_, _21383_, _07012_);
  and (_21421_, _09180_, _07802_);
  or (_21423_, _21421_, _21420_);
  or (_21424_, _21403_, _09827_);
  and (_21425_, _21424_, _05669_);
  and (_21426_, _21425_, _21423_);
  and (_21427_, _21426_, _21419_);
  and (_21428_, _14983_, _07724_);
  or (_21429_, _21428_, _21383_);
  and (_21430_, _21429_, _09833_);
  or (_21431_, _21430_, _06019_);
  or (_21432_, _21431_, _21427_);
  and (_21434_, _21432_, _21390_);
  or (_21435_, _21434_, _06112_);
  and (_21436_, _14876_, _07802_);
  or (_21437_, _21436_, _21383_);
  or (_21438_, _21437_, _08751_);
  and (_21439_, _21438_, _08756_);
  and (_21440_, _21439_, _21435_);
  and (_21441_, _10986_, _07802_);
  or (_21442_, _21441_, _21383_);
  and (_21443_, _21442_, _06284_);
  or (_21445_, _21443_, _21440_);
  and (_21446_, _21445_, _07032_);
  or (_21447_, _21446_, _21388_);
  and (_21448_, _21447_, _06278_);
  and (_21449_, _21395_, _06277_);
  and (_21450_, _21449_, _21384_);
  or (_21451_, _21450_, _06130_);
  or (_21452_, _21451_, _21448_);
  and (_21453_, _14873_, _07724_);
  or (_21454_, _21383_, _08777_);
  or (_21456_, _21454_, _21453_);
  and (_21457_, _21456_, _08782_);
  and (_21458_, _21457_, _21452_);
  nor (_21459_, _10985_, _11359_);
  or (_21460_, _21459_, _21383_);
  and (_21461_, _21460_, _06292_);
  or (_21462_, _21461_, _21458_);
  and (_21463_, _21462_, _06718_);
  and (_21464_, _21392_, _06316_);
  or (_21465_, _21464_, _06047_);
  or (_21467_, _21465_, _21463_);
  and (_21468_, _15055_, _07724_);
  or (_21469_, _21383_, _06048_);
  or (_21470_, _21469_, _21468_);
  and (_21471_, _21470_, _01336_);
  and (_21472_, _21471_, _21467_);
  or (_21473_, _21472_, _21382_);
  and (_43370_, _21473_, _42882_);
  and (_21474_, _01340_, \oc8051_golden_model_1.DPH [5]);
  and (_21475_, _11359_, \oc8051_golden_model_1.DPH [5]);
  and (_21477_, _08652_, _07802_);
  or (_21478_, _21477_, _21475_);
  or (_21479_, _21478_, _06020_);
  and (_21480_, _15093_, _07724_);
  or (_21481_, _21480_, _21475_);
  or (_21482_, _21481_, _06954_);
  and (_21483_, _07802_, \oc8051_golden_model_1.ACC [5]);
  or (_21484_, _21483_, _21475_);
  and (_21485_, _21484_, _06938_);
  and (_21486_, _06939_, \oc8051_golden_model_1.DPH [5]);
  or (_21488_, _21486_, _06102_);
  or (_21489_, _21488_, _21485_);
  and (_21490_, _21489_, _06848_);
  and (_21491_, _21490_, _21482_);
  nor (_21492_, _07977_, _11359_);
  or (_21493_, _21492_, _21475_);
  and (_21494_, _21493_, _06239_);
  or (_21495_, _21494_, _06219_);
  or (_21496_, _21495_, _21491_);
  or (_21497_, _21484_, _06220_);
  and (_21499_, _21497_, _11291_);
  and (_21500_, _21499_, _21496_);
  or (_21501_, _11392_, \oc8051_golden_model_1.DPH [5]);
  nor (_21502_, _11393_, _11291_);
  and (_21503_, _21502_, _21501_);
  or (_21504_, _21503_, _21500_);
  and (_21505_, _21504_, _06111_);
  nor (_21506_, _06359_, _06111_);
  or (_21507_, _21506_, _09818_);
  or (_21508_, _21507_, _21505_);
  or (_21510_, _21475_, _07012_);
  and (_21511_, _09179_, _07802_);
  or (_21512_, _21511_, _21510_);
  or (_21513_, _21493_, _09827_);
  and (_21514_, _21513_, _05669_);
  and (_21515_, _21514_, _21512_);
  and (_21516_, _21515_, _21508_);
  and (_21517_, _15179_, _07724_);
  or (_21518_, _21517_, _21475_);
  and (_21519_, _21518_, _09833_);
  or (_21521_, _21519_, _06019_);
  or (_21522_, _21521_, _21516_);
  and (_21523_, _21522_, _21479_);
  or (_21524_, _21523_, _06112_);
  and (_21525_, _15195_, _07802_);
  or (_21526_, _21525_, _21475_);
  or (_21527_, _21526_, _08751_);
  and (_21528_, _21527_, _08756_);
  and (_21529_, _21528_, _21524_);
  and (_21530_, _12306_, _07802_);
  or (_21532_, _21530_, _21475_);
  and (_21533_, _21532_, _06284_);
  or (_21534_, _21533_, _21529_);
  and (_21535_, _21534_, _07032_);
  or (_21536_, _21475_, _07980_);
  and (_21537_, _21478_, _06108_);
  and (_21538_, _21537_, _21536_);
  or (_21539_, _21538_, _21535_);
  and (_21540_, _21539_, _06278_);
  and (_21541_, _21484_, _06277_);
  and (_21543_, _21541_, _21536_);
  or (_21544_, _21543_, _06130_);
  or (_21545_, _21544_, _21540_);
  and (_21546_, _15194_, _07724_);
  or (_21547_, _21475_, _08777_);
  or (_21548_, _21547_, _21546_);
  and (_21549_, _21548_, _08782_);
  and (_21550_, _21549_, _21545_);
  nor (_21551_, _10982_, _11359_);
  or (_21552_, _21551_, _21475_);
  and (_21554_, _21552_, _06292_);
  or (_21555_, _21554_, _21550_);
  and (_21556_, _21555_, _06718_);
  and (_21557_, _21481_, _06316_);
  or (_21558_, _21557_, _06047_);
  or (_21559_, _21558_, _21556_);
  and (_21560_, _15253_, _07724_);
  or (_21561_, _21475_, _06048_);
  or (_21562_, _21561_, _21560_);
  and (_21563_, _21562_, _01336_);
  and (_21565_, _21563_, _21559_);
  or (_21566_, _21565_, _21474_);
  and (_43371_, _21566_, _42882_);
  and (_21567_, _01340_, \oc8051_golden_model_1.DPH [6]);
  and (_21568_, _11359_, \oc8051_golden_model_1.DPH [6]);
  and (_21569_, _15389_, _07802_);
  or (_21570_, _21569_, _21568_);
  or (_21571_, _21570_, _06020_);
  and (_21572_, _15293_, _07724_);
  or (_21573_, _21572_, _21568_);
  or (_21575_, _21573_, _06954_);
  and (_21576_, _07802_, \oc8051_golden_model_1.ACC [6]);
  or (_21577_, _21576_, _21568_);
  and (_21578_, _21577_, _06938_);
  and (_21579_, _06939_, \oc8051_golden_model_1.DPH [6]);
  or (_21580_, _21579_, _06102_);
  or (_21581_, _21580_, _21578_);
  and (_21582_, _21581_, _06848_);
  and (_21583_, _21582_, _21575_);
  nor (_21584_, _07883_, _11359_);
  or (_21586_, _21584_, _21568_);
  and (_21587_, _21586_, _06239_);
  or (_21588_, _21587_, _06219_);
  or (_21589_, _21588_, _21583_);
  or (_21590_, _21577_, _06220_);
  and (_21591_, _21590_, _11291_);
  and (_21592_, _21591_, _21589_);
  or (_21593_, _11393_, \oc8051_golden_model_1.DPH [6]);
  nor (_21594_, _11394_, _11291_);
  and (_21595_, _21594_, _21593_);
  or (_21597_, _21595_, _21592_);
  and (_21598_, _21597_, _06111_);
  nor (_21599_, _06111_, _06084_);
  or (_21600_, _21599_, _09818_);
  or (_21601_, _21600_, _21598_);
  or (_21602_, _21568_, _07012_);
  and (_21603_, _09178_, _07802_);
  or (_21604_, _21603_, _21602_);
  or (_21605_, _21586_, _09827_);
  and (_21606_, _21605_, _05669_);
  and (_21608_, _21606_, _21604_);
  and (_21609_, _21608_, _21601_);
  and (_21610_, _15382_, _07724_);
  or (_21611_, _21610_, _21568_);
  and (_21612_, _21611_, _09833_);
  or (_21613_, _21612_, _06019_);
  or (_21614_, _21613_, _21609_);
  and (_21615_, _21614_, _21571_);
  or (_21616_, _21615_, _06112_);
  and (_21617_, _15399_, _07724_);
  or (_21619_, _21568_, _08751_);
  or (_21620_, _21619_, _21617_);
  and (_21621_, _21620_, _08756_);
  and (_21622_, _21621_, _21616_);
  and (_21623_, _10980_, _07802_);
  or (_21624_, _21623_, _21568_);
  and (_21625_, _21624_, _06284_);
  or (_21626_, _21625_, _21622_);
  and (_21627_, _21626_, _07032_);
  or (_21628_, _21568_, _07886_);
  and (_21630_, _21570_, _06108_);
  and (_21631_, _21630_, _21628_);
  or (_21632_, _21631_, _21627_);
  and (_21633_, _21632_, _06278_);
  and (_21634_, _21577_, _06277_);
  and (_21635_, _21634_, _21628_);
  or (_21636_, _21635_, _06130_);
  or (_21637_, _21636_, _21633_);
  and (_21638_, _15396_, _07724_);
  or (_21639_, _21568_, _08777_);
  or (_21641_, _21639_, _21638_);
  and (_21642_, _21641_, _08782_);
  and (_21643_, _21642_, _21637_);
  nor (_21644_, _10979_, _11359_);
  or (_21645_, _21644_, _21568_);
  and (_21646_, _21645_, _06292_);
  or (_21647_, _21646_, _21643_);
  and (_21648_, _21647_, _06718_);
  and (_21649_, _21573_, _06316_);
  or (_21650_, _21649_, _06047_);
  or (_21652_, _21650_, _21648_);
  and (_21653_, _15451_, _07724_);
  or (_21654_, _21568_, _06048_);
  or (_21655_, _21654_, _21653_);
  and (_21656_, _21655_, _01336_);
  and (_21657_, _21656_, _21652_);
  or (_21658_, _21657_, _21567_);
  and (_43372_, _21658_, _42882_);
  not (_21659_, \oc8051_golden_model_1.TL1 [0]);
  nor (_21660_, _01336_, _21659_);
  nand (_21662_, _10995_, _07667_);
  nor (_21663_, _07667_, _21659_);
  nor (_21664_, _21663_, _06278_);
  nand (_21665_, _21664_, _21662_);
  and (_21666_, _09120_, _07667_);
  or (_21667_, _21663_, _07012_);
  or (_21668_, _21667_, _21666_);
  and (_21669_, _07667_, _06931_);
  nor (_21670_, _21669_, _21663_);
  nand (_21671_, _21670_, _09815_);
  nor (_21673_, _08127_, _11451_);
  or (_21674_, _21673_, _21663_);
  or (_21675_, _21674_, _06954_);
  and (_21676_, _07667_, \oc8051_golden_model_1.ACC [0]);
  nor (_21677_, _21676_, _21663_);
  nor (_21678_, _21677_, _06939_);
  nor (_21679_, _06938_, _21659_);
  or (_21680_, _21679_, _06102_);
  or (_21681_, _21680_, _21678_);
  and (_21682_, _21681_, _06848_);
  and (_21684_, _21682_, _21675_);
  nor (_21685_, _21670_, _06848_);
  or (_21686_, _21685_, _21684_);
  nand (_21687_, _21686_, _06220_);
  or (_21688_, _21677_, _06220_);
  and (_21689_, _21688_, _09817_);
  nand (_21690_, _21689_, _21687_);
  and (_21691_, _21690_, _21671_);
  and (_21692_, _21691_, _21668_);
  or (_21693_, _21692_, _09833_);
  and (_21695_, _14186_, _07667_);
  or (_21696_, _21663_, _05669_);
  or (_21697_, _21696_, _21695_);
  and (_21698_, _21697_, _06020_);
  and (_21699_, _21698_, _21693_);
  and (_21700_, _07667_, _08672_);
  or (_21701_, _21700_, _21663_);
  and (_21702_, _21701_, _06019_);
  or (_21703_, _21702_, _06112_);
  or (_21704_, _21703_, _21699_);
  and (_21706_, _14086_, _07667_);
  or (_21707_, _21663_, _08751_);
  or (_21708_, _21707_, _21706_);
  and (_21709_, _21708_, _08756_);
  and (_21710_, _21709_, _21704_);
  nor (_21711_, _12302_, _11451_);
  or (_21712_, _21711_, _21663_);
  and (_21713_, _21662_, _06284_);
  and (_21714_, _21713_, _21712_);
  or (_21715_, _21714_, _21710_);
  and (_21717_, _21715_, _07032_);
  nand (_21718_, _21701_, _06108_);
  nor (_21719_, _21718_, _21673_);
  or (_21720_, _21719_, _06277_);
  or (_21721_, _21720_, _21717_);
  and (_21722_, _21721_, _21665_);
  or (_21723_, _21722_, _06130_);
  and (_21724_, _14083_, _07667_);
  or (_21725_, _21663_, _08777_);
  or (_21726_, _21725_, _21724_);
  and (_21728_, _21726_, _08782_);
  and (_21729_, _21728_, _21723_);
  and (_21730_, _21712_, _06292_);
  or (_21731_, _21730_, _19256_);
  or (_21732_, _21731_, _21729_);
  or (_21733_, _21674_, _06408_);
  and (_21734_, _21733_, _01336_);
  and (_21735_, _21734_, _21732_);
  or (_21736_, _21735_, _21660_);
  and (_43374_, _21736_, _42882_);
  not (_21738_, \oc8051_golden_model_1.TL1 [1]);
  nor (_21739_, _01336_, _21738_);
  or (_21740_, _14367_, _11451_);
  or (_21741_, _07667_, \oc8051_golden_model_1.TL1 [1]);
  and (_21742_, _21741_, _09833_);
  and (_21743_, _21742_, _21740_);
  and (_21744_, _09075_, _07667_);
  nor (_21745_, _07667_, _21738_);
  or (_21746_, _21745_, _07012_);
  or (_21747_, _21746_, _21744_);
  and (_21748_, _14284_, _07667_);
  not (_21749_, _21748_);
  and (_21750_, _21749_, _21741_);
  or (_21751_, _21750_, _06954_);
  and (_21752_, _07667_, \oc8051_golden_model_1.ACC [1]);
  or (_21753_, _21752_, _21745_);
  and (_21754_, _21753_, _06938_);
  nor (_21755_, _06938_, _21738_);
  or (_21756_, _21755_, _06102_);
  or (_21757_, _21756_, _21754_);
  and (_21760_, _21757_, _06848_);
  and (_21761_, _21760_, _21751_);
  nor (_21762_, _11451_, _07132_);
  or (_21763_, _21762_, _21745_);
  and (_21764_, _21763_, _06239_);
  or (_21765_, _21764_, _21761_);
  and (_21766_, _21765_, _06220_);
  and (_21767_, _21753_, _06219_);
  or (_21768_, _21767_, _09818_);
  or (_21769_, _21768_, _21766_);
  or (_21771_, _21763_, _09827_);
  and (_21772_, _21771_, _05669_);
  and (_21773_, _21772_, _21769_);
  and (_21774_, _21773_, _21747_);
  or (_21775_, _21774_, _21743_);
  and (_21776_, _21775_, _06020_);
  nand (_21777_, _07667_, _06832_);
  and (_21778_, _21741_, _06019_);
  and (_21779_, _21778_, _21777_);
  or (_21780_, _21779_, _21776_);
  and (_21782_, _21780_, _08751_);
  or (_21783_, _14263_, _11451_);
  and (_21784_, _21741_, _06112_);
  and (_21785_, _21784_, _21783_);
  or (_21786_, _21785_, _06284_);
  or (_21787_, _21786_, _21782_);
  nor (_21788_, _10993_, _11451_);
  or (_21789_, _21788_, _21745_);
  nand (_21790_, _10992_, _07667_);
  and (_21791_, _21790_, _21789_);
  or (_21793_, _21791_, _08756_);
  and (_21794_, _21793_, _07032_);
  and (_21795_, _21794_, _21787_);
  or (_21796_, _14261_, _11451_);
  and (_21797_, _21741_, _06108_);
  and (_21798_, _21797_, _21796_);
  or (_21799_, _21798_, _06277_);
  or (_21800_, _21799_, _21795_);
  nor (_21801_, _21745_, _06278_);
  nand (_21802_, _21801_, _21790_);
  and (_21804_, _21802_, _08777_);
  and (_21805_, _21804_, _21800_);
  or (_21806_, _21777_, _08078_);
  and (_21807_, _21741_, _06130_);
  and (_21808_, _21807_, _21806_);
  or (_21809_, _21808_, _06292_);
  or (_21810_, _21809_, _21805_);
  or (_21811_, _21789_, _08782_);
  and (_21812_, _21811_, _06718_);
  and (_21813_, _21812_, _21810_);
  and (_21815_, _21750_, _06316_);
  or (_21816_, _21815_, _06047_);
  or (_21817_, _21816_, _21813_);
  or (_21818_, _21745_, _06048_);
  or (_21819_, _21818_, _21748_);
  and (_21820_, _21819_, _01336_);
  and (_21821_, _21820_, _21817_);
  or (_21822_, _21821_, _21739_);
  and (_43375_, _21822_, _42882_);
  not (_21823_, \oc8051_golden_model_1.TL1 [2]);
  nor (_21825_, _01336_, _21823_);
  and (_21826_, _09182_, _07667_);
  nor (_21827_, _07667_, _21823_);
  or (_21828_, _21827_, _07012_);
  or (_21829_, _21828_, _21826_);
  nor (_21830_, _11451_, _07530_);
  nor (_21831_, _21830_, _21827_);
  nand (_21832_, _21831_, _09815_);
  and (_21833_, _14493_, _07667_);
  or (_21834_, _21833_, _21827_);
  and (_21836_, _21834_, _06102_);
  nor (_21837_, _06938_, _21823_);
  and (_21838_, _07667_, \oc8051_golden_model_1.ACC [2]);
  nor (_21839_, _21838_, _21827_);
  nor (_21840_, _21839_, _06939_);
  or (_21841_, _21840_, _21837_);
  and (_21842_, _21841_, _06954_);
  or (_21843_, _21842_, _06239_);
  or (_21844_, _21843_, _21836_);
  nand (_21845_, _21831_, _06239_);
  and (_21847_, _21845_, _06220_);
  nand (_21848_, _21847_, _21844_);
  or (_21849_, _21839_, _06220_);
  and (_21850_, _21849_, _09817_);
  nand (_21851_, _21850_, _21848_);
  and (_21852_, _21851_, _21832_);
  and (_21853_, _21852_, _21829_);
  or (_21854_, _21853_, _09833_);
  and (_21855_, _14580_, _07667_);
  or (_21856_, _21855_, _21827_);
  or (_21857_, _21856_, _05669_);
  and (_21858_, _21857_, _06020_);
  and (_21859_, _21858_, _21854_);
  and (_21860_, _07667_, _08730_);
  or (_21861_, _21860_, _21827_);
  and (_21862_, _21861_, _06019_);
  or (_21863_, _21862_, _06112_);
  or (_21864_, _21863_, _21859_);
  and (_21865_, _14596_, _07667_);
  or (_21866_, _21827_, _08751_);
  or (_21869_, _21866_, _21865_);
  and (_21870_, _21869_, _08756_);
  and (_21871_, _21870_, _21864_);
  and (_21872_, _10991_, _07667_);
  or (_21873_, _21872_, _21827_);
  and (_21874_, _21873_, _06284_);
  or (_21875_, _21874_, _21871_);
  and (_21876_, _21875_, _07032_);
  or (_21877_, _21827_, _08177_);
  and (_21878_, _21861_, _06108_);
  and (_21880_, _21878_, _21877_);
  or (_21881_, _21880_, _21876_);
  and (_21882_, _21881_, _06278_);
  nor (_21883_, _21839_, _06278_);
  and (_21884_, _21883_, _21877_);
  or (_21885_, _21884_, _06130_);
  or (_21886_, _21885_, _21882_);
  and (_21887_, _14593_, _07667_);
  or (_21888_, _21827_, _08777_);
  or (_21889_, _21888_, _21887_);
  and (_21891_, _21889_, _08782_);
  and (_21892_, _21891_, _21886_);
  nor (_21893_, _10990_, _11451_);
  or (_21894_, _21893_, _21827_);
  and (_21895_, _21894_, _06292_);
  or (_21896_, _21895_, _21892_);
  and (_21897_, _21896_, _06718_);
  and (_21898_, _21834_, _06316_);
  or (_21899_, _21898_, _06047_);
  or (_21900_, _21899_, _21897_);
  and (_21902_, _14657_, _07667_);
  or (_21903_, _21827_, _06048_);
  or (_21904_, _21903_, _21902_);
  and (_21905_, _21904_, _01336_);
  and (_21906_, _21905_, _21900_);
  or (_21907_, _21906_, _21825_);
  and (_43376_, _21907_, _42882_);
  not (_21908_, \oc8051_golden_model_1.TL1 [3]);
  nor (_21909_, _01336_, _21908_);
  and (_21910_, _09181_, _07667_);
  nor (_21912_, _07667_, _21908_);
  or (_21913_, _21912_, _07012_);
  or (_21914_, _21913_, _21910_);
  nor (_21915_, _11451_, _07353_);
  nor (_21916_, _21915_, _21912_);
  nand (_21917_, _21916_, _09815_);
  and (_21918_, _14672_, _07667_);
  or (_21919_, _21918_, _21912_);
  or (_21920_, _21919_, _06954_);
  and (_21921_, _07667_, \oc8051_golden_model_1.ACC [3]);
  nor (_21923_, _21921_, _21912_);
  nor (_21924_, _21923_, _06939_);
  nor (_21925_, _06938_, _21908_);
  or (_21926_, _21925_, _06102_);
  or (_21927_, _21926_, _21924_);
  and (_21928_, _21927_, _06848_);
  and (_21929_, _21928_, _21920_);
  nor (_21930_, _21916_, _06848_);
  or (_21931_, _21930_, _21929_);
  nand (_21932_, _21931_, _06220_);
  or (_21934_, _21923_, _06220_);
  and (_21935_, _21934_, _09817_);
  nand (_21936_, _21935_, _21932_);
  and (_21937_, _21936_, _21917_);
  and (_21938_, _21937_, _21914_);
  or (_21939_, _21938_, _09833_);
  and (_21940_, _14778_, _07667_);
  or (_21941_, _21912_, _05669_);
  or (_21942_, _21941_, _21940_);
  and (_21943_, _21942_, _06020_);
  and (_21945_, _21943_, _21939_);
  and (_21946_, _07667_, _08662_);
  or (_21947_, _21946_, _21912_);
  and (_21948_, _21947_, _06019_);
  or (_21949_, _21948_, _06112_);
  or (_21950_, _21949_, _21945_);
  and (_21951_, _14793_, _07667_);
  or (_21952_, _21912_, _08751_);
  or (_21953_, _21952_, _21951_);
  and (_21954_, _21953_, _08756_);
  and (_21956_, _21954_, _21950_);
  and (_21957_, _12299_, _07667_);
  or (_21958_, _21957_, _21912_);
  and (_21959_, _21958_, _06284_);
  or (_21960_, _21959_, _21956_);
  and (_21961_, _21960_, _07032_);
  or (_21962_, _21912_, _08029_);
  and (_21963_, _21947_, _06108_);
  and (_21964_, _21963_, _21962_);
  or (_21965_, _21964_, _21961_);
  and (_21967_, _21965_, _06278_);
  nor (_21968_, _21923_, _06278_);
  and (_21969_, _21968_, _21962_);
  or (_21970_, _21969_, _06130_);
  or (_21971_, _21970_, _21967_);
  and (_21972_, _14792_, _07667_);
  or (_21973_, _21912_, _08777_);
  or (_21974_, _21973_, _21972_);
  and (_21975_, _21974_, _08782_);
  and (_21976_, _21975_, _21971_);
  nor (_21978_, _10988_, _11451_);
  or (_21979_, _21978_, _21912_);
  and (_21980_, _21979_, _06292_);
  or (_21981_, _21980_, _21976_);
  and (_21982_, _21981_, _06718_);
  and (_21983_, _21919_, _06316_);
  or (_21984_, _21983_, _06047_);
  or (_21985_, _21984_, _21982_);
  and (_21986_, _14849_, _07667_);
  or (_21987_, _21912_, _06048_);
  or (_21989_, _21987_, _21986_);
  and (_21990_, _21989_, _01336_);
  and (_21991_, _21990_, _21985_);
  or (_21992_, _21991_, _21909_);
  and (_43377_, _21992_, _42882_);
  and (_21993_, _01340_, \oc8051_golden_model_1.TL1 [4]);
  and (_21994_, _11451_, \oc8051_golden_model_1.TL1 [4]);
  and (_21995_, _08665_, _07667_);
  or (_21996_, _21995_, _21994_);
  or (_21997_, _21996_, _06020_);
  and (_21999_, _14887_, _07667_);
  or (_22000_, _21999_, _21994_);
  or (_22001_, _22000_, _06954_);
  and (_22002_, _07667_, \oc8051_golden_model_1.ACC [4]);
  or (_22003_, _22002_, _21994_);
  and (_22004_, _22003_, _06938_);
  and (_22005_, _06939_, \oc8051_golden_model_1.TL1 [4]);
  or (_22006_, _22005_, _06102_);
  or (_22007_, _22006_, _22004_);
  and (_22008_, _22007_, _06848_);
  and (_22010_, _22008_, _22001_);
  nor (_22011_, _08270_, _11451_);
  or (_22012_, _22011_, _21994_);
  and (_22013_, _22012_, _06239_);
  or (_22014_, _22013_, _22010_);
  and (_22015_, _22014_, _06220_);
  and (_22016_, _22003_, _06219_);
  or (_22017_, _22016_, _09818_);
  or (_22018_, _22017_, _22015_);
  and (_22019_, _09180_, _07667_);
  or (_22021_, _21994_, _07012_);
  or (_22022_, _22021_, _22019_);
  or (_22023_, _22012_, _09827_);
  and (_22024_, _22023_, _05669_);
  and (_22025_, _22024_, _22022_);
  and (_22026_, _22025_, _22018_);
  and (_22027_, _14983_, _07667_);
  or (_22028_, _22027_, _21994_);
  and (_22029_, _22028_, _09833_);
  or (_22030_, _22029_, _06019_);
  or (_22032_, _22030_, _22026_);
  and (_22033_, _22032_, _21997_);
  or (_22034_, _22033_, _06112_);
  and (_22035_, _14876_, _07667_);
  or (_22036_, _21994_, _08751_);
  or (_22037_, _22036_, _22035_);
  and (_22038_, _22037_, _08756_);
  and (_22039_, _22038_, _22034_);
  and (_22040_, _10986_, _07667_);
  or (_22041_, _22040_, _21994_);
  and (_22043_, _22041_, _06284_);
  or (_22044_, _22043_, _22039_);
  and (_22045_, _22044_, _07032_);
  or (_22046_, _21994_, _08273_);
  and (_22047_, _21996_, _06108_);
  and (_22048_, _22047_, _22046_);
  or (_22049_, _22048_, _22045_);
  and (_22050_, _22049_, _06278_);
  and (_22051_, _22003_, _06277_);
  and (_22052_, _22051_, _22046_);
  or (_22054_, _22052_, _06130_);
  or (_22055_, _22054_, _22050_);
  and (_22056_, _14873_, _07667_);
  or (_22057_, _21994_, _08777_);
  or (_22058_, _22057_, _22056_);
  and (_22059_, _22058_, _08782_);
  and (_22060_, _22059_, _22055_);
  nor (_22061_, _10985_, _11451_);
  or (_22062_, _22061_, _21994_);
  and (_22063_, _22062_, _06292_);
  or (_22065_, _22063_, _22060_);
  and (_22066_, _22065_, _06718_);
  and (_22067_, _22000_, _06316_);
  or (_22068_, _22067_, _06047_);
  or (_22069_, _22068_, _22066_);
  and (_22070_, _15055_, _07667_);
  or (_22071_, _21994_, _06048_);
  or (_22072_, _22071_, _22070_);
  and (_22073_, _22072_, _01336_);
  and (_22074_, _22073_, _22069_);
  or (_22076_, _22074_, _21993_);
  and (_43378_, _22076_, _42882_);
  and (_22077_, _01340_, \oc8051_golden_model_1.TL1 [5]);
  and (_22078_, _11451_, \oc8051_golden_model_1.TL1 [5]);
  and (_22079_, _08652_, _07667_);
  or (_22080_, _22079_, _22078_);
  or (_22081_, _22080_, _06020_);
  and (_22082_, _15093_, _07667_);
  or (_22083_, _22082_, _22078_);
  or (_22084_, _22083_, _06954_);
  and (_22086_, _07667_, \oc8051_golden_model_1.ACC [5]);
  or (_22087_, _22086_, _22078_);
  and (_22088_, _22087_, _06938_);
  and (_22089_, _06939_, \oc8051_golden_model_1.TL1 [5]);
  or (_22090_, _22089_, _06102_);
  or (_22091_, _22090_, _22088_);
  and (_22092_, _22091_, _06848_);
  and (_22093_, _22092_, _22084_);
  nor (_22094_, _07977_, _11451_);
  or (_22095_, _22094_, _22078_);
  and (_22097_, _22095_, _06239_);
  or (_22098_, _22097_, _22093_);
  and (_22099_, _22098_, _06220_);
  and (_22100_, _22087_, _06219_);
  or (_22101_, _22100_, _09818_);
  or (_22102_, _22101_, _22099_);
  and (_22103_, _09179_, _07667_);
  or (_22104_, _22078_, _07012_);
  or (_22105_, _22104_, _22103_);
  or (_22106_, _22095_, _09827_);
  and (_22108_, _22106_, _05669_);
  and (_22109_, _22108_, _22105_);
  and (_22110_, _22109_, _22102_);
  and (_22111_, _15179_, _07667_);
  or (_22112_, _22111_, _22078_);
  and (_22113_, _22112_, _09833_);
  or (_22114_, _22113_, _06019_);
  or (_22115_, _22114_, _22110_);
  and (_22116_, _22115_, _22081_);
  or (_22117_, _22116_, _06112_);
  and (_22119_, _15195_, _07667_);
  or (_22120_, _22119_, _22078_);
  or (_22121_, _22120_, _08751_);
  and (_22122_, _22121_, _08756_);
  and (_22123_, _22122_, _22117_);
  and (_22124_, _12306_, _07667_);
  or (_22125_, _22124_, _22078_);
  and (_22126_, _22125_, _06284_);
  or (_22127_, _22126_, _22123_);
  and (_22128_, _22127_, _07032_);
  or (_22130_, _22078_, _07980_);
  and (_22131_, _22080_, _06108_);
  and (_22132_, _22131_, _22130_);
  or (_22133_, _22132_, _22128_);
  and (_22134_, _22133_, _06278_);
  and (_22135_, _22087_, _06277_);
  and (_22136_, _22135_, _22130_);
  or (_22137_, _22136_, _06130_);
  or (_22138_, _22137_, _22134_);
  and (_22139_, _15194_, _07667_);
  or (_22141_, _22078_, _08777_);
  or (_22142_, _22141_, _22139_);
  and (_22143_, _22142_, _08782_);
  and (_22144_, _22143_, _22138_);
  nor (_22145_, _10982_, _11451_);
  or (_22146_, _22145_, _22078_);
  and (_22147_, _22146_, _06292_);
  or (_22148_, _22147_, _22144_);
  and (_22149_, _22148_, _06718_);
  and (_22150_, _22083_, _06316_);
  or (_22152_, _22150_, _06047_);
  or (_22153_, _22152_, _22149_);
  and (_22154_, _15253_, _07667_);
  or (_22155_, _22078_, _06048_);
  or (_22156_, _22155_, _22154_);
  and (_22157_, _22156_, _01336_);
  and (_22158_, _22157_, _22153_);
  or (_22159_, _22158_, _22077_);
  and (_43380_, _22159_, _42882_);
  and (_22160_, _01340_, \oc8051_golden_model_1.TL1 [6]);
  and (_22162_, _11451_, \oc8051_golden_model_1.TL1 [6]);
  and (_22163_, _15389_, _07667_);
  or (_22164_, _22163_, _22162_);
  or (_22165_, _22164_, _06020_);
  and (_22166_, _15293_, _07667_);
  or (_22167_, _22166_, _22162_);
  or (_22168_, _22167_, _06954_);
  and (_22169_, _07667_, \oc8051_golden_model_1.ACC [6]);
  or (_22170_, _22169_, _22162_);
  and (_22171_, _22170_, _06938_);
  and (_22173_, _06939_, \oc8051_golden_model_1.TL1 [6]);
  or (_22174_, _22173_, _06102_);
  or (_22175_, _22174_, _22171_);
  and (_22176_, _22175_, _06848_);
  and (_22177_, _22176_, _22168_);
  nor (_22178_, _07883_, _11451_);
  or (_22179_, _22178_, _22162_);
  and (_22180_, _22179_, _06239_);
  or (_22181_, _22180_, _22177_);
  and (_22182_, _22181_, _06220_);
  and (_22184_, _22170_, _06219_);
  or (_22185_, _22184_, _09818_);
  or (_22186_, _22185_, _22182_);
  and (_22187_, _09178_, _07667_);
  or (_22188_, _22162_, _07012_);
  or (_22189_, _22188_, _22187_);
  or (_22190_, _22179_, _09827_);
  and (_22191_, _22190_, _05669_);
  and (_22192_, _22191_, _22189_);
  and (_22193_, _22192_, _22186_);
  and (_22195_, _15382_, _07667_);
  or (_22196_, _22195_, _22162_);
  and (_22197_, _22196_, _09833_);
  or (_22198_, _22197_, _06019_);
  or (_22199_, _22198_, _22193_);
  and (_22200_, _22199_, _22165_);
  or (_22201_, _22200_, _06112_);
  and (_22202_, _15399_, _07667_);
  or (_22203_, _22162_, _08751_);
  or (_22204_, _22203_, _22202_);
  and (_22206_, _22204_, _08756_);
  and (_22207_, _22206_, _22201_);
  and (_22208_, _10980_, _07667_);
  or (_22209_, _22208_, _22162_);
  and (_22210_, _22209_, _06284_);
  or (_22211_, _22210_, _22207_);
  and (_22212_, _22211_, _07032_);
  or (_22213_, _22162_, _07886_);
  and (_22214_, _22164_, _06108_);
  and (_22215_, _22214_, _22213_);
  or (_22218_, _22215_, _22212_);
  and (_22219_, _22218_, _06278_);
  and (_22220_, _22170_, _06277_);
  and (_22221_, _22220_, _22213_);
  or (_22222_, _22221_, _06130_);
  or (_22223_, _22222_, _22219_);
  and (_22224_, _15396_, _07667_);
  or (_22225_, _22162_, _08777_);
  or (_22226_, _22225_, _22224_);
  and (_22227_, _22226_, _08782_);
  and (_22229_, _22227_, _22223_);
  nor (_22230_, _10979_, _11451_);
  or (_22231_, _22230_, _22162_);
  and (_22232_, _22231_, _06292_);
  or (_22233_, _22232_, _22229_);
  and (_22234_, _22233_, _06718_);
  and (_22235_, _22167_, _06316_);
  or (_22236_, _22235_, _06047_);
  or (_22237_, _22236_, _22234_);
  and (_22238_, _15451_, _07667_);
  or (_22240_, _22162_, _06048_);
  or (_22241_, _22240_, _22238_);
  and (_22242_, _22241_, _01336_);
  and (_22243_, _22242_, _22237_);
  or (_22244_, _22243_, _22160_);
  and (_43381_, _22244_, _42882_);
  not (_22245_, \oc8051_golden_model_1.TL0 [0]);
  nor (_22246_, _01336_, _22245_);
  nand (_22247_, _10995_, _07659_);
  nor (_22248_, _07659_, _22245_);
  nor (_22250_, _22248_, _06278_);
  nand (_22251_, _22250_, _22247_);
  and (_22252_, _09120_, _07659_);
  or (_22253_, _22248_, _07012_);
  or (_22254_, _22253_, _22252_);
  and (_22255_, _07659_, _06931_);
  nor (_22256_, _22255_, _22248_);
  nand (_22257_, _22256_, _09815_);
  nor (_22258_, _08127_, _11528_);
  or (_22259_, _22258_, _22248_);
  and (_22261_, _22259_, _06102_);
  nor (_22262_, _06938_, _22245_);
  and (_22263_, _07659_, \oc8051_golden_model_1.ACC [0]);
  nor (_22264_, _22263_, _22248_);
  nor (_22265_, _22264_, _06939_);
  or (_22266_, _22265_, _22262_);
  and (_22267_, _22266_, _06954_);
  or (_22268_, _22267_, _06239_);
  or (_22269_, _22268_, _22261_);
  nand (_22270_, _22256_, _06239_);
  and (_22272_, _22270_, _06220_);
  nand (_22273_, _22272_, _22269_);
  or (_22274_, _22264_, _06220_);
  and (_22275_, _22274_, _09817_);
  nand (_22276_, _22275_, _22273_);
  and (_22277_, _22276_, _22257_);
  and (_22278_, _22277_, _22254_);
  or (_22279_, _22278_, _09833_);
  and (_22280_, _14186_, _07659_);
  or (_22281_, _22248_, _05669_);
  or (_22283_, _22281_, _22280_);
  and (_22284_, _22283_, _06020_);
  and (_22285_, _22284_, _22279_);
  and (_22286_, _07659_, _08672_);
  or (_22287_, _22286_, _22248_);
  and (_22288_, _22287_, _06019_);
  or (_22289_, _22288_, _06112_);
  or (_22290_, _22289_, _22285_);
  and (_22291_, _14086_, _07659_);
  or (_22292_, _22291_, _22248_);
  or (_22294_, _22292_, _08751_);
  and (_22295_, _22294_, _08756_);
  and (_22296_, _22295_, _22290_);
  nor (_22297_, _12302_, _11528_);
  or (_22298_, _22297_, _22248_);
  and (_22299_, _22247_, _06284_);
  and (_22300_, _22299_, _22298_);
  or (_22301_, _22300_, _22296_);
  and (_22302_, _22301_, _07032_);
  nand (_22303_, _22287_, _06108_);
  nor (_22304_, _22303_, _22258_);
  or (_22305_, _22304_, _06277_);
  or (_22306_, _22305_, _22302_);
  and (_22307_, _22306_, _22251_);
  or (_22308_, _22307_, _06130_);
  and (_22309_, _14083_, _07659_);
  or (_22310_, _22248_, _08777_);
  or (_22311_, _22310_, _22309_);
  and (_22312_, _22311_, _08782_);
  and (_22313_, _22312_, _22308_);
  and (_22316_, _22298_, _06292_);
  or (_22317_, _22316_, _19256_);
  or (_22318_, _22317_, _22313_);
  or (_22319_, _22259_, _06408_);
  and (_22320_, _22319_, _01336_);
  and (_22321_, _22320_, _22318_);
  or (_22322_, _22321_, _22246_);
  and (_43382_, _22322_, _42882_);
  not (_22323_, \oc8051_golden_model_1.TL0 [1]);
  nor (_22324_, _01336_, _22323_);
  or (_22326_, _14367_, _11528_);
  or (_22327_, _07659_, \oc8051_golden_model_1.TL0 [1]);
  and (_22328_, _22327_, _09833_);
  and (_22329_, _22328_, _22326_);
  and (_22330_, _09075_, _07659_);
  nor (_22331_, _07659_, _22323_);
  or (_22332_, _22331_, _07012_);
  or (_22333_, _22332_, _22330_);
  and (_22334_, _14284_, _07659_);
  not (_22335_, _22334_);
  and (_22337_, _22335_, _22327_);
  and (_22338_, _22337_, _06102_);
  nor (_22339_, _06938_, _22323_);
  and (_22340_, _07659_, \oc8051_golden_model_1.ACC [1]);
  or (_22341_, _22340_, _22331_);
  and (_22342_, _22341_, _06938_);
  or (_22343_, _22342_, _22339_);
  and (_22344_, _22343_, _06954_);
  or (_22345_, _22344_, _06239_);
  or (_22346_, _22345_, _22338_);
  nor (_22348_, _11528_, _07132_);
  or (_22349_, _22348_, _22331_);
  or (_22350_, _22349_, _06848_);
  and (_22351_, _22350_, _06220_);
  and (_22352_, _22351_, _22346_);
  and (_22353_, _22341_, _06219_);
  or (_22354_, _22353_, _09818_);
  or (_22355_, _22354_, _22352_);
  or (_22356_, _22349_, _09827_);
  and (_22357_, _22356_, _05669_);
  and (_22359_, _22357_, _22355_);
  and (_22360_, _22359_, _22333_);
  or (_22361_, _22360_, _22329_);
  and (_22362_, _22361_, _06020_);
  nand (_22363_, _07659_, _06832_);
  and (_22364_, _22327_, _06019_);
  and (_22365_, _22364_, _22363_);
  or (_22366_, _22365_, _22362_);
  and (_22367_, _22366_, _08751_);
  or (_22368_, _14263_, _11528_);
  and (_22370_, _22327_, _06112_);
  and (_22371_, _22370_, _22368_);
  or (_22372_, _22371_, _06284_);
  or (_22373_, _22372_, _22367_);
  nor (_22374_, _10993_, _11528_);
  or (_22375_, _22374_, _22331_);
  nand (_22376_, _10992_, _07659_);
  and (_22377_, _22376_, _22375_);
  or (_22378_, _22377_, _08756_);
  and (_22379_, _22378_, _07032_);
  and (_22381_, _22379_, _22373_);
  or (_22382_, _14261_, _11528_);
  and (_22383_, _22327_, _06108_);
  and (_22384_, _22383_, _22382_);
  or (_22385_, _22384_, _06277_);
  or (_22386_, _22385_, _22381_);
  nor (_22387_, _22331_, _06278_);
  nand (_22388_, _22387_, _22376_);
  and (_22389_, _22388_, _08777_);
  and (_22390_, _22389_, _22386_);
  or (_22392_, _22363_, _08078_);
  and (_22393_, _22327_, _06130_);
  and (_22394_, _22393_, _22392_);
  or (_22395_, _22394_, _06292_);
  or (_22396_, _22395_, _22390_);
  or (_22397_, _22375_, _08782_);
  and (_22398_, _22397_, _06718_);
  and (_22399_, _22398_, _22396_);
  and (_22400_, _22337_, _06316_);
  or (_22401_, _22400_, _06047_);
  or (_22403_, _22401_, _22399_);
  or (_22404_, _22331_, _06048_);
  or (_22405_, _22404_, _22334_);
  and (_22406_, _22405_, _01336_);
  and (_22407_, _22406_, _22403_);
  or (_22408_, _22407_, _22324_);
  and (_43384_, _22408_, _42882_);
  not (_22409_, \oc8051_golden_model_1.TL0 [2]);
  nor (_22410_, _01336_, _22409_);
  and (_22411_, _09182_, _07659_);
  nor (_22413_, _07659_, _22409_);
  or (_22414_, _22413_, _07012_);
  or (_22415_, _22414_, _22411_);
  nor (_22416_, _11528_, _07530_);
  nor (_22417_, _22416_, _22413_);
  nand (_22418_, _22417_, _09815_);
  and (_22419_, _14493_, _07659_);
  or (_22420_, _22419_, _22413_);
  and (_22421_, _22420_, _06102_);
  nor (_22422_, _06938_, _22409_);
  and (_22424_, _07659_, \oc8051_golden_model_1.ACC [2]);
  nor (_22425_, _22424_, _22413_);
  nor (_22426_, _22425_, _06939_);
  or (_22427_, _22426_, _22422_);
  and (_22428_, _22427_, _06954_);
  or (_22429_, _22428_, _06239_);
  or (_22430_, _22429_, _22421_);
  nand (_22431_, _22417_, _06239_);
  and (_22432_, _22431_, _06220_);
  nand (_22433_, _22432_, _22430_);
  or (_22435_, _22425_, _06220_);
  and (_22436_, _22435_, _09817_);
  nand (_22437_, _22436_, _22433_);
  and (_22438_, _22437_, _22418_);
  and (_22439_, _22438_, _22415_);
  or (_22440_, _22439_, _09833_);
  and (_22441_, _14580_, _07659_);
  or (_22442_, _22441_, _22413_);
  or (_22443_, _22442_, _05669_);
  and (_22444_, _22443_, _06020_);
  and (_22446_, _22444_, _22440_);
  and (_22447_, _07659_, _08730_);
  or (_22448_, _22447_, _22413_);
  and (_22449_, _22448_, _06019_);
  or (_22450_, _22449_, _06112_);
  or (_22451_, _22450_, _22446_);
  and (_22452_, _14596_, _07659_);
  or (_22453_, _22413_, _08751_);
  or (_22454_, _22453_, _22452_);
  and (_22455_, _22454_, _08756_);
  and (_22457_, _22455_, _22451_);
  and (_22458_, _10991_, _07659_);
  or (_22459_, _22458_, _22413_);
  and (_22460_, _22459_, _06284_);
  or (_22461_, _22460_, _22457_);
  and (_22462_, _22461_, _07032_);
  or (_22463_, _22413_, _08177_);
  and (_22464_, _22448_, _06108_);
  and (_22465_, _22464_, _22463_);
  or (_22466_, _22465_, _22462_);
  and (_22468_, _22466_, _06278_);
  nor (_22469_, _22425_, _06278_);
  and (_22470_, _22469_, _22463_);
  or (_22471_, _22470_, _06130_);
  or (_22472_, _22471_, _22468_);
  and (_22473_, _14593_, _07659_);
  or (_22474_, _22413_, _08777_);
  or (_22475_, _22474_, _22473_);
  and (_22476_, _22475_, _08782_);
  and (_22477_, _22476_, _22472_);
  nor (_22479_, _10990_, _11528_);
  or (_22480_, _22479_, _22413_);
  and (_22481_, _22480_, _06292_);
  or (_22482_, _22481_, _22477_);
  and (_22483_, _22482_, _06718_);
  and (_22484_, _22420_, _06316_);
  or (_22485_, _22484_, _06047_);
  or (_22486_, _22485_, _22483_);
  and (_22487_, _14657_, _07659_);
  or (_22488_, _22413_, _06048_);
  or (_22490_, _22488_, _22487_);
  and (_22491_, _22490_, _01336_);
  and (_22492_, _22491_, _22486_);
  or (_22493_, _22492_, _22410_);
  and (_43385_, _22493_, _42882_);
  not (_22494_, \oc8051_golden_model_1.TL0 [3]);
  nor (_22495_, _01336_, _22494_);
  and (_22496_, _09181_, _07659_);
  nor (_22497_, _07659_, _22494_);
  or (_22498_, _22497_, _07012_);
  or (_22500_, _22498_, _22496_);
  nor (_22501_, _11528_, _07353_);
  nor (_22502_, _22501_, _22497_);
  nand (_22503_, _22502_, _09815_);
  and (_22504_, _14672_, _07659_);
  or (_22505_, _22504_, _22497_);
  or (_22506_, _22505_, _06954_);
  and (_22507_, _07659_, \oc8051_golden_model_1.ACC [3]);
  nor (_22508_, _22507_, _22497_);
  nor (_22509_, _22508_, _06939_);
  nor (_22511_, _06938_, _22494_);
  or (_22512_, _22511_, _06102_);
  or (_22513_, _22512_, _22509_);
  and (_22514_, _22513_, _06848_);
  and (_22515_, _22514_, _22506_);
  nor (_22516_, _22502_, _06848_);
  or (_22517_, _22516_, _22515_);
  nand (_22518_, _22517_, _06220_);
  or (_22519_, _22508_, _06220_);
  and (_22520_, _22519_, _09817_);
  nand (_22522_, _22520_, _22518_);
  and (_22523_, _22522_, _22503_);
  and (_22524_, _22523_, _22500_);
  or (_22525_, _22524_, _09833_);
  and (_22526_, _14778_, _07659_);
  or (_22527_, _22526_, _22497_);
  or (_22528_, _22527_, _05669_);
  and (_22529_, _22528_, _06020_);
  and (_22530_, _22529_, _22525_);
  and (_22531_, _07659_, _08662_);
  or (_22533_, _22531_, _22497_);
  and (_22534_, _22533_, _06019_);
  or (_22535_, _22534_, _06112_);
  or (_22536_, _22535_, _22530_);
  and (_22537_, _14793_, _07659_);
  or (_22538_, _22537_, _22497_);
  or (_22539_, _22538_, _08751_);
  and (_22540_, _22539_, _08756_);
  and (_22541_, _22540_, _22536_);
  and (_22542_, _12299_, _07659_);
  or (_22544_, _22542_, _22497_);
  and (_22545_, _22544_, _06284_);
  or (_22546_, _22545_, _22541_);
  and (_22547_, _22546_, _07032_);
  or (_22548_, _22497_, _08029_);
  and (_22549_, _22533_, _06108_);
  and (_22550_, _22549_, _22548_);
  or (_22551_, _22550_, _22547_);
  and (_22552_, _22551_, _06278_);
  nor (_22553_, _22508_, _06278_);
  and (_22555_, _22553_, _22548_);
  or (_22556_, _22555_, _06130_);
  or (_22557_, _22556_, _22552_);
  and (_22558_, _14792_, _07659_);
  or (_22559_, _22497_, _08777_);
  or (_22560_, _22559_, _22558_);
  and (_22561_, _22560_, _08782_);
  and (_22562_, _22561_, _22557_);
  nor (_22563_, _10988_, _11528_);
  or (_22564_, _22563_, _22497_);
  and (_22566_, _22564_, _06292_);
  or (_22567_, _22566_, _22562_);
  and (_22568_, _22567_, _06718_);
  and (_22569_, _22505_, _06316_);
  or (_22570_, _22569_, _06047_);
  or (_22571_, _22570_, _22568_);
  and (_22572_, _14849_, _07659_);
  or (_22573_, _22497_, _06048_);
  or (_22574_, _22573_, _22572_);
  and (_22575_, _22574_, _01336_);
  and (_22577_, _22575_, _22571_);
  or (_22578_, _22577_, _22495_);
  and (_43386_, _22578_, _42882_);
  and (_22579_, _01340_, \oc8051_golden_model_1.TL0 [4]);
  and (_22580_, _11528_, \oc8051_golden_model_1.TL0 [4]);
  or (_22581_, _22580_, _08273_);
  and (_22582_, _08665_, _07659_);
  or (_22583_, _22582_, _22580_);
  and (_22584_, _22583_, _06108_);
  and (_22585_, _22584_, _22581_);
  or (_22587_, _22583_, _06020_);
  and (_22588_, _14887_, _07659_);
  or (_22589_, _22588_, _22580_);
  or (_22590_, _22589_, _06954_);
  and (_22591_, _07659_, \oc8051_golden_model_1.ACC [4]);
  or (_22592_, _22591_, _22580_);
  and (_22593_, _22592_, _06938_);
  and (_22594_, _06939_, \oc8051_golden_model_1.TL0 [4]);
  or (_22595_, _22594_, _06102_);
  or (_22596_, _22595_, _22593_);
  and (_22597_, _22596_, _06848_);
  and (_22598_, _22597_, _22590_);
  nor (_22599_, _08270_, _11528_);
  or (_22600_, _22599_, _22580_);
  and (_22601_, _22600_, _06239_);
  or (_22602_, _22601_, _22598_);
  and (_22603_, _22602_, _06220_);
  and (_22604_, _22592_, _06219_);
  or (_22605_, _22604_, _09818_);
  or (_22606_, _22605_, _22603_);
  and (_22609_, _09180_, _07659_);
  or (_22610_, _22580_, _07012_);
  or (_22611_, _22610_, _22609_);
  or (_22612_, _22600_, _09827_);
  and (_22613_, _22612_, _05669_);
  and (_22614_, _22613_, _22611_);
  and (_22615_, _22614_, _22606_);
  and (_22616_, _14983_, _07659_);
  or (_22617_, _22616_, _22580_);
  and (_22618_, _22617_, _09833_);
  or (_22620_, _22618_, _06019_);
  or (_22621_, _22620_, _22615_);
  and (_22622_, _22621_, _22587_);
  or (_22623_, _22622_, _06112_);
  and (_22624_, _14876_, _07659_);
  or (_22625_, _22580_, _08751_);
  or (_22626_, _22625_, _22624_);
  and (_22627_, _22626_, _08756_);
  and (_22628_, _22627_, _22623_);
  and (_22629_, _10986_, _07659_);
  or (_22631_, _22629_, _22580_);
  and (_22632_, _22631_, _06284_);
  or (_22633_, _22632_, _22628_);
  and (_22634_, _22633_, _07032_);
  or (_22635_, _22634_, _22585_);
  and (_22636_, _22635_, _06278_);
  and (_22637_, _22592_, _06277_);
  and (_22638_, _22637_, _22581_);
  or (_22639_, _22638_, _06130_);
  or (_22640_, _22639_, _22636_);
  and (_22642_, _14873_, _07659_);
  or (_22643_, _22580_, _08777_);
  or (_22644_, _22643_, _22642_);
  and (_22645_, _22644_, _08782_);
  and (_22646_, _22645_, _22640_);
  nor (_22647_, _10985_, _11528_);
  or (_22648_, _22647_, _22580_);
  and (_22649_, _22648_, _06292_);
  or (_22650_, _22649_, _22646_);
  and (_22651_, _22650_, _06718_);
  and (_22653_, _22589_, _06316_);
  or (_22654_, _22653_, _06047_);
  or (_22655_, _22654_, _22651_);
  and (_22656_, _15055_, _07659_);
  or (_22657_, _22580_, _06048_);
  or (_22658_, _22657_, _22656_);
  and (_22659_, _22658_, _01336_);
  and (_22660_, _22659_, _22655_);
  or (_22661_, _22660_, _22579_);
  and (_43387_, _22661_, _42882_);
  and (_22663_, _01340_, \oc8051_golden_model_1.TL0 [5]);
  and (_22664_, _11528_, \oc8051_golden_model_1.TL0 [5]);
  or (_22665_, _22664_, _07980_);
  and (_22666_, _08652_, _07659_);
  or (_22667_, _22666_, _22664_);
  and (_22668_, _22667_, _06108_);
  and (_22669_, _22668_, _22665_);
  or (_22670_, _22667_, _06020_);
  and (_22671_, _15093_, _07659_);
  or (_22672_, _22671_, _22664_);
  or (_22674_, _22672_, _06954_);
  and (_22675_, _07659_, \oc8051_golden_model_1.ACC [5]);
  or (_22676_, _22675_, _22664_);
  and (_22677_, _22676_, _06938_);
  and (_22678_, _06939_, \oc8051_golden_model_1.TL0 [5]);
  or (_22679_, _22678_, _06102_);
  or (_22680_, _22679_, _22677_);
  and (_22681_, _22680_, _06848_);
  and (_22682_, _22681_, _22674_);
  nor (_22683_, _07977_, _11528_);
  or (_22685_, _22683_, _22664_);
  and (_22686_, _22685_, _06239_);
  or (_22687_, _22686_, _22682_);
  and (_22688_, _22687_, _06220_);
  and (_22689_, _22676_, _06219_);
  or (_22690_, _22689_, _09818_);
  or (_22691_, _22690_, _22688_);
  and (_22692_, _09179_, _07659_);
  or (_22693_, _22664_, _07012_);
  or (_22694_, _22693_, _22692_);
  or (_22696_, _22685_, _09827_);
  and (_22697_, _22696_, _05669_);
  and (_22698_, _22697_, _22694_);
  and (_22699_, _22698_, _22691_);
  and (_22700_, _15179_, _07659_);
  or (_22701_, _22700_, _22664_);
  and (_22702_, _22701_, _09833_);
  or (_22703_, _22702_, _06019_);
  or (_22704_, _22703_, _22699_);
  and (_22705_, _22704_, _22670_);
  or (_22706_, _22705_, _06112_);
  and (_22707_, _15195_, _07659_);
  or (_22708_, _22707_, _22664_);
  or (_22709_, _22708_, _08751_);
  and (_22710_, _22709_, _08756_);
  and (_22711_, _22710_, _22706_);
  and (_22712_, _12306_, _07659_);
  or (_22713_, _22712_, _22664_);
  and (_22714_, _22713_, _06284_);
  or (_22715_, _22714_, _22711_);
  and (_22718_, _22715_, _07032_);
  or (_22719_, _22718_, _22669_);
  and (_22720_, _22719_, _06278_);
  and (_22721_, _22676_, _06277_);
  and (_22722_, _22721_, _22665_);
  or (_22723_, _22722_, _06130_);
  or (_22724_, _22723_, _22720_);
  and (_22725_, _15194_, _07659_);
  or (_22726_, _22664_, _08777_);
  or (_22727_, _22726_, _22725_);
  and (_22729_, _22727_, _08782_);
  and (_22730_, _22729_, _22724_);
  nor (_22731_, _10982_, _11528_);
  or (_22732_, _22731_, _22664_);
  and (_22733_, _22732_, _06292_);
  or (_22734_, _22733_, _22730_);
  and (_22735_, _22734_, _06718_);
  and (_22736_, _22672_, _06316_);
  or (_22737_, _22736_, _06047_);
  or (_22738_, _22737_, _22735_);
  and (_22740_, _15253_, _07659_);
  or (_22741_, _22664_, _06048_);
  or (_22742_, _22741_, _22740_);
  and (_22743_, _22742_, _01336_);
  and (_22744_, _22743_, _22738_);
  or (_22745_, _22744_, _22663_);
  and (_43388_, _22745_, _42882_);
  and (_22746_, _01340_, \oc8051_golden_model_1.TL0 [6]);
  and (_22747_, _11528_, \oc8051_golden_model_1.TL0 [6]);
  or (_22748_, _22747_, _07886_);
  and (_22750_, _15389_, _07659_);
  or (_22751_, _22750_, _22747_);
  and (_22752_, _22751_, _06108_);
  and (_22753_, _22752_, _22748_);
  or (_22754_, _22751_, _06020_);
  and (_22755_, _15293_, _07659_);
  or (_22756_, _22755_, _22747_);
  or (_22757_, _22756_, _06954_);
  and (_22758_, _07659_, \oc8051_golden_model_1.ACC [6]);
  or (_22759_, _22758_, _22747_);
  and (_22761_, _22759_, _06938_);
  and (_22762_, _06939_, \oc8051_golden_model_1.TL0 [6]);
  or (_22763_, _22762_, _06102_);
  or (_22764_, _22763_, _22761_);
  and (_22765_, _22764_, _06848_);
  and (_22766_, _22765_, _22757_);
  nor (_22767_, _07883_, _11528_);
  or (_22768_, _22767_, _22747_);
  and (_22769_, _22768_, _06239_);
  or (_22770_, _22769_, _22766_);
  and (_22772_, _22770_, _06220_);
  and (_22773_, _22759_, _06219_);
  or (_22774_, _22773_, _09818_);
  or (_22775_, _22774_, _22772_);
  and (_22776_, _09178_, _07659_);
  or (_22777_, _22747_, _07012_);
  or (_22778_, _22777_, _22776_);
  or (_22779_, _22768_, _09827_);
  and (_22780_, _22779_, _05669_);
  and (_22781_, _22780_, _22778_);
  and (_22783_, _22781_, _22775_);
  and (_22784_, _15382_, _07659_);
  or (_22785_, _22784_, _22747_);
  and (_22786_, _22785_, _09833_);
  or (_22787_, _22786_, _06019_);
  or (_22788_, _22787_, _22783_);
  and (_22789_, _22788_, _22754_);
  or (_22790_, _22789_, _06112_);
  and (_22791_, _15399_, _07659_);
  or (_22792_, _22747_, _08751_);
  or (_22794_, _22792_, _22791_);
  and (_22795_, _22794_, _08756_);
  and (_22796_, _22795_, _22790_);
  and (_22797_, _10980_, _07659_);
  or (_22798_, _22797_, _22747_);
  and (_22799_, _22798_, _06284_);
  or (_22800_, _22799_, _22796_);
  and (_22801_, _22800_, _07032_);
  or (_22802_, _22801_, _22753_);
  and (_22803_, _22802_, _06278_);
  and (_22805_, _22759_, _06277_);
  and (_22806_, _22805_, _22748_);
  or (_22807_, _22806_, _06130_);
  or (_22808_, _22807_, _22803_);
  and (_22809_, _15396_, _07659_);
  or (_22810_, _22747_, _08777_);
  or (_22811_, _22810_, _22809_);
  and (_22812_, _22811_, _08782_);
  and (_22813_, _22812_, _22808_);
  nor (_22814_, _10979_, _11528_);
  or (_22816_, _22814_, _22747_);
  and (_22817_, _22816_, _06292_);
  or (_22818_, _22817_, _22813_);
  and (_22819_, _22818_, _06718_);
  and (_22820_, _22756_, _06316_);
  or (_22821_, _22820_, _06047_);
  or (_22822_, _22821_, _22819_);
  and (_22823_, _15451_, _07659_);
  or (_22824_, _22747_, _06048_);
  or (_22825_, _22824_, _22823_);
  and (_22827_, _22825_, _01336_);
  and (_22828_, _22827_, _22822_);
  or (_22829_, _22828_, _22746_);
  and (_43389_, _22829_, _42882_);
  not (_22830_, \oc8051_golden_model_1.TCON [0]);
  nor (_22831_, _01336_, _22830_);
  nand (_22832_, _10995_, _07648_);
  nor (_22833_, _07648_, _22830_);
  nor (_22834_, _22833_, _06278_);
  nand (_22835_, _22834_, _22832_);
  and (_22837_, _07648_, _08672_);
  or (_22838_, _22837_, _22833_);
  or (_22839_, _22838_, _06020_);
  and (_22840_, _09120_, _07648_);
  or (_22841_, _22833_, _07012_);
  or (_22842_, _22841_, _22840_);
  nor (_22843_, _08127_, _11605_);
  or (_22844_, _22843_, _22833_);
  or (_22845_, _22844_, _06954_);
  and (_22846_, _07648_, \oc8051_golden_model_1.ACC [0]);
  or (_22848_, _22846_, _22833_);
  and (_22849_, _22848_, _06938_);
  nor (_22850_, _06938_, _22830_);
  or (_22851_, _22850_, _06102_);
  or (_22852_, _22851_, _22849_);
  and (_22853_, _22852_, _06044_);
  and (_22854_, _22853_, _22845_);
  nor (_22855_, _08341_, _22830_);
  and (_22856_, _14102_, _08341_);
  or (_22857_, _22856_, _22855_);
  and (_22859_, _22857_, _06043_);
  or (_22860_, _22859_, _22854_);
  and (_22861_, _22860_, _06848_);
  and (_22862_, _07648_, _06931_);
  or (_22863_, _22862_, _22833_);
  and (_22864_, _22863_, _06239_);
  or (_22865_, _22864_, _06219_);
  or (_22866_, _22865_, _22861_);
  or (_22867_, _22848_, _06220_);
  and (_22868_, _22867_, _06040_);
  and (_22870_, _22868_, _22866_);
  and (_22871_, _22833_, _06039_);
  or (_22872_, _22871_, _06032_);
  or (_22873_, _22872_, _22870_);
  or (_22874_, _22844_, _06033_);
  and (_22875_, _22874_, _06027_);
  and (_22876_, _22875_, _22873_);
  or (_22877_, _22855_, _14131_);
  and (_22878_, _22877_, _06026_);
  and (_22879_, _22878_, _22857_);
  or (_22881_, _22879_, _09818_);
  or (_22882_, _22881_, _22876_);
  or (_22883_, _22863_, _09827_);
  and (_22884_, _22883_, _05669_);
  and (_22885_, _22884_, _22882_);
  and (_22886_, _22885_, _22842_);
  and (_22887_, _14186_, _07648_);
  or (_22888_, _22887_, _22833_);
  and (_22889_, _22888_, _09833_);
  or (_22890_, _22889_, _06019_);
  or (_22892_, _22890_, _22886_);
  and (_22893_, _22892_, _22839_);
  or (_22894_, _22893_, _06112_);
  and (_22895_, _14086_, _07648_);
  or (_22896_, _22833_, _08751_);
  or (_22897_, _22896_, _22895_);
  and (_22898_, _22897_, _08756_);
  and (_22899_, _22898_, _22894_);
  nor (_22900_, _12302_, _11605_);
  or (_22901_, _22900_, _22833_);
  and (_22903_, _22832_, _06284_);
  and (_22904_, _22903_, _22901_);
  or (_22905_, _22904_, _22899_);
  and (_22906_, _22905_, _07032_);
  nand (_22907_, _22838_, _06108_);
  nor (_22908_, _22907_, _22843_);
  or (_22909_, _22908_, _06277_);
  or (_22910_, _22909_, _22906_);
  and (_22911_, _22910_, _22835_);
  or (_22912_, _22911_, _06130_);
  and (_22914_, _14083_, _07648_);
  or (_22915_, _22833_, _08777_);
  or (_22916_, _22915_, _22914_);
  and (_22917_, _22916_, _08782_);
  and (_22918_, _22917_, _22912_);
  and (_22919_, _22901_, _06292_);
  or (_22920_, _22919_, _06316_);
  or (_22921_, _22920_, _22918_);
  or (_22922_, _22844_, _06718_);
  and (_22923_, _22922_, _22921_);
  or (_22924_, _22923_, _05652_);
  or (_22925_, _22833_, _05653_);
  and (_22926_, _22925_, _22924_);
  or (_22927_, _22926_, _06047_);
  or (_22928_, _22844_, _06048_);
  and (_22929_, _22928_, _01336_);
  and (_22930_, _22929_, _22927_);
  or (_22931_, _22930_, _22831_);
  and (_43391_, _22931_, _42882_);
  and (_22932_, _01340_, \oc8051_golden_model_1.TCON [1]);
  and (_22935_, _11605_, \oc8051_golden_model_1.TCON [1]);
  nor (_22936_, _10993_, _11605_);
  or (_22937_, _22936_, _22935_);
  or (_22938_, _22937_, _08782_);
  or (_22939_, _14367_, _11605_);
  or (_22940_, _07648_, \oc8051_golden_model_1.TCON [1]);
  and (_22941_, _22940_, _09833_);
  and (_22942_, _22941_, _22939_);
  nor (_22943_, _11605_, _07132_);
  or (_22944_, _22943_, _22935_);
  or (_22946_, _22944_, _06848_);
  and (_22947_, _14284_, _07648_);
  not (_22948_, _22947_);
  and (_22949_, _22948_, _22940_);
  or (_22950_, _22949_, _06954_);
  and (_22951_, _07648_, \oc8051_golden_model_1.ACC [1]);
  or (_22952_, _22951_, _22935_);
  and (_22953_, _22952_, _06938_);
  and (_22954_, _06939_, \oc8051_golden_model_1.TCON [1]);
  or (_22955_, _22954_, _06102_);
  or (_22957_, _22955_, _22953_);
  and (_22958_, _22957_, _06044_);
  and (_22959_, _22958_, _22950_);
  and (_22960_, _11624_, \oc8051_golden_model_1.TCON [1]);
  and (_22961_, _14266_, _08341_);
  or (_22962_, _22961_, _22960_);
  and (_22963_, _22962_, _06043_);
  or (_22964_, _22963_, _06239_);
  or (_22965_, _22964_, _22959_);
  and (_22966_, _22965_, _22946_);
  or (_22968_, _22966_, _06219_);
  or (_22969_, _22952_, _06220_);
  and (_22970_, _22969_, _06040_);
  and (_22971_, _22970_, _22968_);
  and (_22972_, _14273_, _08341_);
  or (_22973_, _22972_, _22960_);
  and (_22974_, _22973_, _06039_);
  or (_22975_, _22974_, _06032_);
  or (_22976_, _22975_, _22971_);
  and (_22977_, _22961_, _14302_);
  or (_22979_, _22960_, _06033_);
  or (_22980_, _22979_, _22977_);
  and (_22981_, _22980_, _06027_);
  and (_22982_, _22981_, _22976_);
  or (_22983_, _22960_, _14267_);
  and (_22984_, _22983_, _06026_);
  and (_22985_, _22984_, _22962_);
  or (_22986_, _22985_, _09818_);
  or (_22987_, _22986_, _22982_);
  and (_22988_, _09075_, _07648_);
  or (_22990_, _22935_, _07012_);
  or (_22991_, _22990_, _22988_);
  or (_22992_, _22944_, _09827_);
  and (_22993_, _22992_, _05669_);
  and (_22994_, _22993_, _22991_);
  and (_22995_, _22994_, _22987_);
  or (_22996_, _22995_, _22942_);
  and (_22997_, _22996_, _06020_);
  nand (_22998_, _07648_, _06832_);
  and (_22999_, _22940_, _06019_);
  and (_23001_, _22999_, _22998_);
  or (_23002_, _23001_, _22997_);
  and (_23003_, _23002_, _08751_);
  or (_23004_, _14263_, _11605_);
  and (_23005_, _22940_, _06112_);
  and (_23006_, _23005_, _23004_);
  or (_23007_, _23006_, _06284_);
  or (_23008_, _23007_, _23003_);
  and (_23009_, _10994_, _07648_);
  or (_23010_, _23009_, _22935_);
  or (_23012_, _23010_, _08756_);
  and (_23013_, _23012_, _07032_);
  and (_23014_, _23013_, _23008_);
  or (_23015_, _14261_, _11605_);
  and (_23016_, _22940_, _06108_);
  and (_23017_, _23016_, _23015_);
  or (_23018_, _23017_, _06277_);
  or (_23019_, _23018_, _23014_);
  and (_23020_, _22951_, _08078_);
  or (_23021_, _22935_, _06278_);
  or (_23023_, _23021_, _23020_);
  and (_23024_, _23023_, _08777_);
  and (_23025_, _23024_, _23019_);
  or (_23026_, _22998_, _08078_);
  and (_23027_, _22940_, _06130_);
  and (_23028_, _23027_, _23026_);
  or (_23029_, _23028_, _06292_);
  or (_23030_, _23029_, _23025_);
  and (_23031_, _23030_, _22938_);
  or (_23032_, _23031_, _06316_);
  or (_23034_, _22949_, _06718_);
  and (_23035_, _23034_, _05653_);
  and (_23036_, _23035_, _23032_);
  and (_23037_, _22973_, _05652_);
  or (_23038_, _23037_, _06047_);
  or (_23039_, _23038_, _23036_);
  or (_23040_, _22935_, _06048_);
  or (_23041_, _23040_, _22947_);
  and (_23042_, _23041_, _01336_);
  and (_23043_, _23042_, _23039_);
  or (_23044_, _23043_, _22932_);
  and (_43392_, _23044_, _42882_);
  and (_23045_, _01340_, \oc8051_golden_model_1.TCON [2]);
  and (_23046_, _11605_, \oc8051_golden_model_1.TCON [2]);
  and (_23047_, _07648_, _08730_);
  or (_23048_, _23047_, _23046_);
  or (_23049_, _23048_, _06020_);
  nor (_23050_, _11605_, _07530_);
  or (_23051_, _23050_, _23046_);
  and (_23052_, _23051_, _06239_);
  and (_23054_, _11624_, \oc8051_golden_model_1.TCON [2]);
  and (_23055_, _14497_, _08341_);
  or (_23056_, _23055_, _23054_);
  or (_23057_, _23056_, _06044_);
  and (_23058_, _14493_, _07648_);
  or (_23059_, _23058_, _23046_);
  and (_23060_, _23059_, _06102_);
  and (_23061_, _06939_, \oc8051_golden_model_1.TCON [2]);
  and (_23062_, _07648_, \oc8051_golden_model_1.ACC [2]);
  or (_23063_, _23062_, _23046_);
  and (_23065_, _23063_, _06938_);
  or (_23066_, _23065_, _23061_);
  and (_23067_, _23066_, _06954_);
  or (_23068_, _23067_, _06043_);
  or (_23069_, _23068_, _23060_);
  and (_23070_, _23069_, _23057_);
  and (_23071_, _23070_, _06848_);
  or (_23072_, _23071_, _23052_);
  or (_23073_, _23072_, _06219_);
  or (_23074_, _23063_, _06220_);
  and (_23076_, _23074_, _06040_);
  and (_23077_, _23076_, _23073_);
  and (_23078_, _14479_, _08341_);
  or (_23079_, _23078_, _23054_);
  and (_23080_, _23079_, _06039_);
  or (_23081_, _23080_, _06032_);
  or (_23082_, _23081_, _23077_);
  or (_23083_, _23054_, _14512_);
  and (_23084_, _23083_, _23056_);
  or (_23085_, _23084_, _06033_);
  and (_23086_, _23085_, _06027_);
  and (_23087_, _23086_, _23082_);
  or (_23088_, _23054_, _14525_);
  and (_23089_, _23088_, _06026_);
  and (_23090_, _23089_, _23056_);
  or (_23091_, _23090_, _09818_);
  or (_23092_, _23091_, _23087_);
  and (_23093_, _09182_, _07648_);
  or (_23094_, _23046_, _07012_);
  or (_23095_, _23094_, _23093_);
  or (_23097_, _23051_, _09827_);
  and (_23098_, _23097_, _05669_);
  and (_23099_, _23098_, _23095_);
  and (_23100_, _23099_, _23092_);
  and (_23101_, _14580_, _07648_);
  or (_23102_, _23101_, _23046_);
  and (_23103_, _23102_, _09833_);
  or (_23104_, _23103_, _06019_);
  or (_23105_, _23104_, _23100_);
  and (_23106_, _23105_, _23049_);
  or (_23107_, _23106_, _06112_);
  and (_23108_, _14596_, _07648_);
  or (_23109_, _23108_, _23046_);
  or (_23110_, _23109_, _08751_);
  and (_23111_, _23110_, _08756_);
  and (_23112_, _23111_, _23107_);
  and (_23113_, _10991_, _07648_);
  or (_23114_, _23113_, _23046_);
  and (_23115_, _23114_, _06284_);
  or (_23116_, _23115_, _23112_);
  and (_23118_, _23116_, _07032_);
  or (_23119_, _23046_, _08177_);
  and (_23120_, _23048_, _06108_);
  and (_23121_, _23120_, _23119_);
  or (_23122_, _23121_, _23118_);
  and (_23123_, _23122_, _06278_);
  and (_23124_, _23063_, _06277_);
  and (_23125_, _23124_, _23119_);
  or (_23126_, _23125_, _06130_);
  or (_23127_, _23126_, _23123_);
  and (_23129_, _14593_, _07648_);
  or (_23130_, _23046_, _08777_);
  or (_23131_, _23130_, _23129_);
  and (_23132_, _23131_, _08782_);
  and (_23133_, _23132_, _23127_);
  nor (_23134_, _10990_, _11605_);
  or (_23135_, _23134_, _23046_);
  and (_23136_, _23135_, _06292_);
  or (_23137_, _23136_, _06316_);
  or (_23138_, _23137_, _23133_);
  or (_23139_, _23059_, _06718_);
  and (_23140_, _23139_, _05653_);
  and (_23141_, _23140_, _23138_);
  and (_23142_, _23079_, _05652_);
  or (_23143_, _23142_, _06047_);
  or (_23144_, _23143_, _23141_);
  and (_23145_, _14657_, _07648_);
  or (_23146_, _23046_, _06048_);
  or (_23147_, _23146_, _23145_);
  and (_23148_, _23147_, _01336_);
  and (_23150_, _23148_, _23144_);
  or (_23151_, _23150_, _23045_);
  and (_43393_, _23151_, _42882_);
  and (_23152_, _01340_, \oc8051_golden_model_1.TCON [3]);
  and (_23153_, _11605_, \oc8051_golden_model_1.TCON [3]);
  and (_23154_, _07648_, _08662_);
  or (_23155_, _23154_, _23153_);
  or (_23156_, _23155_, _06020_);
  and (_23157_, _14672_, _07648_);
  or (_23158_, _23157_, _23153_);
  or (_23160_, _23158_, _06954_);
  and (_23161_, _07648_, \oc8051_golden_model_1.ACC [3]);
  or (_23162_, _23161_, _23153_);
  and (_23163_, _23162_, _06938_);
  and (_23164_, _06939_, \oc8051_golden_model_1.TCON [3]);
  or (_23165_, _23164_, _06102_);
  or (_23166_, _23165_, _23163_);
  and (_23167_, _23166_, _06044_);
  and (_23168_, _23167_, _23160_);
  and (_23169_, _11624_, \oc8051_golden_model_1.TCON [3]);
  and (_23170_, _14683_, _08341_);
  or (_23171_, _23170_, _23169_);
  and (_23172_, _23171_, _06043_);
  or (_23173_, _23172_, _06239_);
  or (_23174_, _23173_, _23168_);
  nor (_23175_, _11605_, _07353_);
  or (_23176_, _23175_, _23153_);
  or (_23177_, _23176_, _06848_);
  and (_23178_, _23177_, _23174_);
  or (_23179_, _23178_, _06219_);
  or (_23180_, _23162_, _06220_);
  and (_23181_, _23180_, _06040_);
  and (_23182_, _23181_, _23179_);
  and (_23183_, _14681_, _08341_);
  or (_23184_, _23183_, _23169_);
  and (_23185_, _23184_, _06039_);
  or (_23186_, _23185_, _06032_);
  or (_23187_, _23186_, _23182_);
  or (_23188_, _23169_, _14708_);
  and (_23189_, _23188_, _23171_);
  or (_23192_, _23189_, _06033_);
  and (_23193_, _23192_, _06027_);
  and (_23194_, _23193_, _23187_);
  and (_23195_, _14724_, _08341_);
  or (_23196_, _23195_, _23169_);
  and (_23197_, _23196_, _06026_);
  or (_23198_, _23197_, _09818_);
  or (_23199_, _23198_, _23194_);
  and (_23200_, _09181_, _07648_);
  or (_23201_, _23153_, _07012_);
  or (_23202_, _23201_, _23200_);
  or (_23203_, _23176_, _09827_);
  and (_23204_, _23203_, _05669_);
  and (_23205_, _23204_, _23202_);
  and (_23206_, _23205_, _23199_);
  and (_23207_, _14778_, _07648_);
  or (_23208_, _23207_, _23153_);
  and (_23209_, _23208_, _09833_);
  or (_23210_, _23209_, _06019_);
  or (_23211_, _23210_, _23206_);
  and (_23213_, _23211_, _23156_);
  or (_23214_, _23213_, _06112_);
  and (_23215_, _14793_, _07648_);
  or (_23216_, _23153_, _08751_);
  or (_23217_, _23216_, _23215_);
  and (_23218_, _23217_, _08756_);
  and (_23219_, _23218_, _23214_);
  and (_23220_, _12299_, _07648_);
  or (_23221_, _23220_, _23153_);
  and (_23222_, _23221_, _06284_);
  or (_23224_, _23222_, _23219_);
  and (_23225_, _23224_, _07032_);
  or (_23226_, _23153_, _08029_);
  and (_23227_, _23155_, _06108_);
  and (_23228_, _23227_, _23226_);
  or (_23229_, _23228_, _23225_);
  and (_23230_, _23229_, _06278_);
  and (_23231_, _23162_, _06277_);
  and (_23232_, _23231_, _23226_);
  or (_23233_, _23232_, _06130_);
  or (_23234_, _23233_, _23230_);
  and (_23235_, _14792_, _07648_);
  or (_23236_, _23153_, _08777_);
  or (_23237_, _23236_, _23235_);
  and (_23238_, _23237_, _08782_);
  and (_23239_, _23238_, _23234_);
  nor (_23240_, _10988_, _11605_);
  or (_23241_, _23240_, _23153_);
  and (_23242_, _23241_, _06292_);
  or (_23243_, _23242_, _06316_);
  or (_23245_, _23243_, _23239_);
  or (_23246_, _23158_, _06718_);
  and (_23247_, _23246_, _05653_);
  and (_23248_, _23247_, _23245_);
  and (_23249_, _23184_, _05652_);
  or (_23250_, _23249_, _06047_);
  or (_23251_, _23250_, _23248_);
  and (_23252_, _14849_, _07648_);
  or (_23253_, _23153_, _06048_);
  or (_23254_, _23253_, _23252_);
  and (_23256_, _23254_, _01336_);
  and (_23257_, _23256_, _23251_);
  or (_23258_, _23257_, _23152_);
  and (_43394_, _23258_, _42882_);
  and (_23259_, _01340_, \oc8051_golden_model_1.TCON [4]);
  and (_23260_, _11605_, \oc8051_golden_model_1.TCON [4]);
  and (_23261_, _08665_, _07648_);
  or (_23262_, _23261_, _23260_);
  or (_23263_, _23262_, _06020_);
  and (_23264_, _14887_, _07648_);
  or (_23265_, _23264_, _23260_);
  or (_23266_, _23265_, _06954_);
  and (_23267_, _07648_, \oc8051_golden_model_1.ACC [4]);
  or (_23268_, _23267_, _23260_);
  and (_23269_, _23268_, _06938_);
  and (_23270_, _06939_, \oc8051_golden_model_1.TCON [4]);
  or (_23271_, _23270_, _06102_);
  or (_23272_, _23271_, _23269_);
  and (_23273_, _23272_, _06044_);
  and (_23274_, _23273_, _23266_);
  and (_23276_, _11624_, \oc8051_golden_model_1.TCON [4]);
  and (_23277_, _14878_, _08341_);
  or (_23278_, _23277_, _23276_);
  and (_23279_, _23278_, _06043_);
  or (_23280_, _23279_, _06239_);
  or (_23281_, _23280_, _23274_);
  nor (_23282_, _08270_, _11605_);
  or (_23283_, _23282_, _23260_);
  or (_23284_, _23283_, _06848_);
  and (_23285_, _23284_, _23281_);
  or (_23287_, _23285_, _06219_);
  or (_23288_, _23268_, _06220_);
  and (_23289_, _23288_, _06040_);
  and (_23290_, _23289_, _23287_);
  and (_23291_, _14882_, _08341_);
  or (_23292_, _23291_, _23276_);
  and (_23293_, _23292_, _06039_);
  or (_23294_, _23293_, _06032_);
  or (_23295_, _23294_, _23290_);
  or (_23296_, _23276_, _14914_);
  and (_23297_, _23296_, _23278_);
  or (_23298_, _23297_, _06033_);
  and (_23299_, _23298_, _06027_);
  and (_23300_, _23299_, _23295_);
  or (_23301_, _23276_, _14879_);
  and (_23302_, _23301_, _06026_);
  and (_23303_, _23302_, _23278_);
  or (_23304_, _23303_, _09818_);
  or (_23305_, _23304_, _23300_);
  and (_23306_, _09180_, _07648_);
  or (_23308_, _23260_, _07012_);
  or (_23309_, _23308_, _23306_);
  or (_23310_, _23283_, _09827_);
  and (_23311_, _23310_, _05669_);
  and (_23312_, _23311_, _23309_);
  and (_23313_, _23312_, _23305_);
  and (_23314_, _14983_, _07648_);
  or (_23315_, _23314_, _23260_);
  and (_23316_, _23315_, _09833_);
  or (_23317_, _23316_, _06019_);
  or (_23319_, _23317_, _23313_);
  and (_23320_, _23319_, _23263_);
  or (_23321_, _23320_, _06112_);
  and (_23322_, _14876_, _07648_);
  or (_23323_, _23260_, _08751_);
  or (_23324_, _23323_, _23322_);
  and (_23325_, _23324_, _08756_);
  and (_23326_, _23325_, _23321_);
  and (_23327_, _10986_, _07648_);
  or (_23328_, _23327_, _23260_);
  and (_23329_, _23328_, _06284_);
  or (_23330_, _23329_, _23326_);
  and (_23331_, _23330_, _07032_);
  or (_23332_, _23260_, _08273_);
  and (_23333_, _23262_, _06108_);
  and (_23334_, _23333_, _23332_);
  or (_23335_, _23334_, _23331_);
  and (_23336_, _23335_, _06278_);
  and (_23337_, _23268_, _06277_);
  and (_23338_, _23337_, _23332_);
  or (_23340_, _23338_, _06130_);
  or (_23341_, _23340_, _23336_);
  and (_23342_, _14873_, _07648_);
  or (_23343_, _23260_, _08777_);
  or (_23344_, _23343_, _23342_);
  and (_23345_, _23344_, _08782_);
  and (_23346_, _23345_, _23341_);
  nor (_23347_, _10985_, _11605_);
  or (_23348_, _23347_, _23260_);
  and (_23349_, _23348_, _06292_);
  or (_23351_, _23349_, _06316_);
  or (_23352_, _23351_, _23346_);
  or (_23353_, _23265_, _06718_);
  and (_23354_, _23353_, _05653_);
  and (_23355_, _23354_, _23352_);
  and (_23356_, _23292_, _05652_);
  or (_23357_, _23356_, _06047_);
  or (_23358_, _23357_, _23355_);
  and (_23359_, _15055_, _07648_);
  or (_23360_, _23260_, _06048_);
  or (_23361_, _23360_, _23359_);
  and (_23362_, _23361_, _01336_);
  and (_23363_, _23362_, _23358_);
  or (_23364_, _23363_, _23259_);
  and (_43395_, _23364_, _42882_);
  and (_23365_, _01340_, \oc8051_golden_model_1.TCON [5]);
  and (_23366_, _11605_, \oc8051_golden_model_1.TCON [5]);
  and (_23367_, _08652_, _07648_);
  or (_23368_, _23367_, _23366_);
  or (_23369_, _23368_, _06020_);
  and (_23371_, _15093_, _07648_);
  or (_23372_, _23371_, _23366_);
  or (_23373_, _23372_, _06954_);
  and (_23374_, _07648_, \oc8051_golden_model_1.ACC [5]);
  or (_23375_, _23374_, _23366_);
  and (_23376_, _23375_, _06938_);
  and (_23377_, _06939_, \oc8051_golden_model_1.TCON [5]);
  or (_23378_, _23377_, _06102_);
  or (_23379_, _23378_, _23376_);
  and (_23380_, _23379_, _06044_);
  and (_23382_, _23380_, _23373_);
  and (_23383_, _11624_, \oc8051_golden_model_1.TCON [5]);
  and (_23384_, _15073_, _08341_);
  or (_23385_, _23384_, _23383_);
  and (_23386_, _23385_, _06043_);
  or (_23387_, _23386_, _06239_);
  or (_23388_, _23387_, _23382_);
  nor (_23389_, _07977_, _11605_);
  or (_23390_, _23389_, _23366_);
  or (_23391_, _23390_, _06848_);
  and (_23392_, _23391_, _23388_);
  or (_23393_, _23392_, _06219_);
  or (_23394_, _23375_, _06220_);
  and (_23395_, _23394_, _06040_);
  and (_23396_, _23395_, _23393_);
  and (_23397_, _15077_, _08341_);
  or (_23398_, _23397_, _23383_);
  and (_23399_, _23398_, _06039_);
  or (_23400_, _23399_, _06032_);
  or (_23401_, _23400_, _23396_);
  or (_23403_, _23383_, _15110_);
  and (_23404_, _23403_, _23385_);
  or (_23405_, _23404_, _06033_);
  and (_23406_, _23405_, _06027_);
  and (_23407_, _23406_, _23401_);
  or (_23408_, _23383_, _15074_);
  and (_23409_, _23408_, _06026_);
  and (_23410_, _23409_, _23385_);
  or (_23411_, _23410_, _09818_);
  or (_23412_, _23411_, _23407_);
  and (_23414_, _09179_, _07648_);
  or (_23415_, _23366_, _07012_);
  or (_23416_, _23415_, _23414_);
  or (_23417_, _23390_, _09827_);
  and (_23418_, _23417_, _05669_);
  and (_23419_, _23418_, _23416_);
  and (_23420_, _23419_, _23412_);
  and (_23421_, _15179_, _07648_);
  or (_23422_, _23421_, _23366_);
  and (_23423_, _23422_, _09833_);
  or (_23424_, _23423_, _06019_);
  or (_23425_, _23424_, _23420_);
  and (_23426_, _23425_, _23369_);
  or (_23427_, _23426_, _06112_);
  and (_23428_, _15195_, _07648_);
  or (_23429_, _23428_, _23366_);
  or (_23430_, _23429_, _08751_);
  and (_23431_, _23430_, _08756_);
  and (_23432_, _23431_, _23427_);
  and (_23433_, _12306_, _07648_);
  or (_23435_, _23433_, _23366_);
  and (_23436_, _23435_, _06284_);
  or (_23437_, _23436_, _23432_);
  and (_23438_, _23437_, _07032_);
  or (_23439_, _23366_, _07980_);
  and (_23440_, _23368_, _06108_);
  and (_23441_, _23440_, _23439_);
  or (_23442_, _23441_, _23438_);
  and (_23443_, _23442_, _06278_);
  and (_23444_, _23375_, _06277_);
  and (_23446_, _23444_, _23439_);
  or (_23447_, _23446_, _06130_);
  or (_23448_, _23447_, _23443_);
  and (_23449_, _15194_, _07648_);
  or (_23450_, _23366_, _08777_);
  or (_23451_, _23450_, _23449_);
  and (_23452_, _23451_, _08782_);
  and (_23453_, _23452_, _23448_);
  nor (_23454_, _10982_, _11605_);
  or (_23455_, _23454_, _23366_);
  and (_23456_, _23455_, _06292_);
  or (_23457_, _23456_, _06316_);
  or (_23458_, _23457_, _23453_);
  or (_23459_, _23372_, _06718_);
  and (_23460_, _23459_, _05653_);
  and (_23461_, _23460_, _23458_);
  and (_23462_, _23398_, _05652_);
  or (_23463_, _23462_, _06047_);
  or (_23464_, _23463_, _23461_);
  and (_23465_, _15253_, _07648_);
  or (_23467_, _23366_, _06048_);
  or (_23468_, _23467_, _23465_);
  and (_23469_, _23468_, _01336_);
  and (_23470_, _23469_, _23464_);
  or (_23471_, _23470_, _23365_);
  and (_43396_, _23471_, _42882_);
  and (_23472_, _01340_, \oc8051_golden_model_1.TCON [6]);
  and (_23473_, _11605_, \oc8051_golden_model_1.TCON [6]);
  and (_23474_, _15389_, _07648_);
  or (_23475_, _23474_, _23473_);
  or (_23477_, _23475_, _06020_);
  and (_23478_, _15293_, _07648_);
  or (_23479_, _23478_, _23473_);
  or (_23480_, _23479_, _06954_);
  and (_23481_, _07648_, \oc8051_golden_model_1.ACC [6]);
  or (_23482_, _23481_, _23473_);
  and (_23483_, _23482_, _06938_);
  and (_23484_, _06939_, \oc8051_golden_model_1.TCON [6]);
  or (_23485_, _23484_, _06102_);
  or (_23486_, _23485_, _23483_);
  and (_23488_, _23486_, _06044_);
  and (_23489_, _23488_, _23480_);
  and (_23490_, _11624_, \oc8051_golden_model_1.TCON [6]);
  and (_23491_, _15280_, _08341_);
  or (_23492_, _23491_, _23490_);
  and (_23493_, _23492_, _06043_);
  or (_23494_, _23493_, _06239_);
  or (_23495_, _23494_, _23489_);
  nor (_23496_, _07883_, _11605_);
  or (_23497_, _23496_, _23473_);
  or (_23498_, _23497_, _06848_);
  and (_23499_, _23498_, _23495_);
  or (_23500_, _23499_, _06219_);
  or (_23501_, _23482_, _06220_);
  and (_23502_, _23501_, _06040_);
  and (_23503_, _23502_, _23500_);
  and (_23504_, _15278_, _08341_);
  or (_23505_, _23504_, _23490_);
  and (_23506_, _23505_, _06039_);
  or (_23507_, _23506_, _06032_);
  or (_23509_, _23507_, _23503_);
  or (_23510_, _23490_, _15310_);
  and (_23511_, _23510_, _23492_);
  or (_23512_, _23511_, _06033_);
  and (_23513_, _23512_, _06027_);
  and (_23514_, _23513_, _23509_);
  or (_23515_, _23490_, _15326_);
  and (_23516_, _23515_, _06026_);
  and (_23517_, _23516_, _23492_);
  or (_23518_, _23517_, _09818_);
  or (_23520_, _23518_, _23514_);
  and (_23521_, _09178_, _07648_);
  or (_23522_, _23473_, _07012_);
  or (_23523_, _23522_, _23521_);
  or (_23524_, _23497_, _09827_);
  and (_23525_, _23524_, _05669_);
  and (_23526_, _23525_, _23523_);
  and (_23527_, _23526_, _23520_);
  and (_23528_, _15382_, _07648_);
  or (_23529_, _23528_, _23473_);
  and (_23531_, _23529_, _09833_);
  or (_23532_, _23531_, _06019_);
  or (_23533_, _23532_, _23527_);
  and (_23534_, _23533_, _23477_);
  or (_23535_, _23534_, _06112_);
  and (_23536_, _15399_, _07648_);
  or (_23537_, _23473_, _08751_);
  or (_23538_, _23537_, _23536_);
  and (_23539_, _23538_, _08756_);
  and (_23540_, _23539_, _23535_);
  and (_23541_, _10980_, _07648_);
  or (_23542_, _23541_, _23473_);
  and (_23543_, _23542_, _06284_);
  or (_23544_, _23543_, _23540_);
  and (_23545_, _23544_, _07032_);
  or (_23546_, _23473_, _07886_);
  and (_23547_, _23475_, _06108_);
  and (_23548_, _23547_, _23546_);
  or (_23549_, _23548_, _23545_);
  and (_23550_, _23549_, _06278_);
  and (_23552_, _23482_, _06277_);
  and (_23553_, _23552_, _23546_);
  or (_23554_, _23553_, _06130_);
  or (_23555_, _23554_, _23550_);
  and (_23556_, _15396_, _07648_);
  or (_23557_, _23473_, _08777_);
  or (_23558_, _23557_, _23556_);
  and (_23559_, _23558_, _08782_);
  and (_23560_, _23559_, _23555_);
  nor (_23561_, _10979_, _11605_);
  or (_23563_, _23561_, _23473_);
  and (_23564_, _23563_, _06292_);
  or (_23565_, _23564_, _06316_);
  or (_23566_, _23565_, _23560_);
  or (_23567_, _23479_, _06718_);
  and (_23568_, _23567_, _05653_);
  and (_23569_, _23568_, _23566_);
  and (_23570_, _23505_, _05652_);
  or (_23571_, _23570_, _06047_);
  or (_23572_, _23571_, _23569_);
  and (_23573_, _15451_, _07648_);
  or (_23574_, _23473_, _06048_);
  or (_23575_, _23574_, _23573_);
  and (_23576_, _23575_, _01336_);
  and (_23577_, _23576_, _23572_);
  or (_23578_, _23577_, _23472_);
  and (_43397_, _23578_, _42882_);
  not (_23579_, \oc8051_golden_model_1.TH1 [0]);
  nor (_23580_, _01336_, _23579_);
  nand (_23581_, _10995_, _07670_);
  nor (_23583_, _07670_, _23579_);
  nor (_23584_, _23583_, _06278_);
  nand (_23585_, _23584_, _23581_);
  and (_23586_, _09120_, _07670_);
  or (_23587_, _23583_, _07012_);
  or (_23588_, _23587_, _23586_);
  and (_23589_, _07670_, _06931_);
  nor (_23590_, _23589_, _23583_);
  nand (_23591_, _23590_, _09815_);
  nor (_23592_, _08127_, _11707_);
  or (_23594_, _23592_, _23583_);
  or (_23595_, _23594_, _06954_);
  and (_23596_, _07670_, \oc8051_golden_model_1.ACC [0]);
  nor (_23597_, _23596_, _23583_);
  nor (_23598_, _23597_, _06939_);
  nor (_23599_, _06938_, _23579_);
  or (_23600_, _23599_, _06102_);
  or (_23601_, _23600_, _23598_);
  and (_23602_, _23601_, _06848_);
  and (_23603_, _23602_, _23595_);
  nor (_23605_, _23590_, _06848_);
  or (_23606_, _23605_, _23603_);
  nand (_23607_, _23606_, _06220_);
  or (_23608_, _23597_, _06220_);
  and (_23609_, _23608_, _09817_);
  nand (_23610_, _23609_, _23607_);
  and (_23611_, _23610_, _23591_);
  and (_23612_, _23611_, _23588_);
  or (_23613_, _23612_, _09833_);
  and (_23614_, _14186_, _07670_);
  or (_23616_, _23614_, _23583_);
  or (_23617_, _23616_, _05669_);
  and (_23618_, _23617_, _06020_);
  and (_23619_, _23618_, _23613_);
  and (_23620_, _07670_, _08672_);
  or (_23621_, _23620_, _23583_);
  and (_23622_, _23621_, _06019_);
  or (_23623_, _23622_, _06112_);
  or (_23624_, _23623_, _23619_);
  and (_23625_, _14086_, _07670_);
  or (_23627_, _23583_, _08751_);
  or (_23628_, _23627_, _23625_);
  and (_23629_, _23628_, _08756_);
  and (_23630_, _23629_, _23624_);
  nor (_23631_, _12302_, _11707_);
  or (_23632_, _23631_, _23583_);
  and (_23633_, _23581_, _06284_);
  and (_23634_, _23633_, _23632_);
  or (_23635_, _23634_, _23630_);
  and (_23636_, _23635_, _07032_);
  nand (_23638_, _23621_, _06108_);
  nor (_23639_, _23638_, _23592_);
  or (_23640_, _23639_, _06277_);
  or (_23641_, _23640_, _23636_);
  and (_23642_, _23641_, _23585_);
  or (_23643_, _23642_, _06130_);
  and (_23644_, _14083_, _07670_);
  or (_23645_, _23583_, _08777_);
  or (_23646_, _23645_, _23644_);
  and (_23647_, _23646_, _08782_);
  and (_23649_, _23647_, _23643_);
  and (_23650_, _23632_, _06292_);
  or (_23651_, _23650_, _19256_);
  or (_23652_, _23651_, _23649_);
  or (_23653_, _23594_, _06408_);
  and (_23654_, _23653_, _01336_);
  and (_23655_, _23654_, _23652_);
  or (_23656_, _23655_, _23580_);
  and (_43399_, _23656_, _42882_);
  not (_23657_, \oc8051_golden_model_1.TH1 [1]);
  nor (_23659_, _01336_, _23657_);
  or (_23660_, _14367_, _11707_);
  or (_23661_, _07670_, \oc8051_golden_model_1.TH1 [1]);
  and (_23662_, _23661_, _09833_);
  and (_23663_, _23662_, _23660_);
  and (_23664_, _09075_, _07670_);
  nor (_23665_, _07670_, _23657_);
  or (_23666_, _23665_, _07012_);
  or (_23667_, _23666_, _23664_);
  and (_23668_, _14284_, _07670_);
  not (_23670_, _23668_);
  and (_23671_, _23670_, _23661_);
  or (_23672_, _23671_, _06954_);
  and (_23673_, _07670_, \oc8051_golden_model_1.ACC [1]);
  or (_23674_, _23673_, _23665_);
  and (_23675_, _23674_, _06938_);
  nor (_23676_, _06938_, _23657_);
  or (_23677_, _23676_, _06102_);
  or (_23678_, _23677_, _23675_);
  and (_23679_, _23678_, _06848_);
  and (_23680_, _23679_, _23672_);
  nor (_23681_, _11707_, _07132_);
  or (_23682_, _23681_, _23665_);
  and (_23683_, _23682_, _06239_);
  or (_23684_, _23683_, _23680_);
  and (_23685_, _23684_, _06220_);
  and (_23686_, _23674_, _06219_);
  or (_23687_, _23686_, _09818_);
  or (_23688_, _23687_, _23685_);
  or (_23689_, _23682_, _09827_);
  and (_23690_, _23689_, _05669_);
  and (_23691_, _23690_, _23688_);
  and (_23692_, _23691_, _23667_);
  or (_23693_, _23692_, _23663_);
  and (_23694_, _23693_, _06020_);
  nand (_23695_, _07670_, _06832_);
  and (_23696_, _23661_, _06019_);
  and (_23697_, _23696_, _23695_);
  or (_23698_, _23697_, _23694_);
  and (_23699_, _23698_, _08751_);
  or (_23701_, _14263_, _11707_);
  and (_23702_, _23661_, _06112_);
  and (_23703_, _23702_, _23701_);
  or (_23704_, _23703_, _06284_);
  or (_23705_, _23704_, _23699_);
  nor (_23706_, _10993_, _11707_);
  or (_23707_, _23706_, _23665_);
  nand (_23708_, _10992_, _07670_);
  and (_23709_, _23708_, _23707_);
  or (_23710_, _23709_, _08756_);
  and (_23712_, _23710_, _07032_);
  and (_23713_, _23712_, _23705_);
  or (_23714_, _14261_, _11707_);
  and (_23715_, _23661_, _06108_);
  and (_23716_, _23715_, _23714_);
  or (_23717_, _23716_, _06277_);
  or (_23718_, _23717_, _23713_);
  nor (_23719_, _23665_, _06278_);
  nand (_23720_, _23719_, _23708_);
  and (_23721_, _23720_, _08777_);
  and (_23723_, _23721_, _23718_);
  or (_23724_, _23695_, _08078_);
  and (_23725_, _23661_, _06130_);
  and (_23726_, _23725_, _23724_);
  or (_23727_, _23726_, _06292_);
  or (_23728_, _23727_, _23723_);
  or (_23729_, _23707_, _08782_);
  and (_23730_, _23729_, _06718_);
  and (_23731_, _23730_, _23728_);
  and (_23732_, _23671_, _06316_);
  or (_23734_, _23732_, _06047_);
  or (_23735_, _23734_, _23731_);
  or (_23736_, _23665_, _06048_);
  or (_23737_, _23736_, _23668_);
  and (_23738_, _23737_, _01336_);
  and (_23739_, _23738_, _23735_);
  or (_23740_, _23739_, _23659_);
  and (_43400_, _23740_, _42882_);
  not (_23741_, \oc8051_golden_model_1.TH1 [2]);
  nor (_23742_, _01336_, _23741_);
  and (_23744_, _09182_, _07670_);
  nor (_23745_, _07670_, _23741_);
  or (_23746_, _23745_, _07012_);
  or (_23747_, _23746_, _23744_);
  nor (_23748_, _11707_, _07530_);
  nor (_23749_, _23748_, _23745_);
  nand (_23750_, _23749_, _09815_);
  and (_23751_, _14493_, _07670_);
  or (_23752_, _23751_, _23745_);
  or (_23753_, _23752_, _06954_);
  and (_23755_, _07670_, \oc8051_golden_model_1.ACC [2]);
  nor (_23756_, _23755_, _23745_);
  nor (_23757_, _23756_, _06939_);
  nor (_23758_, _06938_, _23741_);
  or (_23759_, _23758_, _06102_);
  or (_23760_, _23759_, _23757_);
  and (_23761_, _23760_, _06848_);
  and (_23762_, _23761_, _23753_);
  nor (_23763_, _23749_, _06848_);
  or (_23764_, _23763_, _23762_);
  nand (_23766_, _23764_, _06220_);
  or (_23767_, _23756_, _06220_);
  and (_23768_, _23767_, _09817_);
  nand (_23769_, _23768_, _23766_);
  and (_23770_, _23769_, _23750_);
  and (_23771_, _23770_, _23747_);
  or (_23772_, _23771_, _09833_);
  and (_23773_, _14580_, _07670_);
  or (_23774_, _23745_, _05669_);
  or (_23775_, _23774_, _23773_);
  and (_23777_, _23775_, _06020_);
  and (_23778_, _23777_, _23772_);
  and (_23779_, _07670_, _08730_);
  or (_23780_, _23779_, _23745_);
  and (_23781_, _23780_, _06019_);
  or (_23782_, _23781_, _06112_);
  or (_23783_, _23782_, _23778_);
  and (_23784_, _14596_, _07670_);
  or (_23785_, _23784_, _23745_);
  or (_23786_, _23785_, _08751_);
  and (_23788_, _23786_, _08756_);
  and (_23789_, _23788_, _23783_);
  and (_23790_, _10991_, _07670_);
  or (_23791_, _23790_, _23745_);
  and (_23792_, _23791_, _06284_);
  or (_23793_, _23792_, _23789_);
  and (_23794_, _23793_, _07032_);
  or (_23795_, _23745_, _08177_);
  and (_23796_, _23780_, _06108_);
  and (_23797_, _23796_, _23795_);
  or (_23799_, _23797_, _23794_);
  and (_23800_, _23799_, _06278_);
  nor (_23801_, _23756_, _06278_);
  and (_23802_, _23801_, _23795_);
  or (_23803_, _23802_, _06130_);
  or (_23804_, _23803_, _23800_);
  and (_23805_, _14593_, _07670_);
  or (_23806_, _23745_, _08777_);
  or (_23807_, _23806_, _23805_);
  and (_23808_, _23807_, _08782_);
  and (_23810_, _23808_, _23804_);
  nor (_23811_, _10990_, _11707_);
  or (_23812_, _23811_, _23745_);
  and (_23813_, _23812_, _06292_);
  or (_23814_, _23813_, _23810_);
  and (_23815_, _23814_, _06718_);
  and (_23816_, _23752_, _06316_);
  or (_23817_, _23816_, _06047_);
  or (_23818_, _23817_, _23815_);
  and (_23819_, _14657_, _07670_);
  or (_23821_, _23745_, _06048_);
  or (_23822_, _23821_, _23819_);
  and (_23823_, _23822_, _01336_);
  and (_23824_, _23823_, _23818_);
  or (_23825_, _23824_, _23742_);
  and (_43401_, _23825_, _42882_);
  not (_23826_, \oc8051_golden_model_1.TH1 [3]);
  nor (_23827_, _01336_, _23826_);
  nor (_23828_, _07670_, _23826_);
  or (_23829_, _23828_, _08029_);
  and (_23831_, _07670_, _08662_);
  or (_23832_, _23831_, _23828_);
  and (_23833_, _23832_, _06108_);
  and (_23834_, _23833_, _23829_);
  and (_23835_, _09181_, _07670_);
  or (_23836_, _23828_, _07012_);
  or (_23837_, _23836_, _23835_);
  nor (_23838_, _11707_, _07353_);
  nor (_23839_, _23838_, _23828_);
  nand (_23840_, _23839_, _09815_);
  and (_23842_, _14672_, _07670_);
  or (_23843_, _23842_, _23828_);
  or (_23844_, _23843_, _06954_);
  and (_23845_, _07670_, \oc8051_golden_model_1.ACC [3]);
  nor (_23846_, _23845_, _23828_);
  nor (_23847_, _23846_, _06939_);
  nor (_23848_, _06938_, _23826_);
  or (_23849_, _23848_, _06102_);
  or (_23850_, _23849_, _23847_);
  and (_23851_, _23850_, _06848_);
  and (_23853_, _23851_, _23844_);
  nor (_23854_, _23839_, _06848_);
  or (_23855_, _23854_, _23853_);
  nand (_23856_, _23855_, _06220_);
  or (_23857_, _23846_, _06220_);
  and (_23858_, _23857_, _09817_);
  nand (_23859_, _23858_, _23856_);
  and (_23860_, _23859_, _23840_);
  and (_23861_, _23860_, _23837_);
  or (_23862_, _23861_, _09833_);
  and (_23864_, _14778_, _07670_);
  or (_23865_, _23864_, _23828_);
  or (_23866_, _23865_, _05669_);
  and (_23867_, _23866_, _06020_);
  and (_23868_, _23867_, _23862_);
  and (_23869_, _23832_, _06019_);
  or (_23870_, _23869_, _06112_);
  or (_23871_, _23870_, _23868_);
  and (_23872_, _14793_, _07670_);
  or (_23873_, _23828_, _08751_);
  or (_23875_, _23873_, _23872_);
  and (_23876_, _23875_, _08756_);
  and (_23877_, _23876_, _23871_);
  and (_23878_, _12299_, _07670_);
  or (_23879_, _23878_, _23828_);
  and (_23880_, _23879_, _06284_);
  or (_23881_, _23880_, _23877_);
  and (_23882_, _23881_, _07032_);
  or (_23883_, _23882_, _23834_);
  and (_23884_, _23883_, _06278_);
  nor (_23885_, _23846_, _06278_);
  and (_23886_, _23885_, _23829_);
  or (_23887_, _23886_, _06130_);
  or (_23888_, _23887_, _23884_);
  and (_23889_, _14792_, _07670_);
  or (_23890_, _23828_, _08777_);
  or (_23891_, _23890_, _23889_);
  and (_23892_, _23891_, _08782_);
  and (_23893_, _23892_, _23888_);
  nor (_23894_, _10988_, _11707_);
  or (_23897_, _23894_, _23828_);
  and (_23898_, _23897_, _06292_);
  or (_23899_, _23898_, _23893_);
  and (_23900_, _23899_, _06718_);
  and (_23901_, _23843_, _06316_);
  or (_23902_, _23901_, _06047_);
  or (_23903_, _23902_, _23900_);
  and (_23904_, _14849_, _07670_);
  or (_23905_, _23828_, _06048_);
  or (_23906_, _23905_, _23904_);
  and (_23908_, _23906_, _01336_);
  and (_23909_, _23908_, _23903_);
  or (_23910_, _23909_, _23827_);
  and (_43403_, _23910_, _42882_);
  and (_23911_, _01340_, \oc8051_golden_model_1.TH1 [4]);
  and (_23912_, _11707_, \oc8051_golden_model_1.TH1 [4]);
  or (_23913_, _23912_, _08273_);
  and (_23914_, _08665_, _07670_);
  or (_23915_, _23914_, _23912_);
  and (_23916_, _23915_, _06108_);
  and (_23918_, _23916_, _23913_);
  or (_23919_, _23915_, _06020_);
  and (_23920_, _14887_, _07670_);
  or (_23921_, _23920_, _23912_);
  or (_23922_, _23921_, _06954_);
  and (_23923_, _07670_, \oc8051_golden_model_1.ACC [4]);
  or (_23924_, _23923_, _23912_);
  and (_23925_, _23924_, _06938_);
  and (_23926_, _06939_, \oc8051_golden_model_1.TH1 [4]);
  or (_23927_, _23926_, _06102_);
  or (_23929_, _23927_, _23925_);
  and (_23930_, _23929_, _06848_);
  and (_23931_, _23930_, _23922_);
  nor (_23932_, _08270_, _11707_);
  or (_23933_, _23932_, _23912_);
  and (_23934_, _23933_, _06239_);
  or (_23935_, _23934_, _23931_);
  and (_23936_, _23935_, _06220_);
  and (_23937_, _23924_, _06219_);
  or (_23938_, _23937_, _09818_);
  or (_23940_, _23938_, _23936_);
  and (_23941_, _09180_, _07670_);
  or (_23942_, _23912_, _07012_);
  or (_23943_, _23942_, _23941_);
  or (_23944_, _23933_, _09827_);
  and (_23945_, _23944_, _05669_);
  and (_23946_, _23945_, _23943_);
  and (_23947_, _23946_, _23940_);
  and (_23948_, _14983_, _07670_);
  or (_23949_, _23948_, _23912_);
  and (_23951_, _23949_, _09833_);
  or (_23952_, _23951_, _06019_);
  or (_23953_, _23952_, _23947_);
  and (_23954_, _23953_, _23919_);
  or (_23955_, _23954_, _06112_);
  and (_23956_, _14876_, _07670_);
  or (_23957_, _23912_, _08751_);
  or (_23958_, _23957_, _23956_);
  and (_23959_, _23958_, _08756_);
  and (_23960_, _23959_, _23955_);
  and (_23962_, _10986_, _07670_);
  or (_23963_, _23962_, _23912_);
  and (_23964_, _23963_, _06284_);
  or (_23965_, _23964_, _23960_);
  and (_23966_, _23965_, _07032_);
  or (_23967_, _23966_, _23918_);
  and (_23968_, _23967_, _06278_);
  and (_23969_, _23924_, _06277_);
  and (_23970_, _23969_, _23913_);
  or (_23971_, _23970_, _06130_);
  or (_23973_, _23971_, _23968_);
  and (_23974_, _14873_, _07670_);
  or (_23975_, _23912_, _08777_);
  or (_23976_, _23975_, _23974_);
  and (_23977_, _23976_, _08782_);
  and (_23978_, _23977_, _23973_);
  nor (_23979_, _10985_, _11707_);
  or (_23980_, _23979_, _23912_);
  and (_23981_, _23980_, _06292_);
  or (_23982_, _23981_, _23978_);
  and (_23984_, _23982_, _06718_);
  and (_23985_, _23921_, _06316_);
  or (_23986_, _23985_, _06047_);
  or (_23987_, _23986_, _23984_);
  and (_23988_, _15055_, _07670_);
  or (_23989_, _23912_, _06048_);
  or (_23990_, _23989_, _23988_);
  and (_23991_, _23990_, _01336_);
  and (_23992_, _23991_, _23987_);
  or (_23993_, _23992_, _23911_);
  and (_43404_, _23993_, _42882_);
  and (_23995_, _01340_, \oc8051_golden_model_1.TH1 [5]);
  and (_23996_, _11707_, \oc8051_golden_model_1.TH1 [5]);
  or (_23997_, _23996_, _07980_);
  and (_23998_, _08652_, _07670_);
  or (_23999_, _23998_, _23996_);
  and (_24000_, _23999_, _06108_);
  and (_24001_, _24000_, _23997_);
  or (_24002_, _23999_, _06020_);
  and (_24003_, _15093_, _07670_);
  or (_24005_, _24003_, _23996_);
  or (_24006_, _24005_, _06954_);
  and (_24007_, _07670_, \oc8051_golden_model_1.ACC [5]);
  or (_24008_, _24007_, _23996_);
  and (_24009_, _24008_, _06938_);
  and (_24010_, _06939_, \oc8051_golden_model_1.TH1 [5]);
  or (_24011_, _24010_, _06102_);
  or (_24012_, _24011_, _24009_);
  and (_24013_, _24012_, _06848_);
  and (_24014_, _24013_, _24006_);
  nor (_24016_, _07977_, _11707_);
  or (_24017_, _24016_, _23996_);
  and (_24018_, _24017_, _06239_);
  or (_24019_, _24018_, _24014_);
  and (_24020_, _24019_, _06220_);
  and (_24021_, _24008_, _06219_);
  or (_24022_, _24021_, _09818_);
  or (_24023_, _24022_, _24020_);
  and (_24024_, _09179_, _07670_);
  or (_24025_, _23996_, _07012_);
  or (_24027_, _24025_, _24024_);
  or (_24028_, _24017_, _09827_);
  and (_24029_, _24028_, _05669_);
  and (_24030_, _24029_, _24027_);
  and (_24031_, _24030_, _24023_);
  and (_24032_, _15179_, _07670_);
  or (_24033_, _24032_, _23996_);
  and (_24034_, _24033_, _09833_);
  or (_24035_, _24034_, _06019_);
  or (_24036_, _24035_, _24031_);
  and (_24038_, _24036_, _24002_);
  or (_24039_, _24038_, _06112_);
  and (_24040_, _15195_, _07670_);
  or (_24041_, _23996_, _08751_);
  or (_24042_, _24041_, _24040_);
  and (_24043_, _24042_, _08756_);
  and (_24044_, _24043_, _24039_);
  and (_24045_, _12306_, _07670_);
  or (_24046_, _24045_, _23996_);
  and (_24047_, _24046_, _06284_);
  or (_24049_, _24047_, _24044_);
  and (_24050_, _24049_, _07032_);
  or (_24051_, _24050_, _24001_);
  and (_24052_, _24051_, _06278_);
  and (_24053_, _24008_, _06277_);
  and (_24054_, _24053_, _23997_);
  or (_24055_, _24054_, _06130_);
  or (_24056_, _24055_, _24052_);
  and (_24057_, _15194_, _07670_);
  or (_24058_, _23996_, _08777_);
  or (_24060_, _24058_, _24057_);
  and (_24061_, _24060_, _08782_);
  and (_24062_, _24061_, _24056_);
  nor (_24063_, _10982_, _11707_);
  or (_24064_, _24063_, _23996_);
  and (_24065_, _24064_, _06292_);
  or (_24066_, _24065_, _24062_);
  and (_24067_, _24066_, _06718_);
  and (_24068_, _24005_, _06316_);
  or (_24069_, _24068_, _06047_);
  or (_24070_, _24069_, _24067_);
  and (_24071_, _15253_, _07670_);
  or (_24072_, _23996_, _06048_);
  or (_24073_, _24072_, _24071_);
  and (_24074_, _24073_, _01336_);
  and (_24075_, _24074_, _24070_);
  or (_24076_, _24075_, _23995_);
  and (_43405_, _24076_, _42882_);
  and (_24077_, _01340_, \oc8051_golden_model_1.TH1 [6]);
  and (_24078_, _11707_, \oc8051_golden_model_1.TH1 [6]);
  or (_24081_, _24078_, _07886_);
  and (_24082_, _15389_, _07670_);
  or (_24083_, _24082_, _24078_);
  and (_24084_, _24083_, _06108_);
  and (_24085_, _24084_, _24081_);
  or (_24086_, _24083_, _06020_);
  and (_24087_, _15293_, _07670_);
  or (_24088_, _24087_, _24078_);
  or (_24089_, _24088_, _06954_);
  and (_24090_, _07670_, \oc8051_golden_model_1.ACC [6]);
  or (_24092_, _24090_, _24078_);
  and (_24093_, _24092_, _06938_);
  and (_24094_, _06939_, \oc8051_golden_model_1.TH1 [6]);
  or (_24095_, _24094_, _06102_);
  or (_24096_, _24095_, _24093_);
  and (_24097_, _24096_, _06848_);
  and (_24098_, _24097_, _24089_);
  nor (_24099_, _07883_, _11707_);
  or (_24100_, _24099_, _24078_);
  and (_24101_, _24100_, _06239_);
  or (_24103_, _24101_, _24098_);
  and (_24104_, _24103_, _06220_);
  and (_24105_, _24092_, _06219_);
  or (_24106_, _24105_, _09818_);
  or (_24107_, _24106_, _24104_);
  and (_24108_, _09178_, _07670_);
  or (_24109_, _24078_, _07012_);
  or (_24110_, _24109_, _24108_);
  or (_24111_, _24100_, _09827_);
  and (_24112_, _24111_, _05669_);
  and (_24114_, _24112_, _24110_);
  and (_24115_, _24114_, _24107_);
  and (_24116_, _15382_, _07670_);
  or (_24117_, _24116_, _24078_);
  and (_24118_, _24117_, _09833_);
  or (_24119_, _24118_, _06019_);
  or (_24120_, _24119_, _24115_);
  and (_24121_, _24120_, _24086_);
  or (_24122_, _24121_, _06112_);
  and (_24123_, _15399_, _07670_);
  or (_24125_, _24123_, _24078_);
  or (_24126_, _24125_, _08751_);
  and (_24127_, _24126_, _08756_);
  and (_24128_, _24127_, _24122_);
  and (_24129_, _10980_, _07670_);
  or (_24130_, _24129_, _24078_);
  and (_24131_, _24130_, _06284_);
  or (_24132_, _24131_, _24128_);
  and (_24133_, _24132_, _07032_);
  or (_24134_, _24133_, _24085_);
  and (_24136_, _24134_, _06278_);
  and (_24137_, _24092_, _06277_);
  and (_24138_, _24137_, _24081_);
  or (_24139_, _24138_, _06130_);
  or (_24140_, _24139_, _24136_);
  and (_24141_, _15396_, _07670_);
  or (_24142_, _24078_, _08777_);
  or (_24143_, _24142_, _24141_);
  and (_24144_, _24143_, _08782_);
  and (_24145_, _24144_, _24140_);
  nor (_24147_, _10979_, _11707_);
  or (_24148_, _24147_, _24078_);
  and (_24149_, _24148_, _06292_);
  or (_24150_, _24149_, _24145_);
  and (_24151_, _24150_, _06718_);
  and (_24152_, _24088_, _06316_);
  or (_24153_, _24152_, _06047_);
  or (_24154_, _24153_, _24151_);
  and (_24155_, _15451_, _07670_);
  or (_24156_, _24078_, _06048_);
  or (_24158_, _24156_, _24155_);
  and (_24159_, _24158_, _01336_);
  and (_24160_, _24159_, _24154_);
  or (_24161_, _24160_, _24077_);
  and (_43406_, _24161_, _42882_);
  not (_24162_, \oc8051_golden_model_1.TH0 [0]);
  nor (_24163_, _01336_, _24162_);
  nand (_24164_, _10995_, _07663_);
  nor (_24165_, _07663_, _24162_);
  nor (_24166_, _24165_, _06278_);
  nand (_24168_, _24166_, _24164_);
  and (_24169_, _09120_, _07663_);
  or (_24170_, _24165_, _07012_);
  or (_24171_, _24170_, _24169_);
  and (_24172_, _07663_, _06931_);
  nor (_24173_, _24172_, _24165_);
  nand (_24174_, _24173_, _09815_);
  nor (_24175_, _08127_, _11784_);
  or (_24176_, _24175_, _24165_);
  and (_24177_, _24176_, _06102_);
  nor (_24179_, _06938_, _24162_);
  and (_24180_, _07663_, \oc8051_golden_model_1.ACC [0]);
  nor (_24181_, _24180_, _24165_);
  nor (_24182_, _24181_, _06939_);
  or (_24183_, _24182_, _24179_);
  and (_24184_, _24183_, _06954_);
  or (_24185_, _24184_, _06239_);
  or (_24186_, _24185_, _24177_);
  nand (_24187_, _24173_, _06239_);
  and (_24188_, _24187_, _06220_);
  nand (_24190_, _24188_, _24186_);
  or (_24191_, _24181_, _06220_);
  and (_24192_, _24191_, _09817_);
  nand (_24193_, _24192_, _24190_);
  and (_24194_, _24193_, _24174_);
  and (_24195_, _24194_, _24171_);
  or (_24196_, _24195_, _09833_);
  and (_24197_, _14186_, _07663_);
  or (_24198_, _24165_, _05669_);
  or (_24199_, _24198_, _24197_);
  and (_24201_, _24199_, _06020_);
  and (_24202_, _24201_, _24196_);
  and (_24203_, _07663_, _08672_);
  or (_24204_, _24203_, _24165_);
  and (_24205_, _24204_, _06019_);
  or (_24206_, _24205_, _06112_);
  or (_24207_, _24206_, _24202_);
  and (_24208_, _14086_, _07663_);
  or (_24209_, _24165_, _08751_);
  or (_24210_, _24209_, _24208_);
  and (_24212_, _24210_, _08756_);
  and (_24213_, _24212_, _24207_);
  nor (_24214_, _12302_, _11784_);
  or (_24215_, _24214_, _24165_);
  and (_24216_, _24164_, _06284_);
  and (_24217_, _24216_, _24215_);
  or (_24218_, _24217_, _24213_);
  and (_24219_, _24218_, _07032_);
  nand (_24220_, _24204_, _06108_);
  nor (_24221_, _24220_, _24175_);
  or (_24223_, _24221_, _06277_);
  or (_24224_, _24223_, _24219_);
  and (_24225_, _24224_, _24168_);
  or (_24226_, _24225_, _06130_);
  and (_24227_, _14083_, _07663_);
  or (_24228_, _24165_, _08777_);
  or (_24229_, _24228_, _24227_);
  and (_24230_, _24229_, _08782_);
  and (_24231_, _24230_, _24226_);
  and (_24232_, _24215_, _06292_);
  or (_24234_, _24232_, _19256_);
  or (_24235_, _24234_, _24231_);
  or (_24236_, _24176_, _06408_);
  and (_24237_, _24236_, _01336_);
  and (_24238_, _24237_, _24235_);
  or (_24239_, _24238_, _24163_);
  and (_43408_, _24239_, _42882_);
  not (_24240_, \oc8051_golden_model_1.TH0 [1]);
  nor (_24241_, _01336_, _24240_);
  or (_24242_, _14367_, _11784_);
  or (_24244_, _07663_, \oc8051_golden_model_1.TH0 [1]);
  and (_24245_, _24244_, _09833_);
  and (_24246_, _24245_, _24242_);
  and (_24247_, _09075_, _07663_);
  nor (_24248_, _07663_, _24240_);
  or (_24249_, _24248_, _07012_);
  or (_24250_, _24249_, _24247_);
  and (_24251_, _14284_, _07663_);
  not (_24252_, _24251_);
  and (_24253_, _24252_, _24244_);
  or (_24255_, _24253_, _06954_);
  and (_24256_, _07663_, \oc8051_golden_model_1.ACC [1]);
  or (_24257_, _24256_, _24248_);
  and (_24258_, _24257_, _06938_);
  nor (_24259_, _06938_, _24240_);
  or (_24260_, _24259_, _06102_);
  or (_24261_, _24260_, _24258_);
  and (_24262_, _24261_, _06848_);
  and (_24263_, _24262_, _24255_);
  nor (_24264_, _11784_, _07132_);
  or (_24266_, _24264_, _24248_);
  and (_24267_, _24266_, _06239_);
  or (_24268_, _24267_, _24263_);
  and (_24269_, _24268_, _06220_);
  and (_24270_, _24257_, _06219_);
  or (_24271_, _24270_, _09818_);
  or (_24272_, _24271_, _24269_);
  or (_24273_, _24266_, _09827_);
  and (_24274_, _24273_, _05669_);
  and (_24275_, _24274_, _24272_);
  and (_24277_, _24275_, _24250_);
  or (_24278_, _24277_, _24246_);
  and (_24279_, _24278_, _06020_);
  nand (_24280_, _07663_, _06832_);
  and (_24281_, _24244_, _06019_);
  and (_24282_, _24281_, _24280_);
  or (_24283_, _24282_, _24279_);
  and (_24284_, _24283_, _08751_);
  or (_24285_, _14263_, _11784_);
  and (_24286_, _24244_, _06112_);
  and (_24288_, _24286_, _24285_);
  or (_24289_, _24288_, _06284_);
  or (_24290_, _24289_, _24284_);
  nor (_24291_, _10993_, _11784_);
  or (_24292_, _24291_, _24248_);
  nand (_24293_, _10992_, _07663_);
  and (_24294_, _24293_, _24292_);
  or (_24295_, _24294_, _08756_);
  and (_24296_, _24295_, _07032_);
  and (_24297_, _24296_, _24290_);
  or (_24299_, _14261_, _11784_);
  and (_24300_, _24244_, _06108_);
  and (_24301_, _24300_, _24299_);
  or (_24302_, _24301_, _06277_);
  or (_24303_, _24302_, _24297_);
  nor (_24304_, _24248_, _06278_);
  nand (_24305_, _24304_, _24293_);
  and (_24306_, _24305_, _08777_);
  and (_24307_, _24306_, _24303_);
  or (_24308_, _24280_, _08078_);
  and (_24310_, _24244_, _06130_);
  and (_24311_, _24310_, _24308_);
  or (_24312_, _24311_, _06292_);
  or (_24313_, _24312_, _24307_);
  or (_24314_, _24292_, _08782_);
  and (_24315_, _24314_, _06718_);
  and (_24316_, _24315_, _24313_);
  and (_24317_, _24253_, _06316_);
  or (_24318_, _24317_, _06047_);
  or (_24319_, _24318_, _24316_);
  or (_24321_, _24248_, _06048_);
  or (_24322_, _24321_, _24251_);
  and (_24323_, _24322_, _01336_);
  and (_24324_, _24323_, _24319_);
  or (_24325_, _24324_, _24241_);
  and (_43409_, _24325_, _42882_);
  not (_24326_, \oc8051_golden_model_1.TH0 [2]);
  nor (_24327_, _01336_, _24326_);
  and (_24328_, _09182_, _07663_);
  nor (_24329_, _07663_, _24326_);
  or (_24331_, _24329_, _07012_);
  or (_24332_, _24331_, _24328_);
  nor (_24333_, _11784_, _07530_);
  nor (_24334_, _24333_, _24329_);
  nand (_24335_, _24334_, _09815_);
  and (_24336_, _14493_, _07663_);
  or (_24337_, _24336_, _24329_);
  or (_24338_, _24337_, _06954_);
  and (_24339_, _07663_, \oc8051_golden_model_1.ACC [2]);
  nor (_24340_, _24339_, _24329_);
  nor (_24342_, _24340_, _06939_);
  nor (_24343_, _06938_, _24326_);
  or (_24344_, _24343_, _06102_);
  or (_24345_, _24344_, _24342_);
  and (_24346_, _24345_, _06848_);
  and (_24347_, _24346_, _24338_);
  nor (_24348_, _24334_, _06848_);
  or (_24349_, _24348_, _24347_);
  nand (_24350_, _24349_, _06220_);
  or (_24351_, _24340_, _06220_);
  and (_24353_, _24351_, _09817_);
  nand (_24354_, _24353_, _24350_);
  and (_24355_, _24354_, _24335_);
  and (_24356_, _24355_, _24332_);
  or (_24357_, _24356_, _09833_);
  and (_24358_, _14580_, _07663_);
  or (_24359_, _24358_, _24329_);
  or (_24360_, _24359_, _05669_);
  and (_24361_, _24360_, _06020_);
  and (_24362_, _24361_, _24357_);
  and (_24364_, _07663_, _08730_);
  or (_24365_, _24364_, _24329_);
  and (_24366_, _24365_, _06019_);
  or (_24367_, _24366_, _06112_);
  or (_24368_, _24367_, _24362_);
  and (_24369_, _14596_, _07663_);
  or (_24370_, _24369_, _24329_);
  or (_24371_, _24370_, _08751_);
  and (_24372_, _24371_, _08756_);
  and (_24373_, _24372_, _24368_);
  and (_24376_, _10991_, _07663_);
  or (_24377_, _24376_, _24329_);
  and (_24378_, _24377_, _06284_);
  or (_24379_, _24378_, _24373_);
  and (_24380_, _24379_, _07032_);
  or (_24381_, _24329_, _08177_);
  and (_24382_, _24365_, _06108_);
  and (_24383_, _24382_, _24381_);
  or (_24384_, _24383_, _24380_);
  and (_24385_, _24384_, _06278_);
  nor (_24387_, _24340_, _06278_);
  and (_24388_, _24387_, _24381_);
  or (_24389_, _24388_, _06130_);
  or (_24390_, _24389_, _24385_);
  and (_24391_, _14593_, _07663_);
  or (_24392_, _24329_, _08777_);
  or (_24393_, _24392_, _24391_);
  and (_24394_, _24393_, _08782_);
  and (_24395_, _24394_, _24390_);
  nor (_24396_, _10990_, _11784_);
  or (_24398_, _24396_, _24329_);
  and (_24399_, _24398_, _06292_);
  or (_24400_, _24399_, _24395_);
  and (_24401_, _24400_, _06718_);
  and (_24402_, _24337_, _06316_);
  or (_24403_, _24402_, _06047_);
  or (_24404_, _24403_, _24401_);
  and (_24405_, _14657_, _07663_);
  or (_24406_, _24329_, _06048_);
  or (_24407_, _24406_, _24405_);
  and (_24409_, _24407_, _01336_);
  and (_24410_, _24409_, _24404_);
  or (_24411_, _24410_, _24327_);
  and (_43410_, _24411_, _42882_);
  not (_24412_, \oc8051_golden_model_1.TH0 [3]);
  nor (_24413_, _01336_, _24412_);
  nor (_24414_, _07663_, _24412_);
  or (_24415_, _24414_, _08029_);
  and (_24416_, _07663_, _08662_);
  or (_24417_, _24416_, _24414_);
  and (_24419_, _24417_, _06108_);
  and (_24420_, _24419_, _24415_);
  and (_24421_, _09181_, _07663_);
  or (_24422_, _24414_, _07012_);
  or (_24423_, _24422_, _24421_);
  nor (_24424_, _11784_, _07353_);
  nor (_24425_, _24424_, _24414_);
  nand (_24426_, _24425_, _09815_);
  and (_24427_, _14672_, _07663_);
  or (_24428_, _24427_, _24414_);
  or (_24430_, _24428_, _06954_);
  and (_24431_, _07663_, \oc8051_golden_model_1.ACC [3]);
  nor (_24432_, _24431_, _24414_);
  nor (_24433_, _24432_, _06939_);
  nor (_24434_, _06938_, _24412_);
  or (_24435_, _24434_, _06102_);
  or (_24436_, _24435_, _24433_);
  and (_24437_, _24436_, _06848_);
  and (_24438_, _24437_, _24430_);
  nor (_24439_, _24425_, _06848_);
  or (_24441_, _24439_, _24438_);
  nand (_24442_, _24441_, _06220_);
  or (_24443_, _24432_, _06220_);
  and (_24444_, _24443_, _09817_);
  nand (_24445_, _24444_, _24442_);
  and (_24446_, _24445_, _24426_);
  and (_24447_, _24446_, _24423_);
  or (_24448_, _24447_, _09833_);
  and (_24449_, _14778_, _07663_);
  or (_24450_, _24414_, _05669_);
  or (_24452_, _24450_, _24449_);
  and (_24453_, _24452_, _06020_);
  and (_24454_, _24453_, _24448_);
  and (_24455_, _24417_, _06019_);
  or (_24456_, _24455_, _06112_);
  or (_24457_, _24456_, _24454_);
  and (_24458_, _14793_, _07663_);
  or (_24459_, _24414_, _08751_);
  or (_24460_, _24459_, _24458_);
  and (_24461_, _24460_, _08756_);
  and (_24463_, _24461_, _24457_);
  and (_24464_, _12299_, _07663_);
  or (_24465_, _24464_, _24414_);
  and (_24466_, _24465_, _06284_);
  or (_24467_, _24466_, _24463_);
  and (_24468_, _24467_, _07032_);
  or (_24469_, _24468_, _24420_);
  and (_24470_, _24469_, _06278_);
  nor (_24471_, _24432_, _06278_);
  and (_24472_, _24471_, _24415_);
  or (_24474_, _24472_, _06130_);
  or (_24475_, _24474_, _24470_);
  and (_24476_, _14792_, _07663_);
  or (_24477_, _24414_, _08777_);
  or (_24478_, _24477_, _24476_);
  and (_24479_, _24478_, _08782_);
  and (_24480_, _24479_, _24475_);
  nor (_24481_, _10988_, _11784_);
  or (_24482_, _24481_, _24414_);
  and (_24483_, _24482_, _06292_);
  or (_24485_, _24483_, _24480_);
  and (_24486_, _24485_, _06718_);
  and (_24487_, _24428_, _06316_);
  or (_24488_, _24487_, _06047_);
  or (_24489_, _24488_, _24486_);
  and (_24490_, _14849_, _07663_);
  or (_24491_, _24414_, _06048_);
  or (_24492_, _24491_, _24490_);
  and (_24493_, _24492_, _01336_);
  and (_24494_, _24493_, _24489_);
  or (_24496_, _24494_, _24413_);
  and (_43411_, _24496_, _42882_);
  and (_24497_, _01340_, \oc8051_golden_model_1.TH0 [4]);
  and (_24498_, _11784_, \oc8051_golden_model_1.TH0 [4]);
  or (_24499_, _24498_, _08273_);
  and (_24500_, _08665_, _07663_);
  or (_24501_, _24500_, _24498_);
  and (_24502_, _24501_, _06108_);
  and (_24503_, _24502_, _24499_);
  or (_24504_, _24501_, _06020_);
  and (_24506_, _14887_, _07663_);
  or (_24507_, _24506_, _24498_);
  or (_24508_, _24507_, _06954_);
  and (_24509_, _07663_, \oc8051_golden_model_1.ACC [4]);
  or (_24510_, _24509_, _24498_);
  and (_24511_, _24510_, _06938_);
  and (_24512_, _06939_, \oc8051_golden_model_1.TH0 [4]);
  or (_24513_, _24512_, _06102_);
  or (_24514_, _24513_, _24511_);
  and (_24515_, _24514_, _06848_);
  and (_24517_, _24515_, _24508_);
  nor (_24518_, _08270_, _11784_);
  or (_24519_, _24518_, _24498_);
  and (_24520_, _24519_, _06239_);
  or (_24521_, _24520_, _24517_);
  and (_24522_, _24521_, _06220_);
  and (_24523_, _24510_, _06219_);
  or (_24524_, _24523_, _09818_);
  or (_24525_, _24524_, _24522_);
  and (_24526_, _09180_, _07663_);
  or (_24528_, _24498_, _07012_);
  or (_24529_, _24528_, _24526_);
  or (_24530_, _24519_, _09827_);
  and (_24531_, _24530_, _05669_);
  and (_24532_, _24531_, _24529_);
  and (_24533_, _24532_, _24525_);
  and (_24534_, _14983_, _07663_);
  or (_24535_, _24534_, _24498_);
  and (_24536_, _24535_, _09833_);
  or (_24537_, _24536_, _06019_);
  or (_24539_, _24537_, _24533_);
  and (_24540_, _24539_, _24504_);
  or (_24541_, _24540_, _06112_);
  and (_24542_, _14876_, _07663_);
  or (_24543_, _24542_, _24498_);
  or (_24544_, _24543_, _08751_);
  and (_24545_, _24544_, _08756_);
  and (_24546_, _24545_, _24541_);
  and (_24547_, _10986_, _07663_);
  or (_24548_, _24547_, _24498_);
  and (_24550_, _24548_, _06284_);
  or (_24551_, _24550_, _24546_);
  and (_24552_, _24551_, _07032_);
  or (_24553_, _24552_, _24503_);
  and (_24554_, _24553_, _06278_);
  and (_24555_, _24510_, _06277_);
  and (_24556_, _24555_, _24499_);
  or (_24557_, _24556_, _06130_);
  or (_24558_, _24557_, _24554_);
  and (_24559_, _14873_, _07663_);
  or (_24561_, _24498_, _08777_);
  or (_24562_, _24561_, _24559_);
  and (_24563_, _24562_, _08782_);
  and (_24564_, _24563_, _24558_);
  nor (_24565_, _10985_, _11784_);
  or (_24566_, _24565_, _24498_);
  and (_24567_, _24566_, _06292_);
  or (_24568_, _24567_, _24564_);
  and (_24569_, _24568_, _06718_);
  and (_24570_, _24507_, _06316_);
  or (_24572_, _24570_, _06047_);
  or (_24573_, _24572_, _24569_);
  and (_24574_, _15055_, _07663_);
  or (_24575_, _24498_, _06048_);
  or (_24576_, _24575_, _24574_);
  and (_24577_, _24576_, _01336_);
  and (_24578_, _24577_, _24573_);
  or (_24579_, _24578_, _24497_);
  and (_43412_, _24579_, _42882_);
  and (_24580_, _01340_, \oc8051_golden_model_1.TH0 [5]);
  and (_24582_, _11784_, \oc8051_golden_model_1.TH0 [5]);
  or (_24583_, _24582_, _07980_);
  and (_24584_, _08652_, _07663_);
  or (_24585_, _24584_, _24582_);
  and (_24586_, _24585_, _06108_);
  and (_24587_, _24586_, _24583_);
  or (_24588_, _24585_, _06020_);
  and (_24589_, _15093_, _07663_);
  or (_24590_, _24589_, _24582_);
  or (_24591_, _24590_, _06954_);
  and (_24593_, _07663_, \oc8051_golden_model_1.ACC [5]);
  or (_24594_, _24593_, _24582_);
  and (_24595_, _24594_, _06938_);
  and (_24596_, _06939_, \oc8051_golden_model_1.TH0 [5]);
  or (_24597_, _24596_, _06102_);
  or (_24598_, _24597_, _24595_);
  and (_24599_, _24598_, _06848_);
  and (_24600_, _24599_, _24591_);
  nor (_24601_, _07977_, _11784_);
  or (_24602_, _24601_, _24582_);
  and (_24603_, _24602_, _06239_);
  or (_24604_, _24603_, _24600_);
  and (_24605_, _24604_, _06220_);
  and (_24606_, _24594_, _06219_);
  or (_24607_, _24606_, _09818_);
  or (_24608_, _24607_, _24605_);
  and (_24609_, _09179_, _07663_);
  or (_24610_, _24582_, _07012_);
  or (_24611_, _24610_, _24609_);
  or (_24612_, _24602_, _09827_);
  and (_24615_, _24612_, _05669_);
  and (_24616_, _24615_, _24611_);
  and (_24617_, _24616_, _24608_);
  and (_24618_, _15179_, _07663_);
  or (_24619_, _24618_, _24582_);
  and (_24620_, _24619_, _09833_);
  or (_24621_, _24620_, _06019_);
  or (_24622_, _24621_, _24617_);
  and (_24623_, _24622_, _24588_);
  or (_24624_, _24623_, _06112_);
  and (_24626_, _15195_, _07663_);
  or (_24627_, _24582_, _08751_);
  or (_24628_, _24627_, _24626_);
  and (_24629_, _24628_, _08756_);
  and (_24630_, _24629_, _24624_);
  and (_24631_, _12306_, _07663_);
  or (_24632_, _24631_, _24582_);
  and (_24633_, _24632_, _06284_);
  or (_24634_, _24633_, _24630_);
  and (_24635_, _24634_, _07032_);
  or (_24637_, _24635_, _24587_);
  and (_24638_, _24637_, _06278_);
  and (_24639_, _24594_, _06277_);
  and (_24640_, _24639_, _24583_);
  or (_24641_, _24640_, _06130_);
  or (_24642_, _24641_, _24638_);
  and (_24643_, _15194_, _07663_);
  or (_24644_, _24582_, _08777_);
  or (_24645_, _24644_, _24643_);
  and (_24646_, _24645_, _08782_);
  and (_24648_, _24646_, _24642_);
  nor (_24649_, _10982_, _11784_);
  or (_24650_, _24649_, _24582_);
  and (_24651_, _24650_, _06292_);
  or (_24652_, _24651_, _24648_);
  and (_24653_, _24652_, _06718_);
  and (_24654_, _24590_, _06316_);
  or (_24655_, _24654_, _06047_);
  or (_24656_, _24655_, _24653_);
  and (_24657_, _15253_, _07663_);
  or (_24659_, _24582_, _06048_);
  or (_24660_, _24659_, _24657_);
  and (_24661_, _24660_, _01336_);
  and (_24662_, _24661_, _24656_);
  or (_24663_, _24662_, _24580_);
  and (_43413_, _24663_, _42882_);
  and (_24664_, _01340_, \oc8051_golden_model_1.TH0 [6]);
  and (_24665_, _11784_, \oc8051_golden_model_1.TH0 [6]);
  or (_24666_, _24665_, _07886_);
  and (_24667_, _15389_, _07663_);
  or (_24669_, _24667_, _24665_);
  and (_24670_, _24669_, _06108_);
  and (_24671_, _24670_, _24666_);
  or (_24672_, _24669_, _06020_);
  and (_24673_, _15293_, _07663_);
  or (_24674_, _24673_, _24665_);
  or (_24675_, _24674_, _06954_);
  and (_24676_, _07663_, \oc8051_golden_model_1.ACC [6]);
  or (_24677_, _24676_, _24665_);
  and (_24678_, _24677_, _06938_);
  and (_24680_, _06939_, \oc8051_golden_model_1.TH0 [6]);
  or (_24681_, _24680_, _06102_);
  or (_24682_, _24681_, _24678_);
  and (_24683_, _24682_, _06848_);
  and (_24684_, _24683_, _24675_);
  nor (_24685_, _07883_, _11784_);
  or (_24686_, _24685_, _24665_);
  and (_24687_, _24686_, _06239_);
  or (_24688_, _24687_, _24684_);
  and (_24689_, _24688_, _06220_);
  and (_24691_, _24677_, _06219_);
  or (_24692_, _24691_, _09818_);
  or (_24693_, _24692_, _24689_);
  and (_24694_, _09178_, _07663_);
  or (_24695_, _24665_, _07012_);
  or (_24696_, _24695_, _24694_);
  or (_24697_, _24686_, _09827_);
  and (_24698_, _24697_, _05669_);
  and (_24699_, _24698_, _24696_);
  and (_24700_, _24699_, _24693_);
  and (_24702_, _15382_, _07663_);
  or (_24703_, _24702_, _24665_);
  and (_24704_, _24703_, _09833_);
  or (_24705_, _24704_, _06019_);
  or (_24706_, _24705_, _24700_);
  and (_24707_, _24706_, _24672_);
  or (_24708_, _24707_, _06112_);
  and (_24709_, _15399_, _07663_);
  or (_24710_, _24665_, _08751_);
  or (_24711_, _24710_, _24709_);
  and (_24713_, _24711_, _08756_);
  and (_24714_, _24713_, _24708_);
  and (_24715_, _10980_, _07663_);
  or (_24716_, _24715_, _24665_);
  and (_24717_, _24716_, _06284_);
  or (_24718_, _24717_, _24714_);
  and (_24719_, _24718_, _07032_);
  or (_24720_, _24719_, _24671_);
  and (_24721_, _24720_, _06278_);
  and (_24722_, _24677_, _06277_);
  and (_24724_, _24722_, _24666_);
  or (_24725_, _24724_, _06130_);
  or (_24726_, _24725_, _24721_);
  and (_24727_, _15396_, _07663_);
  or (_24728_, _24665_, _08777_);
  or (_24729_, _24728_, _24727_);
  and (_24730_, _24729_, _08782_);
  and (_24731_, _24730_, _24726_);
  nor (_24732_, _10979_, _11784_);
  or (_24733_, _24732_, _24665_);
  and (_24735_, _24733_, _06292_);
  or (_24736_, _24735_, _24731_);
  and (_24737_, _24736_, _06718_);
  and (_24738_, _24674_, _06316_);
  or (_24739_, _24738_, _06047_);
  or (_24740_, _24739_, _24737_);
  and (_24741_, _15451_, _07663_);
  or (_24742_, _24665_, _06048_);
  or (_24743_, _24742_, _24741_);
  and (_24744_, _24743_, _01336_);
  and (_24746_, _24744_, _24740_);
  or (_24747_, _24746_, _24664_);
  and (_43414_, _24747_, _42882_);
  nor (_24748_, _06119_, _05751_);
  not (_24749_, _24748_);
  and (_24750_, _24749_, _06633_);
  and (_24751_, _12779_, _12771_);
  nor (_24752_, _24751_, _05346_);
  and (_24753_, _12749_, _12756_);
  nor (_24754_, _24753_, _05346_);
  and (_24756_, _11872_, _11016_);
  nor (_24757_, _24756_, _05346_);
  and (_24758_, _12523_, _10855_);
  not (_24759_, _05740_);
  nor (_24760_, _06633_, _24759_);
  nor (_24761_, _10612_, _05346_);
  and (_24762_, _10612_, _05346_);
  nor (_24763_, _24762_, _24761_);
  nor (_24764_, _24763_, _12498_);
  not (_24765_, _05736_);
  and (_24767_, _12002_, _07032_);
  nor (_24768_, _24767_, _05346_);
  not (_24769_, _05727_);
  nor (_24770_, _12006_, _06112_);
  nor (_24771_, _24770_, _05346_);
  and (_24772_, _06019_, _05346_);
  nor (_24773_, _06110_, _09833_);
  and (_24774_, _24773_, _12389_);
  nor (_24775_, _24774_, _05346_);
  nor (_24776_, _06633_, _05694_);
  and (_24778_, _12239_, _12231_);
  nor (_24779_, _24778_, _05346_);
  and (_24780_, _06633_, _06943_);
  nor (_24781_, _12205_, _05346_);
  nor (_24782_, _12214_, _05346_);
  and (_24783_, _12214_, _05346_);
  nor (_24784_, _24783_, _24782_);
  and (_24785_, _12205_, _07233_);
  not (_24786_, _24785_);
  nor (_24787_, _24786_, _24784_);
  nor (_24789_, _24787_, _24781_);
  not (_24790_, _24789_);
  nor (_24791_, _24790_, _24780_);
  nor (_24792_, _24791_, _08384_);
  and (_24793_, _12197_, \oc8051_golden_model_1.PC [0]);
  and (_24794_, _06016_, _05346_);
  nor (_24795_, _24794_, _11928_);
  and (_24796_, _24795_, _12199_);
  or (_24797_, _24796_, _24793_);
  nor (_24798_, _24797_, _08383_);
  nor (_24800_, _24798_, _24792_);
  nor (_24801_, _24800_, _06948_);
  and (_24802_, _06948_, \oc8051_golden_model_1.PC [0]);
  nor (_24803_, _24802_, _24801_);
  and (_24804_, _24803_, _06954_);
  not (_24805_, _12182_);
  and (_24806_, _06633_, \oc8051_golden_model_1.PC [0]);
  nor (_24807_, _24806_, _12088_);
  not (_24808_, _24807_);
  and (_24809_, _24808_, _12187_);
  and (_24811_, _12189_, \oc8051_golden_model_1.PC [0]);
  or (_24812_, _24811_, _06954_);
  nor (_24813_, _24812_, _24809_);
  nor (_24814_, _24813_, _24805_);
  not (_24815_, _24814_);
  nor (_24816_, _24815_, _24804_);
  nor (_24817_, _12182_, _05346_);
  nor (_24818_, _24817_, _07272_);
  not (_24819_, _24818_);
  nor (_24820_, _24819_, _24816_);
  nor (_24822_, _06633_, _05690_);
  not (_24823_, _24778_);
  nor (_24824_, _24823_, _24822_);
  not (_24825_, _24824_);
  nor (_24826_, _24825_, _24820_);
  or (_24827_, _24826_, _12243_);
  nor (_24828_, _24827_, _24779_);
  nor (_24829_, _24828_, _24776_);
  or (_24830_, _24829_, _12256_);
  and (_24831_, _12289_, \oc8051_golden_model_1.PC [0]);
  nor (_24833_, _24807_, _12289_);
  or (_24834_, _24833_, _12255_);
  or (_24835_, _24834_, _24831_);
  and (_24836_, _24835_, _12258_);
  and (_24837_, _24836_, _24830_);
  nor (_24838_, _24837_, _06121_);
  and (_24839_, _12172_, _05346_);
  and (_24840_, _24807_, _12174_);
  or (_24841_, _24840_, _12258_);
  or (_24842_, _24841_, _24839_);
  and (_24844_, _24842_, _24838_);
  and (_24845_, _12310_, _05346_);
  nor (_24846_, _24808_, _12310_);
  nor (_24847_, _24846_, _24845_);
  nor (_24848_, _24847_, _06509_);
  nor (_24849_, _24848_, _24844_);
  nor (_24850_, _24849_, _06115_);
  and (_24851_, _12329_, _05346_);
  nor (_24852_, _24808_, _12329_);
  or (_24853_, _24852_, _24851_);
  and (_24855_, _24853_, _06115_);
  or (_24856_, _24855_, _24850_);
  and (_24857_, _24856_, _12013_);
  and (_24858_, _12012_, _05346_);
  or (_24859_, _24858_, _24857_);
  and (_24860_, _24859_, _05686_);
  nor (_24861_, _06633_, _05686_);
  nor (_24862_, _24861_, _12355_);
  not (_24863_, _24862_);
  nor (_24864_, _24863_, _24860_);
  not (_24866_, _05702_);
  nor (_24867_, _12351_, _05346_);
  nor (_24868_, _24867_, _24866_);
  not (_24869_, _24868_);
  nor (_24870_, _24869_, _24864_);
  nor (_24871_, _06633_, _05702_);
  and (_24872_, _12362_, _05675_);
  not (_24873_, _24872_);
  nor (_24874_, _24873_, _24871_);
  not (_24875_, _24874_);
  nor (_24877_, _24875_, _24870_);
  nor (_24878_, _24872_, _05346_);
  nor (_24879_, _24878_, _06023_);
  not (_24880_, _24879_);
  nor (_24881_, _24880_, _24877_);
  not (_24882_, _24774_);
  nor (_24883_, _06633_, _05673_);
  nor (_24884_, _24883_, _24882_);
  not (_24885_, _24884_);
  nor (_24886_, _24885_, _24881_);
  nor (_24888_, _24886_, _24775_);
  and (_24889_, _24888_, _05720_);
  nor (_24890_, _06633_, _05720_);
  or (_24891_, _24890_, _24889_);
  and (_24892_, _24891_, _12398_);
  and (_24893_, _24795_, _12397_);
  or (_24894_, _24893_, _24892_);
  and (_24895_, _24894_, _06020_);
  or (_24896_, _24895_, _24772_);
  and (_24897_, _24896_, _12413_);
  and (_24899_, _12412_, _05681_);
  or (_24900_, _24899_, _24897_);
  and (_24901_, _24900_, _13587_);
  nor (_24902_, _06633_, _13587_);
  or (_24903_, _24902_, _24901_);
  and (_24904_, _24903_, _12454_);
  not (_24905_, _24770_);
  nor (_24906_, _24795_, _11071_);
  and (_24907_, _11071_, _05346_);
  nor (_24908_, _24907_, _12454_);
  not (_24910_, _24908_);
  nor (_24911_, _24910_, _24906_);
  nor (_24912_, _24911_, _24905_);
  not (_24913_, _24912_);
  nor (_24914_, _24913_, _24904_);
  nor (_24915_, _24914_, _24771_);
  and (_24916_, _24915_, _24769_);
  nor (_24917_, _06633_, _24769_);
  or (_24918_, _24917_, _24916_);
  and (_24919_, _24918_, _12477_);
  not (_24921_, _24767_);
  nor (_24922_, _24795_, _12459_);
  nor (_24923_, _11071_, \oc8051_golden_model_1.PC [0]);
  nor (_24924_, _24923_, _12477_);
  not (_24925_, _24924_);
  nor (_24926_, _24925_, _24922_);
  nor (_24927_, _24926_, _24921_);
  not (_24928_, _24927_);
  nor (_24929_, _24928_, _24919_);
  nor (_24930_, _24929_, _24768_);
  and (_24932_, _24930_, _24765_);
  nor (_24933_, _06633_, _24765_);
  or (_24934_, _24933_, _24932_);
  and (_24935_, _24934_, _12498_);
  and (_24936_, _11993_, _08777_);
  not (_24937_, _24936_);
  or (_24938_, _24937_, _24935_);
  nor (_24939_, _24938_, _24764_);
  nor (_24940_, _24936_, _05346_);
  nor (_24941_, _24940_, _05740_);
  not (_24943_, _24941_);
  nor (_24944_, _24943_, _24939_);
  nor (_24945_, _24944_, _24760_);
  nor (_24946_, _24945_, _11982_);
  nor (_24947_, _10607_, _05346_);
  and (_24948_, _10607_, _05346_);
  nor (_24949_, _24948_, _24947_);
  nor (_24950_, _24949_, _12518_);
  nor (_24951_, _24950_, _24946_);
  and (_24952_, _24951_, _24758_);
  nor (_24954_, _24758_, _05346_);
  nor (_24955_, _24954_, _06298_);
  not (_24956_, _24955_);
  nor (_24957_, _24956_, _24952_);
  and (_24958_, _09120_, _06298_);
  or (_24959_, _24958_, _24957_);
  and (_24960_, _24959_, _05734_);
  nor (_24961_, _06633_, _05734_);
  or (_24962_, _24961_, _24960_);
  and (_24963_, _24962_, _06306_);
  and (_24965_, _24808_, _12722_);
  nor (_24966_, _12722_, _05346_);
  or (_24967_, _24966_, _06306_);
  or (_24968_, _24967_, _24965_);
  and (_24969_, _24968_, _24756_);
  not (_24970_, _24969_);
  nor (_24971_, _24970_, _24963_);
  nor (_24972_, _24971_, _24757_);
  and (_24973_, _24972_, _06050_);
  and (_24974_, _09120_, _06049_);
  or (_24976_, _24974_, _24973_);
  and (_24977_, _24976_, _05748_);
  nor (_24978_, _06633_, _05748_);
  nor (_24979_, _24978_, _24977_);
  nor (_24980_, _24979_, _06126_);
  not (_24981_, _24753_);
  and (_24982_, _12722_, \oc8051_golden_model_1.PC [0]);
  nor (_24983_, _24807_, _12722_);
  nor (_24984_, _24983_, _24982_);
  and (_24985_, _24984_, _06126_);
  nor (_24987_, _24985_, _24981_);
  not (_24988_, _24987_);
  nor (_24989_, _24988_, _24980_);
  nor (_24990_, _24989_, _24754_);
  nor (_24991_, _24990_, _07458_);
  and (_24992_, _07458_, _06633_);
  nor (_24993_, _24992_, _05652_);
  not (_24994_, _24993_);
  nor (_24995_, _24994_, _24991_);
  not (_24996_, _24751_);
  and (_24998_, _24984_, _05652_);
  nor (_24999_, _24998_, _24996_);
  not (_25000_, _24999_);
  nor (_25001_, _25000_, _24995_);
  nor (_25002_, _25001_, _24752_);
  nor (_25003_, _24749_, _25002_);
  or (_25004_, _25003_, _12789_);
  nor (_25005_, _25004_, _24750_);
  and (_25006_, _12789_, _05346_);
  or (_25007_, _25006_, _25005_);
  or (_25009_, _25007_, _01340_);
  or (_25010_, _01336_, \oc8051_golden_model_1.PC [0]);
  and (_25011_, _25010_, _42882_);
  and (_43417_, _25011_, _25009_);
  and (_25012_, _12789_, _12086_);
  and (_25013_, _06047_, _05312_);
  nor (_25014_, _12756_, _12086_);
  nor (_25015_, _08286_, _12086_);
  nor (_25016_, _11872_, _12086_);
  nor (_25017_, _12523_, _12086_);
  and (_25019_, _11989_, _05777_);
  nor (_25020_, _12002_, _12086_);
  and (_25021_, _12006_, _05777_);
  nor (_25022_, _08742_, _05312_);
  not (_25023_, _06089_);
  nor (_25024_, _12389_, _12086_);
  nor (_25025_, _12362_, _12086_);
  and (_25026_, _12172_, _05777_);
  nor (_25027_, _12090_, _12088_);
  nor (_25028_, _25027_, _12091_);
  and (_25030_, _25028_, _12174_);
  nor (_25031_, _25030_, _25026_);
  nand (_25032_, _25031_, _06104_);
  and (_25033_, _06948_, _12086_);
  or (_25034_, _12199_, \oc8051_golden_model_1.PC [1]);
  nor (_25035_, _11930_, _11928_);
  nor (_25036_, _25035_, _11931_);
  nand (_25037_, _25036_, _12199_);
  and (_25038_, _25037_, _25034_);
  nand (_25039_, _25038_, _08384_);
  and (_25041_, _06832_, _06943_);
  nor (_25042_, _12205_, _12086_);
  and (_25043_, _07250_, \oc8051_golden_model_1.PC [0]);
  nand (_25044_, _06450_, _06523_);
  and (_25045_, _06530_, _05346_);
  nor (_25046_, _25045_, _25044_);
  nor (_25047_, _25046_, _25043_);
  nor (_25048_, _25047_, _05312_);
  and (_25049_, _25047_, _05312_);
  nor (_25050_, _25049_, _25048_);
  nor (_25052_, _25050_, _24786_);
  nor (_25053_, _25052_, _25042_);
  not (_25054_, _25053_);
  nor (_25055_, _25054_, _25041_);
  nor (_25056_, _25055_, _08384_);
  nor (_25057_, _25056_, _06948_);
  and (_25058_, _25057_, _25039_);
  or (_25059_, _25058_, _25033_);
  nand (_25060_, _25059_, _06954_);
  or (_25061_, _12187_, _12086_);
  not (_25063_, _25028_);
  or (_25064_, _25063_, _12189_);
  nand (_25065_, _25064_, _25061_);
  nand (_25066_, _25065_, _06102_);
  and (_25067_, _25066_, _12182_);
  nand (_25068_, _25067_, _25060_);
  nor (_25069_, _12182_, _12086_);
  nor (_25070_, _25069_, _06043_);
  nand (_25071_, _25070_, _25068_);
  and (_25072_, _06043_, _05312_);
  nor (_25074_, _25072_, _07272_);
  nand (_25075_, _25074_, _25071_);
  and (_25076_, _06832_, _07272_);
  nor (_25077_, _25076_, _06239_);
  nand (_25078_, _25077_, _25075_);
  and (_25079_, _06239_, _05312_);
  nor (_25080_, _25079_, _12232_);
  nand (_25081_, _25080_, _25078_);
  nor (_25082_, _12231_, _12086_);
  nor (_25083_, _25082_, _06219_);
  nand (_25085_, _25083_, _25081_);
  and (_25086_, _06219_, _05312_);
  nor (_25087_, _25086_, _12241_);
  nand (_25088_, _25087_, _25085_);
  nor (_25089_, _12239_, _12086_);
  nor (_25090_, _25089_, _06039_);
  nand (_25091_, _25090_, _25088_);
  and (_25092_, _06039_, _05312_);
  nor (_25093_, _25092_, _12243_);
  nand (_25094_, _25093_, _25091_);
  and (_25096_, _06832_, _12243_);
  nor (_25097_, _25096_, _06038_);
  nand (_25098_, _25097_, _25094_);
  and (_25099_, _06038_, _05312_);
  nor (_25100_, _25099_, _12256_);
  and (_25101_, _25100_, _25098_);
  and (_25102_, _12289_, _05777_);
  nor (_25103_, _25063_, _12289_);
  or (_25104_, _25103_, _25102_);
  nor (_25105_, _25104_, _12255_);
  or (_25107_, _25105_, _25101_);
  nand (_25108_, _25107_, _12258_);
  nand (_25109_, _25108_, _25032_);
  nand (_25110_, _25109_, _06509_);
  nor (_25111_, _25063_, _12310_);
  not (_25112_, _25111_);
  and (_25113_, _12310_, _05777_);
  nor (_25114_, _25113_, _06509_);
  and (_25115_, _25114_, _25112_);
  nor (_25116_, _25115_, _06115_);
  nand (_25118_, _25116_, _25110_);
  and (_25119_, _12329_, _12086_);
  not (_25120_, _25119_);
  nor (_25121_, _25028_, _12329_);
  nor (_25122_, _25121_, _12298_);
  and (_25123_, _25122_, _25120_);
  nor (_25124_, _25123_, _12012_);
  nand (_25125_, _25124_, _25118_);
  and (_25126_, _12012_, _05777_);
  not (_25127_, _25126_);
  and (_25129_, _25127_, _12337_);
  nand (_25130_, _25129_, _25125_);
  and (_25131_, _06032_, _05312_);
  not (_25132_, _25131_);
  not (_25133_, _12344_);
  nor (_25134_, _06832_, _05686_);
  nor (_25135_, _25134_, _25133_);
  and (_25136_, _25135_, _25132_);
  nand (_25137_, _25136_, _25130_);
  nor (_25138_, _12344_, _05312_);
  nor (_25140_, _25138_, _12348_);
  nand (_25141_, _25140_, _25137_);
  and (_25142_, _12350_, _05777_);
  or (_25143_, _25142_, _12351_);
  nand (_25144_, _25143_, _25141_);
  nor (_25145_, _12350_, _12086_);
  nor (_25146_, _25145_, _06251_);
  nand (_25147_, _25146_, _25144_);
  and (_25148_, _06251_, _05312_);
  nor (_25149_, _25148_, _24866_);
  nand (_25150_, _25149_, _25147_);
  and (_25151_, _06832_, _24866_);
  nor (_25152_, _25151_, _06250_);
  nand (_25153_, _25152_, _25150_);
  and (_25154_, _06250_, _05312_);
  nor (_25155_, _25154_, _12368_);
  and (_25156_, _25155_, _25153_);
  or (_25157_, _25156_, _25025_);
  nand (_25158_, _25157_, _12366_);
  nor (_25159_, _12366_, _05312_);
  nor (_25162_, _25159_, _05676_);
  nand (_25163_, _25162_, _25158_);
  nor (_25164_, _05777_, _05675_);
  nor (_25165_, _25164_, _06026_);
  and (_25166_, _25165_, _25163_);
  and (_25167_, _06026_, \oc8051_golden_model_1.PC [1]);
  or (_25168_, _25167_, _25166_);
  nand (_25169_, _25168_, _05673_);
  and (_25170_, _06832_, _06023_);
  nor (_25171_, _25170_, _06110_);
  nand (_25173_, _25171_, _25169_);
  and (_25174_, _06110_, _05777_);
  nor (_25175_, _25174_, _09818_);
  nand (_25176_, _25175_, _25173_);
  nor (_25177_, _09817_, _05312_);
  nor (_25178_, _25177_, _09833_);
  nand (_25179_, _25178_, _25176_);
  nor (_25180_, _12086_, _05669_);
  nor (_25181_, _25180_, _12393_);
  and (_25182_, _25181_, _25179_);
  or (_25184_, _25182_, _25024_);
  nand (_25185_, _25184_, _25023_);
  and (_25186_, _06089_, \oc8051_golden_model_1.PC [1]);
  nor (_25187_, _25186_, _05719_);
  and (_25188_, _25187_, _25185_);
  nor (_25189_, _06832_, _05720_);
  or (_25190_, _25189_, _25188_);
  nand (_25191_, _25190_, _12398_);
  and (_25192_, _25036_, _12397_);
  nor (_25193_, _25192_, _08743_);
  and (_25195_, _25193_, _25191_);
  or (_25196_, _25195_, _25022_);
  nand (_25197_, _25196_, _06020_);
  and (_25198_, _06019_, _12086_);
  nor (_25199_, _25198_, _10661_);
  nand (_25200_, _25199_, _25197_);
  and (_25201_, _10661_, _05312_);
  nor (_25202_, _25201_, _12412_);
  nand (_25203_, _25202_, _25200_);
  nor (_25204_, _12413_, _05775_);
  nor (_25206_, _25204_, _06088_);
  nand (_25207_, _25206_, _25203_);
  and (_25208_, _06088_, _05312_);
  nor (_25209_, _25208_, _05724_);
  nand (_25210_, _25209_, _25207_);
  and (_25211_, _06832_, _05724_);
  nor (_25212_, _25211_, _12453_);
  nand (_25213_, _25212_, _25210_);
  nor (_25214_, _25036_, _11071_);
  and (_25215_, _11071_, \oc8051_golden_model_1.PC [1]);
  nor (_25217_, _25215_, _12454_);
  not (_25218_, _25217_);
  nor (_25219_, _25218_, _25214_);
  nor (_25220_, _25219_, _12006_);
  and (_25221_, _25220_, _25213_);
  or (_25222_, _25221_, _25021_);
  nand (_25223_, _25222_, _12466_);
  nor (_25224_, _12466_, _05312_);
  nor (_25225_, _25224_, _06112_);
  nand (_25226_, _25225_, _25223_);
  and (_25228_, _06112_, _05777_);
  nor (_25229_, _25228_, _06284_);
  and (_25230_, _25229_, _25226_);
  and (_25231_, _06284_, \oc8051_golden_model_1.PC [1]);
  or (_25232_, _25231_, _25230_);
  nand (_25233_, _25232_, _24769_);
  and (_25234_, _06832_, _05727_);
  nor (_25235_, _25234_, _12476_);
  nand (_25236_, _25235_, _25233_);
  nor (_25237_, _25036_, _12459_);
  nor (_25239_, _11071_, _05312_);
  nor (_25240_, _25239_, _12477_);
  not (_25241_, _25240_);
  nor (_25242_, _25241_, _25237_);
  nor (_25243_, _25242_, _12481_);
  and (_25244_, _25243_, _25236_);
  or (_25245_, _25244_, _25020_);
  nand (_25246_, _25245_, _10742_);
  nor (_25247_, _10742_, _05312_);
  nor (_25248_, _25247_, _06108_);
  nand (_25250_, _25248_, _25246_);
  and (_25251_, _06108_, _05777_);
  nor (_25252_, _25251_, _06277_);
  and (_25253_, _25252_, _25250_);
  and (_25254_, _06277_, \oc8051_golden_model_1.PC [1]);
  or (_25255_, _25254_, _25253_);
  nand (_25256_, _25255_, _24765_);
  and (_25257_, _06832_, _05736_);
  nor (_25258_, _25257_, _12497_);
  nand (_25259_, _25258_, _25256_);
  and (_25261_, \oc8051_golden_model_1.PSW [7], _05312_);
  and (_25262_, _25036_, _10606_);
  or (_25263_, _25262_, _25261_);
  and (_25264_, _25263_, _12497_);
  nor (_25265_, _25264_, _11989_);
  and (_25266_, _25265_, _25259_);
  nor (_25267_, _25266_, _25019_);
  nor (_25268_, _07002_, _10394_);
  nor (_25269_, _25268_, _10757_);
  or (_25270_, _25269_, _25267_);
  and (_25272_, _25269_, _05777_);
  nor (_25273_, _25272_, _06669_);
  nand (_25274_, _25273_, _25270_);
  and (_25275_, _06669_, _12086_);
  nor (_25276_, _25275_, _11987_);
  nand (_25277_, _25276_, _25274_);
  nor (_25278_, _11986_, _05312_);
  nor (_25279_, _25278_, _06130_);
  and (_25280_, _25279_, _25277_);
  and (_25281_, _06130_, _05777_);
  or (_25283_, _25281_, _06292_);
  nor (_25284_, _25283_, _25280_);
  and (_25285_, _06292_, \oc8051_golden_model_1.PC [1]);
  or (_25286_, _25285_, _25284_);
  nand (_25287_, _25286_, _24759_);
  and (_25288_, _06832_, _05740_);
  nor (_25289_, _25288_, _11982_);
  nand (_25290_, _25289_, _25287_);
  nor (_25291_, _25036_, _10606_);
  and (_25292_, _10606_, \oc8051_golden_model_1.PC [1]);
  nor (_25294_, _25292_, _12518_);
  not (_25295_, _25294_);
  nor (_25296_, _25295_, _25291_);
  nor (_25297_, _25296_, _12525_);
  and (_25298_, _25297_, _25290_);
  or (_25299_, _25298_, _25017_);
  nand (_25300_, _25299_, _10825_);
  nor (_25301_, _10825_, _05312_);
  nor (_25302_, _25301_, _10854_);
  nand (_25303_, _25302_, _25300_);
  and (_25305_, _10854_, _12086_);
  nor (_25306_, _25305_, _06298_);
  and (_25307_, _25306_, _25303_);
  and (_25308_, _12150_, _06298_);
  or (_25309_, _25308_, _25307_);
  nand (_25310_, _25309_, _05734_);
  and (_25311_, _06832_, _05732_);
  nor (_25312_, _25311_, _06129_);
  nand (_25313_, _25312_, _25310_);
  nor (_25314_, _12722_, _05777_);
  not (_25316_, _25314_);
  and (_25317_, _25063_, _12722_);
  nor (_25318_, _25317_, _06306_);
  and (_25319_, _25318_, _25316_);
  nor (_25320_, _25319_, _12541_);
  and (_25321_, _25320_, _25313_);
  or (_25322_, _25321_, _25016_);
  nand (_25323_, _25322_, _10975_);
  nor (_25324_, _10975_, _05312_);
  nor (_25325_, _25324_, _11015_);
  nand (_25327_, _25325_, _25323_);
  and (_25328_, _11015_, _12086_);
  nor (_25329_, _25328_, _06049_);
  and (_25330_, _25329_, _25327_);
  and (_25331_, _12150_, _06049_);
  or (_25332_, _25331_, _25330_);
  nand (_25333_, _25332_, _05748_);
  and (_25334_, _06832_, _05747_);
  nor (_25335_, _25334_, _06126_);
  nand (_25336_, _25335_, _25333_);
  not (_25338_, _08286_);
  nor (_25339_, _25028_, _12722_);
  and (_25340_, _12722_, _12086_);
  nor (_25341_, _25340_, _25339_);
  and (_25342_, _25341_, _06126_);
  nor (_25343_, _25342_, _25338_);
  and (_25344_, _25343_, _25336_);
  nor (_25345_, _25344_, _25015_);
  not (_25346_, _05495_);
  nor (_25347_, _07248_, _25346_);
  or (_25349_, _25347_, _25345_);
  and (_25350_, _25347_, _05777_);
  nor (_25351_, _25350_, _06316_);
  nand (_25352_, _25351_, _25349_);
  not (_25353_, _12756_);
  and (_25354_, _06316_, _05312_);
  nor (_25355_, _25354_, _25353_);
  and (_25356_, _25355_, _25352_);
  or (_25357_, _25356_, _25014_);
  nand (_25358_, _25357_, _07059_);
  and (_25360_, _07458_, _06832_);
  nor (_25361_, _25360_, _05652_);
  nand (_25362_, _25361_, _25358_);
  and (_25363_, _25341_, _05652_);
  nor (_25364_, _25363_, _12772_);
  nand (_25365_, _25364_, _25362_);
  nor (_25366_, _12771_, _12086_);
  nor (_25367_, _25366_, _06047_);
  and (_25368_, _25367_, _25365_);
  or (_25369_, _25368_, _25013_);
  nand (_25371_, _25369_, _12779_);
  nor (_25372_, _12779_, _05777_);
  nor (_25373_, _25372_, _24749_);
  nand (_25374_, _25373_, _25371_);
  and (_25375_, _24749_, _06832_);
  nor (_25376_, _25375_, _12789_);
  and (_25377_, _25376_, _25374_);
  or (_25378_, _25377_, _25012_);
  or (_25379_, _25378_, _01340_);
  or (_25380_, _01336_, \oc8051_golden_model_1.PC [1]);
  and (_25382_, _25380_, _42882_);
  and (_43418_, _25382_, _25379_);
  and (_25383_, _06047_, _05803_);
  and (_25384_, _06316_, _05803_);
  nor (_25385_, _11872_, _05823_);
  nor (_25386_, _12523_, _05823_);
  nor (_25387_, _11993_, _05823_);
  nor (_25388_, _12002_, _05823_);
  and (_25389_, _12006_, _05824_);
  nor (_25390_, _08741_, _05803_);
  nor (_25392_, _12344_, _05803_);
  and (_25393_, _12012_, _05824_);
  or (_25394_, _12174_, _12083_);
  and (_25395_, _12095_, _12092_);
  nor (_25396_, _25395_, _12096_);
  or (_25397_, _25396_, _12172_);
  nand (_25398_, _25397_, _25394_);
  nand (_25399_, _25398_, _06104_);
  and (_25400_, _06943_, _06445_);
  nor (_25401_, _12205_, _05823_);
  nor (_25403_, _12214_, _05823_);
  and (_25404_, _06938_, _05804_);
  nor (_25405_, _06938_, \oc8051_golden_model_1.PC [2]);
  and (_25406_, _25405_, _07251_);
  nor (_25407_, _25406_, _25404_);
  nor (_25408_, _25407_, _06530_);
  nor (_25409_, _25408_, _25403_);
  nor (_25410_, _25409_, _24786_);
  or (_25411_, _25410_, _25401_);
  nor (_25412_, _25411_, _25400_);
  nor (_25413_, _25412_, _08384_);
  and (_25414_, _11935_, _11932_);
  nor (_25415_, _25414_, _11936_);
  nand (_25416_, _25415_, _12199_);
  or (_25417_, _12199_, _05804_);
  and (_25418_, _25417_, _08384_);
  and (_25419_, _25418_, _25416_);
  or (_25420_, _25419_, _25413_);
  nand (_25421_, _25420_, _06949_);
  and (_25422_, _06948_, _05824_);
  nor (_25425_, _25422_, _06102_);
  nand (_25426_, _25425_, _25421_);
  or (_25427_, _25396_, _12189_);
  or (_25428_, _12187_, _12083_);
  and (_25429_, _25428_, _06102_);
  nand (_25430_, _25429_, _25427_);
  and (_25431_, _25430_, _12182_);
  nand (_25432_, _25431_, _25426_);
  nor (_25433_, _12182_, _05823_);
  nor (_25434_, _25433_, _06043_);
  nand (_25436_, _25434_, _25432_);
  and (_25437_, _06043_, _05803_);
  nor (_25438_, _25437_, _07272_);
  nand (_25439_, _25438_, _25436_);
  and (_25440_, _06445_, _07272_);
  nor (_25441_, _25440_, _06239_);
  nand (_25442_, _25441_, _25439_);
  and (_25443_, _06239_, _05803_);
  nor (_25444_, _25443_, _12232_);
  nand (_25445_, _25444_, _25442_);
  nor (_25447_, _12231_, _05823_);
  nor (_25448_, _25447_, _06219_);
  nand (_25449_, _25448_, _25445_);
  and (_25450_, _06219_, _05803_);
  nor (_25451_, _25450_, _12241_);
  nand (_25452_, _25451_, _25449_);
  nor (_25453_, _12239_, _05823_);
  nor (_25454_, _25453_, _06039_);
  nand (_25455_, _25454_, _25452_);
  and (_25456_, _06039_, _05803_);
  nor (_25458_, _25456_, _12243_);
  nand (_25459_, _25458_, _25455_);
  and (_25460_, _06445_, _12243_);
  nor (_25461_, _25460_, _06038_);
  nand (_25462_, _25461_, _25459_);
  and (_25463_, _06038_, _05803_);
  nor (_25464_, _25463_, _12256_);
  and (_25465_, _25464_, _25462_);
  and (_25466_, _12289_, _12083_);
  not (_25467_, _25466_);
  not (_25469_, _25396_);
  nor (_25470_, _25469_, _12289_);
  nor (_25471_, _25470_, _12255_);
  and (_25472_, _25471_, _25467_);
  or (_25473_, _25472_, _25465_);
  nand (_25474_, _25473_, _12258_);
  nand (_25475_, _25474_, _25399_);
  nand (_25476_, _25475_, _06509_);
  nor (_25477_, _25469_, _12310_);
  not (_25478_, _25477_);
  and (_25480_, _12310_, _12083_);
  nor (_25481_, _25480_, _06509_);
  and (_25482_, _25481_, _25478_);
  nor (_25483_, _25482_, _06115_);
  nand (_25484_, _25483_, _25476_);
  and (_25485_, _12329_, _12084_);
  nor (_25486_, _25396_, _12329_);
  or (_25487_, _25486_, _12298_);
  or (_25488_, _25487_, _25485_);
  and (_25489_, _25488_, _12013_);
  and (_25491_, _25489_, _25484_);
  or (_25492_, _25491_, _25393_);
  nand (_25493_, _25492_, _06033_);
  and (_25494_, _06032_, _05804_);
  nor (_25495_, _25494_, _07355_);
  nand (_25496_, _25495_, _25493_);
  nor (_25497_, _06445_, _05686_);
  nor (_25498_, _25497_, _25133_);
  and (_25499_, _25498_, _25496_);
  or (_25500_, _25499_, _25392_);
  nand (_25502_, _25500_, _12351_);
  nor (_25503_, _12351_, _05823_);
  nor (_25504_, _25503_, _06251_);
  nand (_25505_, _25504_, _25502_);
  and (_25506_, _06251_, _05803_);
  nor (_25507_, _25506_, _24866_);
  nand (_25508_, _25507_, _25505_);
  and (_25509_, _06445_, _24866_);
  nor (_25510_, _25509_, _06250_);
  nand (_25511_, _25510_, _25508_);
  and (_25513_, _06250_, _05803_);
  nor (_25514_, _25513_, _12368_);
  and (_25515_, _25514_, _25511_);
  nor (_25516_, _12362_, _05823_);
  or (_25517_, _25516_, _25515_);
  nand (_25518_, _25517_, _12366_);
  nor (_25519_, _12366_, _05803_);
  nor (_25520_, _25519_, _05676_);
  nand (_25521_, _25520_, _25518_);
  nor (_25522_, _05824_, _05675_);
  nor (_25524_, _25522_, _06026_);
  and (_25525_, _25524_, _25521_);
  and (_25526_, _06026_, _05804_);
  or (_25527_, _25526_, _25525_);
  nand (_25528_, _25527_, _05673_);
  and (_25529_, _06445_, _06023_);
  nor (_25530_, _25529_, _06110_);
  nand (_25531_, _25530_, _25528_);
  and (_25532_, _12083_, _06110_);
  nor (_25533_, _25532_, _07011_);
  and (_25535_, _25533_, _09827_);
  nand (_25536_, _25535_, _25531_);
  nor (_25537_, _09817_, _05803_);
  nor (_25538_, _25537_, _09833_);
  nand (_25539_, _25538_, _25536_);
  nor (_25540_, _12084_, _05669_);
  nor (_25541_, _25540_, _12393_);
  nand (_25542_, _25541_, _25539_);
  nor (_25543_, _12389_, _05823_);
  nor (_25544_, _25543_, _06089_);
  and (_25546_, _25544_, _25542_);
  and (_25547_, _06089_, _05803_);
  or (_25548_, _25547_, _05719_);
  nor (_25549_, _25548_, _25546_);
  and (_25550_, _06445_, _05719_);
  or (_25551_, _25550_, _25549_);
  nand (_25552_, _25551_, _12398_);
  not (_25553_, _08740_);
  nor (_25554_, _25415_, _12398_);
  nor (_25555_, _25554_, _25553_);
  nand (_25557_, _25555_, _25552_);
  not (_25558_, _08741_);
  nor (_25559_, _08740_, _05804_);
  nor (_25560_, _25559_, _25558_);
  and (_25561_, _25560_, _25557_);
  or (_25562_, _25561_, _25390_);
  nand (_25563_, _25562_, _06020_);
  and (_25564_, _12084_, _06019_);
  nor (_25565_, _25564_, _10661_);
  nand (_25566_, _25565_, _25563_);
  and (_25568_, _10661_, _05803_);
  nor (_25569_, _25568_, _12412_);
  nand (_25570_, _25569_, _25566_);
  and (_25571_, _12412_, _05818_);
  nor (_25572_, _25571_, _06088_);
  nand (_25573_, _25572_, _25570_);
  and (_25574_, _06088_, _05803_);
  nor (_25575_, _25574_, _05724_);
  nand (_25576_, _25575_, _25573_);
  and (_25577_, _06445_, _05724_);
  nor (_25579_, _25577_, _12453_);
  nand (_25580_, _25579_, _25576_);
  nor (_25581_, _25415_, _11071_);
  and (_25582_, _11071_, _05804_);
  nor (_25583_, _25582_, _12454_);
  not (_25584_, _25583_);
  nor (_25585_, _25584_, _25581_);
  nor (_25586_, _25585_, _12006_);
  and (_25587_, _25586_, _25580_);
  or (_25588_, _25587_, _25389_);
  nand (_25590_, _25588_, _12466_);
  nor (_25591_, _12466_, _05803_);
  nor (_25592_, _25591_, _06112_);
  nand (_25593_, _25592_, _25590_);
  and (_25594_, _12083_, _06112_);
  nor (_25595_, _25594_, _06284_);
  and (_25596_, _25595_, _25593_);
  and (_25597_, _06284_, _05804_);
  or (_25598_, _25597_, _25596_);
  nand (_25599_, _25598_, _24769_);
  and (_25601_, _06445_, _05727_);
  nor (_25602_, _25601_, _12476_);
  nand (_25603_, _25602_, _25599_);
  nor (_25604_, _25415_, _12459_);
  nor (_25605_, _11071_, _05803_);
  nor (_25606_, _25605_, _12477_);
  not (_25607_, _25606_);
  nor (_25608_, _25607_, _25604_);
  nor (_25609_, _25608_, _12481_);
  and (_25610_, _25609_, _25603_);
  or (_25612_, _25610_, _25388_);
  nand (_25613_, _25612_, _10742_);
  nor (_25614_, _10742_, _05803_);
  nor (_25615_, _25614_, _06108_);
  nand (_25616_, _25615_, _25613_);
  and (_25617_, _12083_, _06108_);
  nor (_25618_, _25617_, _06277_);
  and (_25619_, _25618_, _25616_);
  and (_25620_, _06277_, _05804_);
  or (_25621_, _25620_, _25619_);
  nand (_25623_, _25621_, _24765_);
  and (_25624_, _06445_, _05736_);
  nor (_25625_, _25624_, _12497_);
  nand (_25626_, _25625_, _25623_);
  nor (_25627_, _25415_, \oc8051_golden_model_1.PSW [7]);
  nor (_25628_, _05803_, _10606_);
  nor (_25629_, _25628_, _12498_);
  not (_25630_, _25629_);
  nor (_25631_, _25630_, _25627_);
  nor (_25632_, _25631_, _12502_);
  and (_25634_, _25632_, _25626_);
  or (_25635_, _25634_, _25387_);
  nand (_25636_, _25635_, _11986_);
  nor (_25637_, _11986_, _05803_);
  nor (_25638_, _25637_, _06130_);
  and (_25639_, _25638_, _25636_);
  and (_25640_, _12083_, _06130_);
  or (_25641_, _25640_, _06292_);
  nor (_25642_, _25641_, _25639_);
  and (_25643_, _06292_, _05804_);
  or (_25645_, _25643_, _25642_);
  nand (_25646_, _25645_, _24759_);
  and (_25647_, _06445_, _05740_);
  nor (_25648_, _25647_, _11982_);
  nand (_25649_, _25648_, _25646_);
  or (_25650_, _25415_, _10606_);
  or (_25651_, _05803_, \oc8051_golden_model_1.PSW [7]);
  and (_25652_, _25651_, _11982_);
  and (_25653_, _25652_, _25650_);
  nor (_25654_, _25653_, _12525_);
  and (_25656_, _25654_, _25649_);
  or (_25657_, _25656_, _25386_);
  nand (_25658_, _25657_, _10825_);
  nor (_25659_, _10825_, _05803_);
  nor (_25660_, _25659_, _10854_);
  nand (_25661_, _25660_, _25658_);
  and (_25662_, _10854_, _05823_);
  nor (_25663_, _25662_, _06298_);
  and (_25664_, _25663_, _25661_);
  and (_25665_, _09030_, _06298_);
  or (_25667_, _25665_, _25664_);
  nand (_25668_, _25667_, _05734_);
  and (_25669_, _06445_, _05732_);
  nor (_25670_, _25669_, _06129_);
  nand (_25671_, _25670_, _25668_);
  nor (_25672_, _12083_, _12722_);
  and (_25673_, _25469_, _12722_);
  or (_25674_, _25673_, _06306_);
  nor (_25675_, _25674_, _25672_);
  nor (_25676_, _25675_, _12541_);
  and (_25678_, _25676_, _25671_);
  or (_25679_, _25678_, _25385_);
  nand (_25680_, _25679_, _10975_);
  nor (_25681_, _10975_, _05803_);
  nor (_25682_, _25681_, _11015_);
  nand (_25683_, _25682_, _25680_);
  and (_25684_, _11015_, _05823_);
  nor (_25685_, _25684_, _06049_);
  and (_25686_, _25685_, _25683_);
  and (_25687_, _09030_, _06049_);
  or (_25689_, _25687_, _25686_);
  nand (_25690_, _25689_, _05748_);
  and (_25691_, _06445_, _05747_);
  nor (_25692_, _25691_, _06126_);
  nand (_25693_, _25692_, _25690_);
  nor (_25694_, _25396_, _12722_);
  and (_25695_, _12084_, _12722_);
  nor (_25696_, _25695_, _25694_);
  and (_25697_, _25696_, _06126_);
  nor (_25698_, _25697_, _12750_);
  nand (_25700_, _25698_, _25693_);
  nor (_25701_, _12749_, _05823_);
  nor (_25702_, _25701_, _06316_);
  and (_25703_, _25702_, _25700_);
  or (_25704_, _25703_, _25384_);
  nand (_25705_, _25704_, _12756_);
  nor (_25706_, _12756_, _05824_);
  nor (_25707_, _25706_, _07458_);
  nand (_25708_, _25707_, _25705_);
  and (_25709_, _07458_, _06445_);
  nor (_25711_, _25709_, _05652_);
  nand (_25712_, _25711_, _25708_);
  and (_25713_, _25696_, _05652_);
  nor (_25714_, _25713_, _12772_);
  nand (_25715_, _25714_, _25712_);
  nor (_25716_, _12771_, _05823_);
  nor (_25717_, _25716_, _06047_);
  and (_25718_, _25717_, _25715_);
  or (_25719_, _25718_, _25383_);
  nand (_25720_, _25719_, _12779_);
  nor (_25721_, _12779_, _05824_);
  nor (_25722_, _25721_, _24749_);
  nand (_25723_, _25722_, _25720_);
  and (_25724_, _24749_, _06445_);
  nor (_25725_, _25724_, _12789_);
  and (_25726_, _25725_, _25723_);
  and (_25727_, _12789_, _05823_);
  or (_25728_, _25727_, _25726_);
  or (_25729_, _25728_, _01340_);
  or (_25730_, _01336_, \oc8051_golden_model_1.PC [2]);
  and (_25733_, _25730_, _42882_);
  and (_43419_, _25733_, _25729_);
  and (_25734_, _06047_, _05853_);
  nor (_25735_, _11872_, _06150_);
  nor (_25736_, _12523_, _06150_);
  or (_25737_, _11993_, _06150_);
  or (_25738_, _12002_, _06150_);
  nand (_25739_, _12006_, _05870_);
  or (_25740_, _08742_, _05853_);
  nand (_25741_, _12012_, _05870_);
  and (_25743_, _12172_, _12078_);
  or (_25744_, _12081_, _12080_);
  and (_25745_, _25744_, _12097_);
  nor (_25746_, _25744_, _12097_);
  nor (_25747_, _25746_, _25745_);
  and (_25748_, _25747_, _12174_);
  or (_25749_, _25748_, _25743_);
  or (_25750_, _25749_, _12258_);
  and (_25751_, _12289_, _12078_);
  not (_25752_, _25747_);
  nor (_25754_, _25752_, _12289_);
  or (_25755_, _25754_, _25751_);
  or (_25756_, _25755_, _12255_);
  nor (_25757_, _07233_, _06215_);
  not (_25758_, _06530_);
  nand (_25759_, _06938_, _06148_);
  and (_25760_, _25759_, _25758_);
  nor (_25761_, _07250_, _05307_);
  or (_25762_, _25761_, _06938_);
  and (_25763_, _25762_, _25760_);
  or (_25765_, _12214_, _05870_);
  nand (_25766_, _25765_, _12205_);
  or (_25767_, _25766_, _25763_);
  and (_25768_, _25767_, _07233_);
  or (_25769_, _25768_, _25757_);
  or (_25770_, _12205_, _06150_);
  and (_25771_, _25770_, _25769_);
  or (_25772_, _25771_, _08384_);
  or (_25773_, _11925_, _11924_);
  and (_25774_, _25773_, _11937_);
  nor (_25776_, _25773_, _11937_);
  nor (_25777_, _25776_, _25774_);
  and (_25778_, _25777_, _12199_);
  and (_25779_, _12197_, _05853_);
  or (_25780_, _25779_, _08383_);
  or (_25781_, _25780_, _25778_);
  and (_25782_, _25781_, _25772_);
  or (_25783_, _25782_, _06948_);
  nand (_25784_, _06948_, _05870_);
  and (_25785_, _25784_, _06954_);
  and (_25787_, _25785_, _25783_);
  or (_25788_, _12187_, _12078_);
  or (_25789_, _25747_, _12189_);
  and (_25790_, _25789_, _06102_);
  and (_25791_, _25790_, _25788_);
  or (_25792_, _25791_, _24805_);
  or (_25793_, _25792_, _25787_);
  or (_25794_, _12182_, _06150_);
  and (_25795_, _25794_, _06044_);
  and (_25796_, _25795_, _25793_);
  and (_25798_, _06043_, _05853_);
  or (_25799_, _25798_, _07272_);
  or (_25800_, _25799_, _25796_);
  nand (_25801_, _06215_, _07272_);
  and (_25802_, _25801_, _06848_);
  and (_25803_, _25802_, _25800_);
  nand (_25804_, _06239_, _05853_);
  nand (_25805_, _25804_, _12231_);
  or (_25806_, _25805_, _25803_);
  or (_25807_, _12231_, _06150_);
  and (_25809_, _25807_, _06220_);
  and (_25810_, _25809_, _25806_);
  nand (_25811_, _06219_, _05853_);
  nand (_25812_, _25811_, _12239_);
  or (_25813_, _25812_, _25810_);
  or (_25814_, _12239_, _06150_);
  and (_25815_, _25814_, _06040_);
  and (_25816_, _25815_, _25813_);
  and (_25817_, _06039_, _05853_);
  or (_25818_, _25817_, _12243_);
  or (_25820_, _25818_, _25816_);
  nand (_25821_, _06215_, _12243_);
  and (_25822_, _25821_, _07364_);
  and (_25823_, _25822_, _25820_);
  nand (_25824_, _06038_, _05853_);
  nand (_25825_, _25824_, _12255_);
  or (_25826_, _25825_, _25823_);
  and (_25827_, _25826_, _25756_);
  or (_25828_, _25827_, _13850_);
  and (_25829_, _25828_, _25750_);
  or (_25831_, _25829_, _06121_);
  nor (_25832_, _25752_, _12310_);
  and (_25833_, _12310_, _12078_);
  or (_25834_, _25833_, _06509_);
  or (_25835_, _25834_, _25832_);
  and (_25836_, _25835_, _12298_);
  and (_25837_, _25836_, _25831_);
  nand (_25838_, _12329_, _12079_);
  or (_25839_, _25747_, _12329_);
  and (_25840_, _25839_, _06115_);
  and (_25842_, _25840_, _25838_);
  or (_25843_, _25842_, _12012_);
  or (_25844_, _25843_, _25837_);
  and (_25845_, _25844_, _25741_);
  or (_25846_, _25845_, _06032_);
  nand (_25847_, _06032_, _06148_);
  and (_25848_, _25847_, _05686_);
  and (_25849_, _25848_, _25846_);
  nor (_25850_, _06215_, _05686_);
  or (_25851_, _25850_, _25133_);
  or (_25853_, _25851_, _25849_);
  or (_25854_, _12344_, _05853_);
  and (_25855_, _25854_, _25853_);
  or (_25856_, _25855_, _12355_);
  or (_25857_, _12351_, _06150_);
  and (_25858_, _25857_, _13765_);
  and (_25859_, _25858_, _25856_);
  and (_25860_, _06251_, _05853_);
  or (_25861_, _25860_, _24866_);
  or (_25862_, _25861_, _25859_);
  nand (_25864_, _06215_, _24866_);
  and (_25865_, _25864_, _13764_);
  and (_25866_, _25865_, _25862_);
  nand (_25867_, _06250_, _05853_);
  nand (_25868_, _25867_, _12362_);
  or (_25869_, _25868_, _25866_);
  or (_25870_, _12362_, _06150_);
  and (_25871_, _25870_, _25869_);
  or (_25872_, _25871_, _12367_);
  or (_25873_, _12366_, _05853_);
  and (_25875_, _25873_, _05675_);
  and (_25876_, _25875_, _25872_);
  nor (_25877_, _05675_, _05870_);
  or (_25878_, _25877_, _06026_);
  or (_25879_, _25878_, _25876_);
  nand (_25880_, _06026_, _06148_);
  and (_25881_, _25880_, _25879_);
  or (_25882_, _25881_, _06023_);
  nand (_25883_, _06215_, _06023_);
  and (_25884_, _25883_, _06111_);
  and (_25886_, _25884_, _25882_);
  nand (_25887_, _12078_, _06110_);
  nand (_25888_, _25887_, _09817_);
  or (_25889_, _25888_, _25886_);
  or (_25890_, _09817_, _05853_);
  and (_25891_, _25890_, _05669_);
  and (_25892_, _25891_, _25889_);
  or (_25893_, _12079_, _05669_);
  nand (_25894_, _25893_, _12389_);
  or (_25895_, _25894_, _25892_);
  or (_25896_, _12389_, _06150_);
  and (_25897_, _25896_, _25023_);
  and (_25898_, _25897_, _25895_);
  and (_25899_, _06089_, _05853_);
  or (_25900_, _25899_, _05719_);
  or (_25901_, _25900_, _25898_);
  nand (_25902_, _06215_, _05719_);
  and (_25903_, _25902_, _12398_);
  and (_25904_, _25903_, _25901_);
  and (_25905_, _25777_, _12397_);
  or (_25907_, _25905_, _08743_);
  or (_25908_, _25907_, _25904_);
  and (_25909_, _25908_, _25740_);
  or (_25910_, _25909_, _06019_);
  nand (_25911_, _12079_, _06019_);
  and (_25912_, _25911_, _10662_);
  and (_25913_, _25912_, _25910_);
  and (_25914_, _10661_, _05853_);
  or (_25915_, _25914_, _12412_);
  or (_25916_, _25915_, _25913_);
  or (_25918_, _12413_, _05865_);
  and (_25919_, _25918_, _06636_);
  and (_25920_, _25919_, _25916_);
  and (_25921_, _06088_, _05853_);
  or (_25922_, _25921_, _05724_);
  or (_25923_, _25922_, _25920_);
  nand (_25924_, _06215_, _05724_);
  and (_25925_, _25924_, _12454_);
  and (_25926_, _25925_, _25923_);
  or (_25927_, _25777_, _11071_);
  nand (_25928_, _11071_, _06148_);
  and (_25929_, _25928_, _12453_);
  and (_25930_, _25929_, _25927_);
  or (_25931_, _25930_, _12006_);
  or (_25932_, _25931_, _25926_);
  and (_25933_, _25932_, _25739_);
  or (_25934_, _25933_, _12467_);
  or (_25935_, _12466_, _05853_);
  and (_25936_, _25935_, _08751_);
  and (_25937_, _25936_, _25934_);
  and (_25938_, _12078_, _06112_);
  or (_25939_, _25938_, _06284_);
  or (_25940_, _25939_, _25937_);
  nand (_25941_, _06284_, _06148_);
  and (_25942_, _25941_, _25940_);
  or (_25943_, _25942_, _05727_);
  nand (_25944_, _06215_, _05727_);
  and (_25945_, _25944_, _12477_);
  and (_25946_, _25945_, _25943_);
  or (_25947_, _25777_, _12459_);
  or (_25948_, _11071_, _05853_);
  and (_25949_, _25948_, _12476_);
  and (_25950_, _25949_, _25947_);
  or (_25951_, _25950_, _12481_);
  or (_25952_, _25951_, _25946_);
  and (_25953_, _25952_, _25738_);
  or (_25954_, _25953_, _10743_);
  or (_25955_, _10742_, _05853_);
  and (_25956_, _25955_, _07032_);
  and (_25957_, _25956_, _25954_);
  and (_25958_, _12078_, _06108_);
  or (_25959_, _25958_, _06277_);
  or (_25960_, _25959_, _25957_);
  nand (_25961_, _06277_, _06148_);
  and (_25962_, _25961_, _25960_);
  or (_25963_, _25962_, _05736_);
  nand (_25964_, _06215_, _05736_);
  and (_25965_, _25964_, _12498_);
  and (_25966_, _25965_, _25963_);
  or (_25967_, _25777_, \oc8051_golden_model_1.PSW [7]);
  or (_25968_, _05853_, _10606_);
  and (_25969_, _25968_, _12497_);
  and (_25970_, _25969_, _25967_);
  or (_25971_, _25970_, _12502_);
  or (_25972_, _25971_, _25966_);
  nand (_25973_, _25972_, _25737_);
  nand (_25974_, _25973_, _11986_);
  nor (_25975_, _11986_, _05853_);
  nor (_25976_, _25975_, _06130_);
  and (_25977_, _25976_, _25974_);
  and (_25979_, _12078_, _06130_);
  or (_25980_, _25979_, _06292_);
  nor (_25981_, _25980_, _25977_);
  and (_25982_, _06292_, _06148_);
  or (_25983_, _25982_, _25981_);
  nand (_25984_, _25983_, _24759_);
  and (_25985_, _06215_, _05740_);
  nor (_25986_, _25985_, _11982_);
  nand (_25987_, _25986_, _25984_);
  and (_25988_, _05853_, _10606_);
  and (_25990_, _25777_, \oc8051_golden_model_1.PSW [7]);
  or (_25991_, _25990_, _25988_);
  and (_25992_, _25991_, _11982_);
  nor (_25993_, _25992_, _12525_);
  and (_25994_, _25993_, _25987_);
  or (_25995_, _25994_, _25736_);
  nand (_25996_, _25995_, _10825_);
  nor (_25997_, _10825_, _05853_);
  nor (_25998_, _25997_, _10854_);
  nand (_25999_, _25998_, _25996_);
  and (_26000_, _10854_, _06150_);
  nor (_26001_, _26000_, _06298_);
  and (_26002_, _26001_, _25999_);
  and (_26003_, _08985_, _06298_);
  or (_26004_, _26003_, _26002_);
  nand (_26005_, _26004_, _05734_);
  and (_26006_, _06215_, _05732_);
  nor (_26007_, _26006_, _06129_);
  nand (_26008_, _26007_, _26005_);
  and (_26009_, _25752_, _12722_);
  nor (_26011_, _12078_, _12722_);
  or (_26012_, _26011_, _06306_);
  nor (_26013_, _26012_, _26009_);
  nor (_26014_, _26013_, _12541_);
  and (_26015_, _26014_, _26008_);
  or (_26016_, _26015_, _25735_);
  nand (_26017_, _26016_, _10975_);
  nor (_26018_, _10975_, _05853_);
  nor (_26019_, _26018_, _11015_);
  nand (_26020_, _26019_, _26017_);
  and (_26022_, _11015_, _06150_);
  nor (_26023_, _26022_, _06049_);
  and (_26024_, _26023_, _26020_);
  and (_26025_, _08985_, _06049_);
  or (_26026_, _26025_, _26024_);
  nand (_26027_, _26026_, _05748_);
  and (_26028_, _06215_, _05747_);
  nor (_26029_, _26028_, _06126_);
  nand (_26030_, _26029_, _26027_);
  nor (_26031_, _25747_, _12722_);
  and (_26033_, _12079_, _12722_);
  nor (_26034_, _26033_, _26031_);
  and (_26035_, _26034_, _06126_);
  nor (_26036_, _26035_, _12750_);
  nand (_26037_, _26036_, _26030_);
  nor (_26038_, _12749_, _06150_);
  nor (_26039_, _26038_, _06316_);
  nand (_26040_, _26039_, _26037_);
  and (_26041_, _06316_, _05853_);
  nor (_26042_, _26041_, _25353_);
  and (_26043_, _26042_, _26040_);
  nor (_26044_, _12756_, _06150_);
  or (_26045_, _26044_, _26043_);
  nand (_26046_, _26045_, _07059_);
  and (_26047_, _07458_, _06215_);
  nor (_26048_, _26047_, _05652_);
  nand (_26049_, _26048_, _26046_);
  and (_26050_, _26034_, _05652_);
  nor (_26051_, _26050_, _12772_);
  nand (_26052_, _26051_, _26049_);
  nor (_26055_, _12771_, _06150_);
  nor (_26056_, _26055_, _06047_);
  and (_26057_, _26056_, _26052_);
  or (_26058_, _26057_, _25734_);
  nand (_26059_, _26058_, _12779_);
  nor (_26060_, _12779_, _05870_);
  nor (_26061_, _26060_, _24749_);
  nand (_26062_, _26061_, _26059_);
  and (_26063_, _24749_, _06215_);
  nor (_26064_, _26063_, _12789_);
  and (_26065_, _26064_, _26062_);
  and (_26066_, _12789_, _06150_);
  or (_26067_, _26066_, _26065_);
  or (_26068_, _26067_, _01340_);
  or (_26069_, _01336_, \oc8051_golden_model_1.PC [3]);
  and (_26070_, _26069_, _42882_);
  and (_43420_, _26070_, _26068_);
  and (_26071_, _08581_, _07458_);
  nor (_26072_, _11921_, _08742_);
  nor (_26073_, _12344_, _11921_);
  not (_26075_, \oc8051_golden_model_1.PC [4]);
  nor (_26076_, _05331_, _26075_);
  and (_26077_, _05331_, _26075_);
  nor (_26078_, _26077_, _26076_);
  not (_26079_, _26078_);
  and (_26080_, _26079_, _12012_);
  or (_26081_, _12174_, _12074_);
  and (_26082_, _12102_, _12099_);
  nor (_26083_, _26082_, _12103_);
  not (_26084_, _26083_);
  nand (_26086_, _26084_, _12174_);
  nand (_26087_, _26086_, _26081_);
  nand (_26088_, _26087_, _06104_);
  and (_26089_, _11922_, _06039_);
  and (_26090_, _08581_, _06943_);
  not (_26091_, _12205_);
  and (_26092_, _11922_, _06938_);
  nor (_26093_, _26092_, _06530_);
  nor (_26094_, _07250_, _26075_);
  or (_26095_, _26094_, _06938_);
  and (_26097_, _26095_, _26093_);
  nor (_26098_, _26079_, _12214_);
  or (_26099_, _26098_, _06943_);
  nor (_26100_, _26099_, _26097_);
  nor (_26101_, _26100_, _26091_);
  not (_26102_, _26101_);
  nor (_26103_, _26102_, _26090_);
  nor (_26104_, _26079_, _12205_);
  nor (_26105_, _26104_, _08384_);
  not (_26106_, _26105_);
  nor (_26108_, _26106_, _26103_);
  and (_26109_, _11942_, _11939_);
  nor (_26110_, _26109_, _11943_);
  nand (_26111_, _26110_, _12199_);
  or (_26112_, _12199_, _11922_);
  and (_26113_, _26112_, _26111_);
  and (_26114_, _26113_, _08384_);
  or (_26115_, _26114_, _26108_);
  nand (_26116_, _26115_, _06949_);
  and (_26117_, _26079_, _06948_);
  nor (_26119_, _26117_, _06102_);
  nand (_26120_, _26119_, _26116_);
  or (_26121_, _12187_, _12074_);
  or (_26122_, _26083_, _12189_);
  and (_26123_, _26122_, _06102_);
  nand (_26124_, _26123_, _26121_);
  nand (_26125_, _26124_, _26120_);
  nand (_26126_, _26125_, _12182_);
  nor (_26127_, _26079_, _12182_);
  nor (_26128_, _26127_, _06043_);
  nand (_26129_, _26128_, _26126_);
  and (_26130_, _11922_, _06043_);
  nor (_26131_, _26130_, _07272_);
  nand (_26132_, _26131_, _26129_);
  nor (_26133_, _08581_, _05690_);
  nor (_26134_, _26133_, _06239_);
  nand (_26135_, _26134_, _26132_);
  and (_26136_, _11922_, _06239_);
  nor (_26137_, _26136_, _12232_);
  nand (_26138_, _26137_, _26135_);
  nor (_26140_, _26079_, _12231_);
  nor (_26141_, _26140_, _06219_);
  nand (_26142_, _26141_, _26138_);
  and (_26143_, _11922_, _06219_);
  nor (_26144_, _26143_, _12241_);
  nand (_26145_, _26144_, _26142_);
  nor (_26146_, _26079_, _12239_);
  nor (_26147_, _26146_, _06039_);
  and (_26148_, _26147_, _26145_);
  or (_26149_, _26148_, _26089_);
  nand (_26151_, _26149_, _05694_);
  and (_26152_, _08581_, _12243_);
  nor (_26153_, _26152_, _06038_);
  nand (_26154_, _26153_, _26151_);
  and (_26155_, _11921_, _06038_);
  nor (_26156_, _26155_, _12256_);
  and (_26157_, _26156_, _26154_);
  and (_26158_, _12289_, _12074_);
  nor (_26159_, _26084_, _12289_);
  or (_26160_, _26159_, _12255_);
  nor (_26162_, _26160_, _26158_);
  or (_26163_, _26162_, _26157_);
  nand (_26164_, _26163_, _12258_);
  nand (_26165_, _26164_, _26088_);
  nand (_26166_, _26165_, _06509_);
  nor (_26167_, _26084_, _12310_);
  not (_26168_, _26167_);
  and (_26169_, _12310_, _12074_);
  nor (_26170_, _26169_, _06509_);
  and (_26171_, _26170_, _26168_);
  nor (_26173_, _26171_, _06115_);
  nand (_26174_, _26173_, _26166_);
  nor (_26175_, _26083_, _12329_);
  and (_26176_, _12329_, _12075_);
  nor (_26177_, _26176_, _12298_);
  not (_26178_, _26177_);
  nor (_26179_, _26178_, _26175_);
  nor (_26180_, _26179_, _12012_);
  and (_26181_, _26180_, _26174_);
  or (_26182_, _26181_, _26080_);
  nand (_26184_, _26182_, _06033_);
  and (_26185_, _11922_, _06032_);
  nor (_26186_, _26185_, _07355_);
  nand (_26187_, _26186_, _26184_);
  nor (_26188_, _08581_, _05686_);
  nor (_26189_, _26188_, _25133_);
  and (_26190_, _26189_, _26187_);
  or (_26191_, _26190_, _26073_);
  nand (_26192_, _26191_, _12351_);
  nor (_26193_, _26078_, _12351_);
  nor (_26194_, _26193_, _06251_);
  nand (_26195_, _26194_, _26192_);
  and (_26196_, _11921_, _06251_);
  nor (_26197_, _26196_, _24866_);
  nand (_26198_, _26197_, _26195_);
  and (_26199_, _08581_, _24866_);
  nor (_26200_, _26199_, _06250_);
  and (_26201_, _26200_, _26198_);
  and (_26202_, _11921_, _06250_);
  or (_26203_, _26202_, _26201_);
  nand (_26205_, _26203_, _12362_);
  nor (_26206_, _26079_, _12362_);
  nor (_26207_, _26206_, _12367_);
  nand (_26208_, _26207_, _26205_);
  nor (_26209_, _11921_, _12366_);
  nor (_26210_, _26209_, _05676_);
  nand (_26211_, _26210_, _26208_);
  nor (_26212_, _26079_, _05675_);
  nor (_26213_, _26212_, _06026_);
  and (_26214_, _26213_, _26211_);
  and (_26216_, _11922_, _06026_);
  or (_26217_, _26216_, _26214_);
  nand (_26218_, _26217_, _05673_);
  and (_26219_, _08581_, _06023_);
  nor (_26220_, _26219_, _06110_);
  nand (_26221_, _26220_, _26218_);
  and (_26222_, _12074_, _06110_);
  nor (_26223_, _26222_, _09818_);
  nand (_26224_, _26223_, _26221_);
  nor (_26225_, _11921_, _09817_);
  nor (_26227_, _26225_, _09833_);
  nand (_26228_, _26227_, _26224_);
  nor (_26229_, _12075_, _05669_);
  nor (_26230_, _26229_, _12393_);
  nand (_26231_, _26230_, _26228_);
  nor (_26232_, _26078_, _12389_);
  nor (_26233_, _26232_, _06089_);
  nand (_26234_, _26233_, _26231_);
  and (_26235_, _11921_, _06089_);
  nor (_26236_, _26235_, _05719_);
  nand (_26238_, _26236_, _26234_);
  and (_26239_, _08581_, _05719_);
  nor (_26240_, _26239_, _12397_);
  nand (_26241_, _26240_, _26238_);
  and (_26242_, _26110_, _12397_);
  nor (_26243_, _26242_, _08743_);
  and (_26244_, _26243_, _26241_);
  or (_26245_, _26244_, _26072_);
  nand (_26246_, _26245_, _06020_);
  and (_26247_, _12075_, _06019_);
  nor (_26249_, _26247_, _10661_);
  and (_26250_, _26249_, _26246_);
  and (_26251_, _11921_, _10661_);
  or (_26252_, _26251_, _26250_);
  nand (_26253_, _26252_, _12413_);
  and (_26254_, _12431_, _12428_);
  nor (_26255_, _26254_, _12432_);
  and (_26256_, _26255_, _12412_);
  nor (_26257_, _26256_, _06088_);
  and (_26258_, _26257_, _26253_);
  and (_26259_, _11922_, _06088_);
  or (_26260_, _26259_, _26258_);
  nand (_26261_, _26260_, _13587_);
  and (_26262_, _08581_, _05724_);
  nor (_26263_, _26262_, _12453_);
  and (_26264_, _26263_, _26261_);
  and (_26265_, _11921_, _11071_);
  and (_26266_, _26110_, _12459_);
  or (_26267_, _26266_, _26265_);
  and (_26268_, _26267_, _12453_);
  or (_26270_, _26268_, _26264_);
  nand (_26271_, _26270_, _12007_);
  and (_26272_, _26078_, _12006_);
  nor (_26273_, _26272_, _12467_);
  nand (_26274_, _26273_, _26271_);
  nor (_26275_, _12466_, _11921_);
  nor (_26276_, _26275_, _06112_);
  nand (_26277_, _26276_, _26274_);
  and (_26278_, _12074_, _06112_);
  nor (_26279_, _26278_, _06284_);
  and (_26281_, _26279_, _26277_);
  and (_26282_, _11922_, _06284_);
  or (_26283_, _26282_, _26281_);
  nand (_26284_, _26283_, _24769_);
  and (_26285_, _08581_, _05727_);
  nor (_26286_, _26285_, _12476_);
  and (_26287_, _26286_, _26284_);
  nor (_26288_, _11922_, _11071_);
  and (_26289_, _26110_, _11071_);
  or (_26290_, _26289_, _26288_);
  and (_26292_, _26290_, _12476_);
  or (_26293_, _26292_, _26287_);
  nand (_26294_, _26293_, _12002_);
  nor (_26295_, _26079_, _12002_);
  nor (_26296_, _26295_, _10743_);
  nand (_26297_, _26296_, _26294_);
  nor (_26298_, _11921_, _10742_);
  nor (_26299_, _26298_, _06108_);
  nand (_26300_, _26299_, _26297_);
  and (_26301_, _12074_, _06108_);
  nor (_26303_, _26301_, _06277_);
  and (_26304_, _26303_, _26300_);
  and (_26305_, _11922_, _06277_);
  or (_26306_, _26305_, _26304_);
  nand (_26307_, _26306_, _24765_);
  and (_26308_, _08581_, _05736_);
  nor (_26309_, _26308_, _12497_);
  and (_26310_, _26309_, _26307_);
  and (_26311_, _11921_, \oc8051_golden_model_1.PSW [7]);
  and (_26312_, _26110_, _10606_);
  or (_26314_, _26312_, _26311_);
  and (_26315_, _26314_, _12497_);
  or (_26316_, _26315_, _26310_);
  nand (_26317_, _26316_, _11993_);
  nor (_26318_, _26079_, _11993_);
  nor (_26319_, _26318_, _11987_);
  nand (_26320_, _26319_, _26317_);
  nor (_26321_, _11921_, _11986_);
  nor (_26322_, _26321_, _06130_);
  nand (_26323_, _26322_, _26320_);
  and (_26324_, _12074_, _06130_);
  nor (_26325_, _26324_, _06292_);
  and (_26326_, _26325_, _26323_);
  and (_26327_, _11922_, _06292_);
  or (_26328_, _26327_, _26326_);
  nand (_26329_, _26328_, _24759_);
  and (_26330_, _08581_, _05740_);
  nor (_26331_, _26330_, _11982_);
  and (_26332_, _26331_, _26329_);
  and (_26333_, _11921_, _10606_);
  and (_26335_, _26110_, \oc8051_golden_model_1.PSW [7]);
  or (_26336_, _26335_, _26333_);
  and (_26337_, _26336_, _11982_);
  or (_26338_, _26337_, _26332_);
  nand (_26339_, _26338_, _12523_);
  nor (_26340_, _26079_, _12523_);
  nor (_26341_, _26340_, _10826_);
  nand (_26342_, _26341_, _26339_);
  nor (_26343_, _11921_, _10825_);
  nor (_26344_, _26343_, _10854_);
  nand (_26346_, _26344_, _26342_);
  and (_26347_, _26078_, _10854_);
  nor (_26348_, _26347_, _06298_);
  and (_26349_, _26348_, _26346_);
  and (_26350_, _08937_, _06298_);
  or (_26351_, _26350_, _26349_);
  nand (_26352_, _26351_, _05734_);
  and (_26353_, _08581_, _05732_);
  nor (_26354_, _26353_, _06129_);
  and (_26355_, _26354_, _26352_);
  nor (_26357_, _12075_, _12722_);
  and (_26358_, _26083_, _12722_);
  nor (_26359_, _26358_, _26357_);
  nor (_26360_, _26359_, _06306_);
  or (_26361_, _26360_, _26355_);
  nand (_26362_, _26361_, _11872_);
  nor (_26363_, _26079_, _11872_);
  nor (_26364_, _26363_, _10976_);
  nand (_26365_, _26364_, _26362_);
  nor (_26366_, _11921_, _10975_);
  nor (_26368_, _26366_, _11015_);
  nand (_26369_, _26368_, _26365_);
  and (_26370_, _26078_, _11015_);
  nor (_26371_, _26370_, _06049_);
  nand (_26372_, _26371_, _26369_);
  and (_26373_, _08937_, _06049_);
  nor (_26374_, _26373_, _05747_);
  nand (_26375_, _26374_, _26372_);
  nor (_26376_, _08581_, _05748_);
  nor (_26377_, _26376_, _06126_);
  nand (_26379_, _26377_, _26375_);
  nor (_26380_, _26083_, _12722_);
  and (_26381_, _12075_, _12722_);
  nor (_26382_, _26381_, _26380_);
  nor (_26383_, _26382_, _06704_);
  nor (_26384_, _26383_, _12750_);
  nand (_26385_, _26384_, _26379_);
  nor (_26386_, _26079_, _12749_);
  nor (_26387_, _26386_, _06316_);
  nand (_26388_, _26387_, _26385_);
  and (_26390_, _11922_, _06316_);
  nor (_26391_, _26390_, _25353_);
  nand (_26392_, _26391_, _26388_);
  nor (_26393_, _26079_, _12756_);
  nor (_26394_, _26393_, _07458_);
  and (_26395_, _26394_, _26392_);
  or (_26396_, _26395_, _26071_);
  nand (_26397_, _26396_, _05653_);
  nor (_26398_, _26382_, _05653_);
  nor (_26399_, _26398_, _12772_);
  nand (_26401_, _26399_, _26397_);
  nor (_26402_, _26079_, _12771_);
  nor (_26403_, _26402_, _06047_);
  nand (_26404_, _26403_, _26401_);
  not (_26405_, _12779_);
  and (_26406_, _11922_, _06047_);
  nor (_26407_, _26406_, _26405_);
  nand (_26408_, _26407_, _26404_);
  nor (_26409_, _26079_, _12779_);
  nor (_26410_, _26409_, _24749_);
  nand (_26411_, _26410_, _26408_);
  and (_26412_, _24749_, _08581_);
  nor (_26413_, _26412_, _12789_);
  and (_26414_, _26413_, _26411_);
  and (_26415_, _26078_, _12789_);
  or (_26416_, _26415_, _26414_);
  or (_26417_, _26416_, _01340_);
  or (_26418_, _01336_, \oc8051_golden_model_1.PC [4]);
  and (_26419_, _26418_, _42882_);
  and (_43421_, _26419_, _26417_);
  nor (_26421_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_26422_, _11916_, _05346_);
  nor (_26423_, _26422_, _26421_);
  and (_26424_, _26423_, _12789_);
  and (_26425_, _11916_, _06047_);
  nor (_26426_, _26423_, _11872_);
  nor (_26427_, _26423_, _12523_);
  nor (_26428_, _26423_, _11993_);
  nor (_26429_, _26423_, _12002_);
  not (_26430_, _26423_);
  and (_26432_, _26430_, _12006_);
  nor (_26433_, _11916_, _08742_);
  and (_26434_, _26430_, _12012_);
  and (_26435_, _12172_, _12069_);
  or (_26436_, _12071_, _12072_);
  and (_26437_, _26436_, _12104_);
  nor (_26438_, _26436_, _12104_);
  nor (_26439_, _26438_, _26437_);
  and (_26440_, _26439_, _12174_);
  nor (_26441_, _26440_, _26435_);
  nand (_26443_, _26441_, _06104_);
  nor (_26444_, _08612_, _07233_);
  nand (_26445_, _11917_, _06938_);
  and (_26446_, _26445_, _25758_);
  and (_26447_, _07251_, \oc8051_golden_model_1.PC [5]);
  or (_26448_, _26447_, _06938_);
  and (_26449_, _26448_, _26446_);
  or (_26450_, _26430_, _12214_);
  nand (_26451_, _26450_, _12205_);
  or (_26452_, _26451_, _26449_);
  and (_26454_, _26452_, _07233_);
  or (_26455_, _26454_, _26444_);
  or (_26456_, _26423_, _12205_);
  and (_26457_, _26456_, _26455_);
  nor (_26458_, _26457_, _08384_);
  or (_26459_, _11919_, _11918_);
  and (_26460_, _26459_, _11944_);
  nor (_26461_, _26459_, _11944_);
  or (_26462_, _26461_, _26460_);
  or (_26463_, _26462_, _12197_);
  or (_26465_, _12199_, _11917_);
  and (_26466_, _26465_, _08384_);
  and (_26467_, _26466_, _26463_);
  or (_26468_, _26467_, _26458_);
  nand (_26469_, _26468_, _06949_);
  and (_26470_, _26430_, _06948_);
  nor (_26471_, _26470_, _06102_);
  nand (_26472_, _26471_, _26469_);
  or (_26473_, _12187_, _12069_);
  or (_26474_, _26439_, _12189_);
  and (_26475_, _26474_, _06102_);
  nand (_26476_, _26475_, _26473_);
  and (_26477_, _26476_, _12182_);
  nand (_26478_, _26477_, _26472_);
  nor (_26479_, _26423_, _12182_);
  nor (_26480_, _26479_, _06043_);
  nand (_26481_, _26480_, _26478_);
  and (_26482_, _11916_, _06043_);
  nor (_26483_, _26482_, _07272_);
  nand (_26484_, _26483_, _26481_);
  and (_26486_, _08612_, _07272_);
  nor (_26487_, _26486_, _06239_);
  nand (_26488_, _26487_, _26484_);
  and (_26489_, _11916_, _06239_);
  nor (_26490_, _26489_, _12232_);
  nand (_26491_, _26490_, _26488_);
  nor (_26492_, _26423_, _12231_);
  nor (_26493_, _26492_, _06219_);
  nand (_26494_, _26493_, _26491_);
  and (_26495_, _11916_, _06219_);
  nor (_26497_, _26495_, _12241_);
  nand (_26498_, _26497_, _26494_);
  nor (_26499_, _26423_, _12239_);
  nor (_26500_, _26499_, _06039_);
  nand (_26501_, _26500_, _26498_);
  and (_26502_, _11916_, _06039_);
  nor (_26503_, _26502_, _12243_);
  nand (_26504_, _26503_, _26501_);
  and (_26505_, _08612_, _12243_);
  nor (_26506_, _26505_, _06038_);
  nand (_26508_, _26506_, _26504_);
  and (_26509_, _11916_, _06038_);
  nor (_26510_, _26509_, _12256_);
  and (_26511_, _26510_, _26508_);
  and (_26512_, _12289_, _12069_);
  not (_26513_, _26439_);
  nor (_26514_, _26513_, _12289_);
  or (_26515_, _26514_, _26512_);
  nor (_26516_, _26515_, _12255_);
  or (_26517_, _26516_, _26511_);
  nand (_26518_, _26517_, _12258_);
  nand (_26519_, _26518_, _26443_);
  nand (_26520_, _26519_, _06509_);
  nor (_26521_, _26513_, _12310_);
  not (_26522_, _26521_);
  and (_26523_, _12310_, _12069_);
  nor (_26524_, _26523_, _06509_);
  and (_26525_, _26524_, _26522_);
  nor (_26526_, _26525_, _06115_);
  nand (_26527_, _26526_, _26520_);
  nor (_26530_, _26439_, _12329_);
  and (_26531_, _12329_, _12070_);
  nor (_26532_, _26531_, _12298_);
  not (_26533_, _26532_);
  nor (_26534_, _26533_, _26530_);
  nor (_26535_, _26534_, _12012_);
  and (_26536_, _26535_, _26527_);
  or (_26537_, _26536_, _26434_);
  nand (_26538_, _26537_, _06033_);
  and (_26539_, _11917_, _06032_);
  nor (_26541_, _26539_, _07355_);
  nand (_26542_, _26541_, _26538_);
  nor (_26543_, _08612_, _05686_);
  nor (_26544_, _26543_, _25133_);
  and (_26545_, _26544_, _26542_);
  nor (_26546_, _12344_, _11916_);
  or (_26547_, _26546_, _26545_);
  nand (_26548_, _26547_, _12351_);
  nor (_26549_, _26423_, _12351_);
  nor (_26550_, _26549_, _06251_);
  nand (_26552_, _26550_, _26548_);
  and (_26553_, _11916_, _06251_);
  nor (_26554_, _26553_, _24866_);
  nand (_26555_, _26554_, _26552_);
  and (_26556_, _08612_, _24866_);
  nor (_26557_, _26556_, _06250_);
  nand (_26558_, _26557_, _26555_);
  and (_26559_, _11916_, _06250_);
  nor (_26560_, _26559_, _12368_);
  and (_26561_, _26560_, _26558_);
  nor (_26563_, _26423_, _12362_);
  or (_26564_, _26563_, _26561_);
  nand (_26565_, _26564_, _12366_);
  nor (_26566_, _11916_, _12366_);
  nor (_26567_, _26566_, _05676_);
  nand (_26568_, _26567_, _26565_);
  nor (_26569_, _26430_, _05675_);
  nor (_26570_, _26569_, _06026_);
  and (_26571_, _26570_, _26568_);
  and (_26572_, _11917_, _06026_);
  or (_26574_, _26572_, _26571_);
  nand (_26575_, _26574_, _05673_);
  and (_26576_, _08612_, _06023_);
  nor (_26577_, _26576_, _06110_);
  nand (_26578_, _26577_, _26575_);
  and (_26579_, _12069_, _06110_);
  nor (_26580_, _26579_, _09818_);
  nand (_26581_, _26580_, _26578_);
  nor (_26582_, _11916_, _09817_);
  nor (_26583_, _26582_, _09833_);
  nand (_26585_, _26583_, _26581_);
  nor (_26586_, _12070_, _05669_);
  nor (_26587_, _26586_, _12393_);
  nand (_26588_, _26587_, _26585_);
  nor (_26589_, _26423_, _12389_);
  nor (_26590_, _26589_, _06089_);
  nand (_26591_, _26590_, _26588_);
  and (_26592_, _11916_, _06089_);
  nor (_26593_, _26592_, _05719_);
  nand (_26594_, _26593_, _26591_);
  and (_26596_, _08612_, _05719_);
  nor (_26597_, _26596_, _12397_);
  nand (_26598_, _26597_, _26594_);
  nor (_26599_, _26462_, _12398_);
  nor (_26600_, _26599_, _08743_);
  and (_26601_, _26600_, _26598_);
  or (_26602_, _26601_, _26433_);
  nand (_26603_, _26602_, _06020_);
  and (_26604_, _12070_, _06019_);
  nor (_26605_, _26604_, _10661_);
  and (_26607_, _26605_, _26603_);
  and (_26608_, _11916_, _10661_);
  or (_26609_, _26608_, _26607_);
  nand (_26610_, _26609_, _12413_);
  and (_26611_, _12433_, _12426_);
  nor (_26612_, _26611_, _12434_);
  and (_26613_, _26612_, _12412_);
  nor (_26614_, _26613_, _06088_);
  and (_26615_, _26614_, _26610_);
  and (_26616_, _11917_, _06088_);
  or (_26618_, _26616_, _26615_);
  nand (_26619_, _26618_, _13587_);
  and (_26620_, _08612_, _05724_);
  nor (_26621_, _26620_, _12453_);
  nand (_26622_, _26621_, _26619_);
  and (_26623_, _11916_, _11071_);
  nor (_26624_, _26462_, _11071_);
  or (_26625_, _26624_, _26623_);
  and (_26626_, _26625_, _12453_);
  nor (_26627_, _26626_, _12006_);
  and (_26629_, _26627_, _26622_);
  or (_26630_, _26629_, _26432_);
  nand (_26631_, _26630_, _12466_);
  nor (_26632_, _12466_, _11916_);
  nor (_26633_, _26632_, _06112_);
  nand (_26634_, _26633_, _26631_);
  and (_26635_, _12069_, _06112_);
  nor (_26636_, _26635_, _06284_);
  and (_26637_, _26636_, _26634_);
  and (_26638_, _11917_, _06284_);
  or (_26640_, _26638_, _26637_);
  nand (_26641_, _26640_, _24769_);
  and (_26642_, _08612_, _05727_);
  nor (_26643_, _26642_, _12476_);
  nand (_26644_, _26643_, _26641_);
  and (_26645_, _26462_, _11071_);
  nor (_26646_, _11916_, _11071_);
  nor (_26647_, _26646_, _12477_);
  not (_26648_, _26647_);
  nor (_26649_, _26648_, _26645_);
  nor (_26651_, _26649_, _12481_);
  and (_26652_, _26651_, _26644_);
  or (_26653_, _26652_, _26429_);
  nand (_26654_, _26653_, _10742_);
  nor (_26655_, _11916_, _10742_);
  nor (_26656_, _26655_, _06108_);
  nand (_26657_, _26656_, _26654_);
  and (_26658_, _12069_, _06108_);
  nor (_26659_, _26658_, _06277_);
  and (_26660_, _26659_, _26657_);
  and (_26662_, _11917_, _06277_);
  or (_26663_, _26662_, _26660_);
  nand (_26664_, _26663_, _24765_);
  and (_26665_, _08612_, _05736_);
  nor (_26666_, _26665_, _12497_);
  nand (_26667_, _26666_, _26664_);
  and (_26668_, _11916_, \oc8051_golden_model_1.PSW [7]);
  nor (_26669_, _26462_, \oc8051_golden_model_1.PSW [7]);
  or (_26670_, _26669_, _26668_);
  and (_26671_, _26670_, _12497_);
  nor (_26673_, _26671_, _12502_);
  and (_26674_, _26673_, _26667_);
  or (_26675_, _26674_, _26428_);
  nand (_26676_, _26675_, _11986_);
  nor (_26677_, _11916_, _11986_);
  nor (_26678_, _26677_, _06130_);
  nand (_26679_, _26678_, _26676_);
  and (_26680_, _12069_, _06130_);
  nor (_26681_, _26680_, _06292_);
  and (_26682_, _26681_, _26679_);
  and (_26684_, _11917_, _06292_);
  or (_26685_, _26684_, _26682_);
  nand (_26686_, _26685_, _24759_);
  and (_26687_, _08612_, _05740_);
  nor (_26688_, _26687_, _11982_);
  nand (_26689_, _26688_, _26686_);
  nand (_26690_, _26462_, \oc8051_golden_model_1.PSW [7]);
  or (_26691_, _11916_, \oc8051_golden_model_1.PSW [7]);
  and (_26692_, _26691_, _11982_);
  and (_26693_, _26692_, _26690_);
  nor (_26695_, _26693_, _12525_);
  and (_26696_, _26695_, _26689_);
  or (_26697_, _26696_, _26427_);
  nand (_26698_, _26697_, _10825_);
  nor (_26699_, _11916_, _10825_);
  nor (_26700_, _26699_, _10854_);
  nand (_26701_, _26700_, _26698_);
  and (_26702_, _26423_, _10854_);
  nor (_26703_, _26702_, _06298_);
  and (_26704_, _26703_, _26701_);
  and (_26706_, _08888_, _06298_);
  or (_26707_, _26706_, _26704_);
  nand (_26708_, _26707_, _05734_);
  and (_26709_, _08612_, _05732_);
  nor (_26710_, _26709_, _06129_);
  nand (_26711_, _26710_, _26708_);
  and (_26712_, _26513_, _12722_);
  nor (_26713_, _12069_, _12722_);
  or (_26714_, _26713_, _06306_);
  or (_26715_, _26714_, _26712_);
  and (_26717_, _26715_, _11872_);
  and (_26718_, _26717_, _26711_);
  or (_26719_, _26718_, _26426_);
  nand (_26720_, _26719_, _10975_);
  nor (_26721_, _11916_, _10975_);
  nor (_26722_, _26721_, _11015_);
  nand (_26723_, _26722_, _26720_);
  and (_26724_, _26423_, _11015_);
  nor (_26725_, _26724_, _06049_);
  and (_26726_, _26725_, _26723_);
  and (_26728_, _08888_, _06049_);
  or (_26729_, _26728_, _26726_);
  nand (_26730_, _26729_, _05748_);
  and (_26731_, _08612_, _05747_);
  nor (_26732_, _26731_, _06126_);
  nand (_26733_, _26732_, _26730_);
  and (_26734_, _12070_, _12722_);
  nor (_26735_, _26439_, _12722_);
  nor (_26736_, _26735_, _26734_);
  and (_26737_, _26736_, _06126_);
  nor (_26739_, _26737_, _12750_);
  nand (_26740_, _26739_, _26733_);
  nor (_26741_, _26423_, _12749_);
  nor (_26742_, _26741_, _06316_);
  nand (_26743_, _26742_, _26740_);
  and (_26744_, _11916_, _06316_);
  nor (_26745_, _26744_, _25353_);
  and (_26746_, _26745_, _26743_);
  nor (_26747_, _26423_, _12756_);
  or (_26748_, _26747_, _26746_);
  nand (_26749_, _26748_, _07059_);
  and (_26750_, _08612_, _07458_);
  nor (_26751_, _26750_, _05652_);
  nand (_26752_, _26751_, _26749_);
  and (_26753_, _26736_, _05652_);
  nor (_26754_, _26753_, _12772_);
  nand (_26755_, _26754_, _26752_);
  nor (_26756_, _26423_, _12771_);
  nor (_26757_, _26756_, _06047_);
  and (_26758_, _26757_, _26755_);
  or (_26761_, _26758_, _26425_);
  nand (_26762_, _26761_, _12779_);
  nor (_26763_, _26430_, _12779_);
  nor (_26764_, _26763_, _24749_);
  nand (_26765_, _26764_, _26762_);
  and (_26766_, _24749_, _08612_);
  nor (_26767_, _26766_, _12789_);
  and (_26768_, _26767_, _26765_);
  or (_26769_, _26768_, _26424_);
  or (_26770_, _26769_, _01340_);
  or (_26772_, _01336_, \oc8051_golden_model_1.PC [5]);
  and (_26773_, _26772_, _42882_);
  and (_43422_, _26773_, _26770_);
  and (_26774_, _08647_, _07458_);
  and (_26775_, _08386_, _11860_);
  nor (_26776_, _26775_, \oc8051_golden_model_1.PC [6]);
  nor (_26777_, _26776_, _11861_);
  not (_26778_, _26777_);
  and (_26779_, _26778_, _11015_);
  and (_26780_, _12063_, _06130_);
  and (_26782_, _12063_, _06108_);
  and (_26783_, _12063_, _06112_);
  and (_26784_, _11909_, _06088_);
  nor (_26785_, _12344_, _11908_);
  and (_26786_, _26778_, _12012_);
  nor (_26787_, _12106_, _12066_);
  nor (_26788_, _26787_, _12107_);
  or (_26789_, _26788_, _12172_);
  or (_26790_, _12174_, _12062_);
  nand (_26791_, _26790_, _26789_);
  nand (_26793_, _26791_, _06104_);
  and (_26794_, _11909_, _06039_);
  or (_26795_, _26788_, _12189_);
  or (_26796_, _12187_, _12062_);
  and (_26797_, _26796_, _06102_);
  nand (_26798_, _26797_, _26795_);
  and (_26799_, _11946_, _11913_);
  nor (_26800_, _26799_, _11947_);
  nand (_26801_, _26800_, _12199_);
  or (_26802_, _12199_, _11909_);
  and (_26804_, _26802_, _08384_);
  nand (_26805_, _26804_, _26801_);
  not (_26806_, _12219_);
  and (_26807_, _08647_, _06943_);
  and (_26808_, _11909_, _06938_);
  nor (_26809_, _26808_, _06530_);
  and (_26810_, _07251_, \oc8051_golden_model_1.PC [6]);
  or (_26811_, _26810_, _06938_);
  and (_26812_, _26811_, _26809_);
  nor (_26813_, _26778_, _12214_);
  or (_26815_, _26813_, _06943_);
  nor (_26816_, _26815_, _26812_);
  nor (_26817_, _26816_, _26091_);
  not (_26818_, _26817_);
  nor (_26819_, _26818_, _26807_);
  nor (_26820_, _26778_, _12205_);
  nor (_26821_, _26820_, _08384_);
  not (_26822_, _26821_);
  nor (_26823_, _26822_, _26819_);
  nor (_26824_, _26823_, _26806_);
  nand (_26826_, _26824_, _26805_);
  nand (_26827_, _26826_, _26798_);
  nand (_26828_, _26827_, _12182_);
  nor (_26829_, _26778_, _12225_);
  nor (_26830_, _26829_, _06043_);
  nand (_26831_, _26830_, _26828_);
  and (_26832_, _11909_, _06043_);
  nor (_26833_, _26832_, _07272_);
  nand (_26834_, _26833_, _26831_);
  nor (_26835_, _08647_, _05690_);
  nor (_26837_, _26835_, _06239_);
  nand (_26838_, _26837_, _26834_);
  and (_26839_, _11909_, _06239_);
  nor (_26840_, _26839_, _12232_);
  nand (_26841_, _26840_, _26838_);
  nor (_26842_, _26778_, _12231_);
  nor (_26843_, _26842_, _06219_);
  nand (_26844_, _26843_, _26841_);
  and (_26845_, _11909_, _06219_);
  nor (_26846_, _26845_, _12241_);
  nand (_26848_, _26846_, _26844_);
  nor (_26849_, _26778_, _12239_);
  nor (_26850_, _26849_, _06039_);
  and (_26851_, _26850_, _26848_);
  or (_26852_, _26851_, _26794_);
  nand (_26853_, _26852_, _05694_);
  and (_26854_, _08647_, _12243_);
  nor (_26855_, _26854_, _06038_);
  nand (_26856_, _26855_, _26853_);
  and (_26857_, _11908_, _06038_);
  nor (_26859_, _26857_, _12256_);
  and (_26860_, _26859_, _26856_);
  and (_26861_, _12289_, _12062_);
  not (_26862_, _26861_);
  not (_26863_, _26788_);
  nor (_26864_, _26863_, _12289_);
  nor (_26865_, _26864_, _12255_);
  and (_26866_, _26865_, _26862_);
  or (_26867_, _26866_, _26860_);
  nand (_26868_, _26867_, _12258_);
  nand (_26870_, _26868_, _26793_);
  nand (_26871_, _26870_, _06509_);
  nor (_26872_, _26863_, _12310_);
  not (_26873_, _26872_);
  and (_26874_, _12310_, _12062_);
  nor (_26875_, _26874_, _06509_);
  and (_26876_, _26875_, _26873_);
  nor (_26877_, _26876_, _06115_);
  nand (_26878_, _26877_, _26871_);
  and (_26879_, _12329_, _12062_);
  not (_26881_, _12329_);
  and (_26882_, _26788_, _26881_);
  nor (_26883_, _26882_, _26879_);
  nor (_26884_, _26883_, _12298_);
  nor (_26885_, _26884_, _12012_);
  and (_26886_, _26885_, _26878_);
  or (_26887_, _26886_, _26786_);
  nand (_26888_, _26887_, _06033_);
  and (_26889_, _11909_, _06032_);
  nor (_26890_, _26889_, _07355_);
  nand (_26892_, _26890_, _26888_);
  nor (_26893_, _08647_, _05686_);
  nor (_26894_, _26893_, _25133_);
  and (_26895_, _26894_, _26892_);
  or (_26896_, _26895_, _26785_);
  nand (_26897_, _26896_, _12351_);
  nor (_26898_, _26777_, _12351_);
  nor (_26899_, _26898_, _06251_);
  nand (_26900_, _26899_, _26897_);
  and (_26901_, _11908_, _06251_);
  nor (_26903_, _26901_, _24866_);
  nand (_26904_, _26903_, _26900_);
  and (_26905_, _08647_, _24866_);
  nor (_26906_, _26905_, _06250_);
  nand (_26907_, _26906_, _26904_);
  and (_26908_, _11908_, _06250_);
  nor (_26909_, _26908_, _12368_);
  nand (_26910_, _26909_, _26907_);
  nor (_26911_, _26777_, _12362_);
  nor (_26912_, _26911_, _12367_);
  nand (_26914_, _26912_, _26910_);
  nor (_26915_, _11909_, _12366_);
  nor (_26916_, _26915_, _05676_);
  and (_26917_, _26916_, _26914_);
  nor (_26918_, _26777_, _05675_);
  or (_26919_, _26918_, _26917_);
  nand (_26920_, _26919_, _06027_);
  and (_26921_, _11909_, _06026_);
  nor (_26922_, _26921_, _06023_);
  nand (_26923_, _26922_, _26920_);
  nor (_26925_, _08647_, _05673_);
  nor (_26926_, _26925_, _06110_);
  nand (_26927_, _26926_, _26923_);
  and (_26928_, _12063_, _06110_);
  nor (_26929_, _26928_, _09818_);
  nand (_26930_, _26929_, _26927_);
  nor (_26931_, _11909_, _09817_);
  nor (_26932_, _26931_, _09833_);
  nand (_26933_, _26932_, _26930_);
  nor (_26934_, _12062_, _05669_);
  nor (_26936_, _26934_, _12393_);
  nand (_26937_, _26936_, _26933_);
  nor (_26938_, _26778_, _12389_);
  nor (_26939_, _26938_, _06089_);
  nand (_26940_, _26939_, _26937_);
  and (_26941_, _11909_, _06089_);
  nor (_26942_, _26941_, _05719_);
  nand (_26943_, _26942_, _26940_);
  nor (_26944_, _08647_, _05720_);
  nor (_26945_, _26944_, _12397_);
  nand (_26947_, _26945_, _26943_);
  nor (_26948_, _26800_, _12398_);
  nor (_26949_, _26948_, _08743_);
  nand (_26950_, _26949_, _26947_);
  nor (_26951_, _11909_, _08742_);
  nor (_26952_, _26951_, _06019_);
  nand (_26953_, _26952_, _26950_);
  and (_26954_, _12063_, _06019_);
  nor (_26955_, _26954_, _10661_);
  nand (_26956_, _26955_, _26953_);
  and (_26958_, _11908_, _10661_);
  nor (_26959_, _26958_, _12412_);
  and (_26960_, _26959_, _26956_);
  and (_26961_, _12435_, _12422_);
  nor (_26962_, _26961_, _12436_);
  nor (_26963_, _26962_, _12413_);
  or (_26964_, _26963_, _26960_);
  and (_26965_, _26964_, _06636_);
  or (_26966_, _26965_, _26784_);
  nand (_26967_, _26966_, _13587_);
  and (_26969_, _08647_, _05724_);
  nor (_26970_, _26969_, _12453_);
  nand (_26971_, _26970_, _26967_);
  and (_26972_, _11908_, _11071_);
  and (_26973_, _26800_, _12459_);
  or (_26974_, _26973_, _26972_);
  and (_26975_, _26974_, _12453_);
  nor (_26976_, _26975_, _12006_);
  nand (_26977_, _26976_, _26971_);
  and (_26978_, _26778_, _12006_);
  nor (_26980_, _26978_, _12467_);
  nand (_26981_, _26980_, _26977_);
  nor (_26982_, _12466_, _11909_);
  nor (_26983_, _26982_, _06112_);
  and (_26984_, _26983_, _26981_);
  or (_26985_, _26984_, _26783_);
  nand (_26986_, _26985_, _08756_);
  and (_26987_, _11909_, _06284_);
  nor (_26988_, _26987_, _05727_);
  and (_26989_, _26988_, _26986_);
  nor (_26991_, _08647_, _24769_);
  or (_26992_, _26991_, _26989_);
  nand (_26993_, _26992_, _12477_);
  nor (_26994_, _11909_, _11071_);
  and (_26995_, _26800_, _11071_);
  or (_26996_, _26995_, _26994_);
  and (_26997_, _26996_, _12476_);
  nor (_26998_, _26997_, _12481_);
  nand (_26999_, _26998_, _26993_);
  nor (_27000_, _26777_, _12002_);
  nor (_27002_, _27000_, _10743_);
  nand (_27003_, _27002_, _26999_);
  nor (_27004_, _11909_, _10742_);
  nor (_27005_, _27004_, _06108_);
  and (_27006_, _27005_, _27003_);
  or (_27007_, _27006_, _26782_);
  nand (_27008_, _27007_, _06278_);
  and (_27009_, _11909_, _06277_);
  nor (_27010_, _27009_, _05736_);
  and (_27011_, _27010_, _27008_);
  nor (_27013_, _08647_, _24765_);
  or (_27014_, _27013_, _27011_);
  nand (_27015_, _27014_, _12498_);
  and (_27016_, _11908_, \oc8051_golden_model_1.PSW [7]);
  and (_27017_, _26800_, _10606_);
  or (_27018_, _27017_, _27016_);
  and (_27019_, _27018_, _12497_);
  nor (_27020_, _27019_, _12502_);
  nand (_27021_, _27020_, _27015_);
  nor (_27022_, _26777_, _11993_);
  nor (_27024_, _27022_, _11987_);
  nand (_27025_, _27024_, _27021_);
  nor (_27026_, _11909_, _11986_);
  nor (_27027_, _27026_, _06130_);
  and (_27028_, _27027_, _27025_);
  or (_27029_, _27028_, _26780_);
  nand (_27030_, _27029_, _08782_);
  and (_27031_, _11909_, _06292_);
  nor (_27032_, _27031_, _05740_);
  and (_27033_, _27032_, _27030_);
  nor (_27035_, _08647_, _24759_);
  or (_27036_, _27035_, _27033_);
  nand (_27037_, _27036_, _12518_);
  or (_27038_, _26800_, _10606_);
  or (_27039_, _11908_, \oc8051_golden_model_1.PSW [7]);
  and (_27040_, _27039_, _11982_);
  and (_27041_, _27040_, _27038_);
  nor (_27042_, _27041_, _12525_);
  nand (_27043_, _27042_, _27037_);
  nor (_27044_, _26777_, _12523_);
  nor (_27046_, _27044_, _10826_);
  nand (_27047_, _27046_, _27043_);
  nor (_27048_, _11909_, _10825_);
  nor (_27049_, _27048_, _10854_);
  nand (_27050_, _27049_, _27047_);
  and (_27051_, _26778_, _10854_);
  nor (_27052_, _27051_, _06298_);
  nand (_27053_, _27052_, _27050_);
  and (_27054_, _09178_, _06298_);
  nor (_27055_, _27054_, _05732_);
  nand (_27057_, _27055_, _27053_);
  and (_27058_, _08647_, _05732_);
  nor (_27059_, _27058_, _06129_);
  nand (_27060_, _27059_, _27057_);
  and (_27061_, _26863_, _12722_);
  nor (_27062_, _12062_, _12722_);
  or (_27063_, _27062_, _06306_);
  nor (_27064_, _27063_, _27061_);
  nor (_27065_, _27064_, _12541_);
  nand (_27066_, _27065_, _27060_);
  nor (_27068_, _26777_, _11872_);
  nor (_27069_, _27068_, _10976_);
  nand (_27070_, _27069_, _27066_);
  nor (_27071_, _11909_, _10975_);
  nor (_27072_, _27071_, _11015_);
  and (_27073_, _27072_, _27070_);
  or (_27074_, _27073_, _26779_);
  nand (_27075_, _27074_, _06050_);
  and (_27076_, _08843_, _06049_);
  nor (_27077_, _27076_, _05747_);
  nand (_27079_, _27077_, _27075_);
  nor (_27080_, _08647_, _05748_);
  nor (_27081_, _27080_, _06126_);
  and (_27082_, _27081_, _27079_);
  nor (_27083_, _26788_, _12722_);
  and (_27084_, _12063_, _12722_);
  nor (_27085_, _27084_, _27083_);
  nor (_27086_, _27085_, _06704_);
  or (_27087_, _27086_, _27082_);
  and (_27088_, _27087_, _12749_);
  nor (_27090_, _26777_, _12749_);
  or (_27091_, _27090_, _27088_);
  nand (_27092_, _27091_, _06718_);
  and (_27093_, _11909_, _06316_);
  nor (_27094_, _27093_, _25353_);
  nand (_27095_, _27094_, _27092_);
  nor (_27096_, _26778_, _12756_);
  nor (_27097_, _27096_, _07458_);
  and (_27098_, _27097_, _27095_);
  or (_27099_, _27098_, _26774_);
  nand (_27101_, _27099_, _05653_);
  nor (_27102_, _27085_, _05653_);
  nor (_27103_, _27102_, _12772_);
  nand (_27104_, _27103_, _27101_);
  nor (_27105_, _26778_, _12771_);
  nor (_27106_, _27105_, _06047_);
  nand (_27107_, _27106_, _27104_);
  and (_27108_, _11909_, _06047_);
  nor (_27109_, _27108_, _26405_);
  nand (_27110_, _27109_, _27107_);
  nor (_27112_, _26778_, _12779_);
  nor (_27113_, _27112_, _24749_);
  nand (_27114_, _27113_, _27110_);
  and (_27115_, _24749_, _08647_);
  nor (_27116_, _27115_, _12789_);
  and (_27117_, _27116_, _27114_);
  and (_27118_, _26777_, _12789_);
  or (_27119_, _27118_, _27117_);
  or (_27120_, _27119_, _01340_);
  or (_27121_, _01336_, \oc8051_golden_model_1.PC [6]);
  and (_27123_, _27121_, _42882_);
  and (_43423_, _27123_, _27120_);
  and (_27124_, _08391_, _06047_);
  and (_27125_, _08391_, _06316_);
  nor (_27126_, _11861_, \oc8051_golden_model_1.PC [7]);
  nor (_27127_, _27126_, _11862_);
  nor (_27128_, _27127_, _11872_);
  nor (_27129_, _27127_, _12523_);
  nor (_27130_, _27127_, _11993_);
  nor (_27131_, _27127_, _12002_);
  not (_27133_, _27127_);
  and (_27134_, _27133_, _12006_);
  nor (_27135_, _08742_, _08391_);
  nor (_27136_, _12344_, _08391_);
  and (_27137_, _27133_, _12012_);
  nor (_27138_, _08332_, _07233_);
  nand (_27139_, _08524_, _06938_);
  and (_27140_, _27139_, _25758_);
  and (_27141_, _07251_, \oc8051_golden_model_1.PC [7]);
  or (_27142_, _27141_, _06938_);
  and (_27144_, _27142_, _27140_);
  or (_27145_, _27133_, _12214_);
  nand (_27146_, _27145_, _12205_);
  or (_27147_, _27146_, _27144_);
  and (_27148_, _27147_, _07233_);
  or (_27149_, _27148_, _27138_);
  or (_27150_, _27127_, _12205_);
  and (_27151_, _27150_, _27149_);
  nor (_27152_, _27151_, _08384_);
  or (_27153_, _11904_, _11905_);
  and (_27155_, _27153_, _11948_);
  nor (_27156_, _27153_, _11948_);
  nor (_27157_, _27156_, _27155_);
  nand (_27158_, _27157_, _12199_);
  or (_27159_, _12199_, _08524_);
  and (_27160_, _27159_, _08384_);
  and (_27161_, _27160_, _27158_);
  or (_27162_, _27161_, _27152_);
  nand (_27163_, _27162_, _06949_);
  and (_27164_, _27133_, _06948_);
  nor (_27166_, _27164_, _06102_);
  nand (_27167_, _27166_, _27163_);
  or (_27168_, _12187_, _09141_);
  and (_27169_, _12108_, _12059_);
  nor (_27170_, _27169_, _12109_);
  or (_27171_, _27170_, _12189_);
  and (_27172_, _27171_, _06102_);
  nand (_27173_, _27172_, _27168_);
  and (_27174_, _27173_, _12182_);
  nand (_27175_, _27174_, _27167_);
  nor (_27177_, _27127_, _12182_);
  nor (_27178_, _27177_, _06043_);
  nand (_27179_, _27178_, _27175_);
  and (_27180_, _08391_, _06043_);
  nor (_27181_, _27180_, _07272_);
  nand (_27182_, _27181_, _27179_);
  and (_27183_, _08332_, _07272_);
  nor (_27184_, _27183_, _06239_);
  nand (_27185_, _27184_, _27182_);
  and (_27186_, _08391_, _06239_);
  nor (_27188_, _27186_, _12232_);
  nand (_27189_, _27188_, _27185_);
  nor (_27190_, _27127_, _12231_);
  nor (_27191_, _27190_, _06219_);
  nand (_27192_, _27191_, _27189_);
  and (_27193_, _08391_, _06219_);
  nor (_27194_, _27193_, _12241_);
  nand (_27195_, _27194_, _27192_);
  nor (_27196_, _27127_, _12239_);
  nor (_27197_, _27196_, _06039_);
  nand (_27199_, _27197_, _27195_);
  and (_27200_, _08391_, _06039_);
  nor (_27201_, _27200_, _12243_);
  nand (_27202_, _27201_, _27199_);
  and (_27203_, _08332_, _12243_);
  nor (_27204_, _27203_, _06038_);
  nand (_27205_, _27204_, _27202_);
  and (_27206_, _08391_, _06038_);
  nor (_27207_, _27206_, _12256_);
  nand (_27208_, _27207_, _27205_);
  not (_27210_, _27170_);
  nor (_27211_, _27210_, _12289_);
  not (_27212_, _27211_);
  and (_27213_, _12289_, _09141_);
  nor (_27214_, _27213_, _12255_);
  and (_27215_, _27214_, _27212_);
  nor (_27216_, _27215_, _06104_);
  nand (_27217_, _27216_, _27208_);
  or (_27218_, _12174_, _09141_);
  or (_27219_, _27170_, _12172_);
  and (_27221_, _27219_, _06104_);
  nand (_27222_, _27221_, _27218_);
  and (_27223_, _27222_, _06509_);
  nand (_27224_, _27223_, _27217_);
  nor (_27225_, _27210_, _12310_);
  not (_27226_, _27225_);
  and (_27227_, _12310_, _09141_);
  nor (_27228_, _27227_, _06509_);
  and (_27229_, _27228_, _27226_);
  nor (_27230_, _27229_, _06115_);
  nand (_27232_, _27230_, _27224_);
  nor (_27233_, _27170_, _12329_);
  and (_27234_, _12329_, _09142_);
  nor (_27235_, _27234_, _12298_);
  not (_27236_, _27235_);
  nor (_27237_, _27236_, _27233_);
  nor (_27238_, _27237_, _12012_);
  and (_27239_, _27238_, _27232_);
  or (_27240_, _27239_, _27137_);
  nand (_27241_, _27240_, _06033_);
  and (_27243_, _08524_, _06032_);
  nor (_27244_, _27243_, _07355_);
  nand (_27245_, _27244_, _27241_);
  nor (_27246_, _08332_, _05686_);
  nor (_27247_, _27246_, _25133_);
  and (_27248_, _27247_, _27245_);
  or (_27249_, _27248_, _27136_);
  nand (_27250_, _27249_, _12351_);
  nor (_27251_, _27127_, _12351_);
  nor (_27252_, _27251_, _06251_);
  nand (_27254_, _27252_, _27250_);
  and (_27255_, _08391_, _06251_);
  nor (_27256_, _27255_, _24866_);
  nand (_27257_, _27256_, _27254_);
  and (_27258_, _08332_, _24866_);
  nor (_27259_, _27258_, _06250_);
  nand (_27260_, _27259_, _27257_);
  and (_27261_, _08391_, _06250_);
  nor (_27262_, _27261_, _12368_);
  and (_27263_, _27262_, _27260_);
  nor (_27265_, _27127_, _12362_);
  or (_27266_, _27265_, _27263_);
  nand (_27267_, _27266_, _12366_);
  nor (_27268_, _12366_, _08391_);
  nor (_27269_, _27268_, _05676_);
  nand (_27270_, _27269_, _27267_);
  nor (_27271_, _27133_, _05675_);
  nor (_27272_, _27271_, _06026_);
  and (_27273_, _27272_, _27270_);
  and (_27274_, _08524_, _06026_);
  or (_27276_, _27274_, _27273_);
  nand (_27277_, _27276_, _05673_);
  and (_27278_, _08332_, _06023_);
  nor (_27279_, _27278_, _06110_);
  nand (_27280_, _27279_, _27277_);
  and (_27281_, _09141_, _06110_);
  nor (_27282_, _27281_, _09818_);
  nand (_27283_, _27282_, _27280_);
  nor (_27284_, _09817_, _08391_);
  nor (_27285_, _27284_, _09833_);
  nand (_27287_, _27285_, _27283_);
  nor (_27288_, _09142_, _05669_);
  nor (_27289_, _27288_, _12393_);
  nand (_27290_, _27289_, _27287_);
  nor (_27291_, _27127_, _12389_);
  nor (_27292_, _27291_, _06089_);
  nand (_27293_, _27292_, _27290_);
  and (_27294_, _08391_, _06089_);
  nor (_27295_, _27294_, _05719_);
  nand (_27296_, _27295_, _27293_);
  and (_27298_, _08332_, _05719_);
  nor (_27299_, _27298_, _12397_);
  nand (_27300_, _27299_, _27296_);
  and (_27301_, _27157_, _12397_);
  nor (_27302_, _27301_, _08743_);
  and (_27303_, _27302_, _27300_);
  or (_27304_, _27303_, _27135_);
  nand (_27305_, _27304_, _06020_);
  and (_27306_, _09142_, _06019_);
  nor (_27307_, _27306_, _10661_);
  and (_27309_, _27307_, _27305_);
  and (_27310_, _10661_, _08391_);
  or (_27311_, _27310_, _27309_);
  nand (_27312_, _27311_, _12413_);
  or (_27313_, _12417_, _12418_);
  nor (_27314_, _27313_, _12437_);
  and (_27315_, _27313_, _12437_);
  nor (_27316_, _27315_, _27314_);
  and (_27317_, _27316_, _12412_);
  nor (_27318_, _27317_, _06088_);
  and (_27320_, _27318_, _27312_);
  and (_27321_, _08524_, _06088_);
  or (_27322_, _27321_, _27320_);
  nand (_27323_, _27322_, _13587_);
  and (_27324_, _08332_, _05724_);
  nor (_27325_, _27324_, _12453_);
  nand (_27326_, _27325_, _27323_);
  and (_27327_, _11071_, _08391_);
  and (_27328_, _27157_, _12459_);
  or (_27329_, _27328_, _27327_);
  and (_27330_, _27329_, _12453_);
  nor (_27331_, _27330_, _12006_);
  and (_27332_, _27331_, _27326_);
  or (_27333_, _27332_, _27134_);
  nand (_27334_, _27333_, _12466_);
  nor (_27335_, _12466_, _08391_);
  nor (_27336_, _27335_, _06112_);
  nand (_27337_, _27336_, _27334_);
  and (_27338_, _09141_, _06112_);
  nor (_27339_, _27338_, _06284_);
  and (_27342_, _27339_, _27337_);
  and (_27343_, _08524_, _06284_);
  or (_27344_, _27343_, _27342_);
  nand (_27345_, _27344_, _24769_);
  and (_27346_, _08332_, _05727_);
  nor (_27347_, _27346_, _12476_);
  nand (_27348_, _27347_, _27345_);
  nor (_27349_, _27157_, _12459_);
  nor (_27350_, _11071_, _08391_);
  nor (_27351_, _27350_, _12477_);
  not (_27353_, _27351_);
  nor (_27354_, _27353_, _27349_);
  nor (_27355_, _27354_, _12481_);
  and (_27356_, _27355_, _27348_);
  or (_27357_, _27356_, _27131_);
  nand (_27358_, _27357_, _10742_);
  nor (_27359_, _10742_, _08391_);
  nor (_27360_, _27359_, _06108_);
  nand (_27361_, _27360_, _27358_);
  and (_27362_, _09141_, _06108_);
  nor (_27364_, _27362_, _06277_);
  and (_27365_, _27364_, _27361_);
  and (_27366_, _08524_, _06277_);
  or (_27367_, _27366_, _27365_);
  nand (_27368_, _27367_, _24765_);
  and (_27369_, _08332_, _05736_);
  nor (_27370_, _27369_, _12497_);
  nand (_27371_, _27370_, _27368_);
  and (_27372_, _08391_, \oc8051_golden_model_1.PSW [7]);
  and (_27373_, _27157_, _10606_);
  or (_27375_, _27373_, _27372_);
  and (_27376_, _27375_, _12497_);
  nor (_27377_, _27376_, _12502_);
  and (_27378_, _27377_, _27371_);
  or (_27379_, _27378_, _27130_);
  nand (_27380_, _27379_, _11986_);
  nor (_27381_, _11986_, _08391_);
  nor (_27382_, _27381_, _06130_);
  nand (_27383_, _27382_, _27380_);
  and (_27384_, _09141_, _06130_);
  nor (_27386_, _27384_, _06292_);
  and (_27387_, _27386_, _27383_);
  and (_27388_, _08524_, _06292_);
  or (_27389_, _27388_, _27387_);
  nand (_27390_, _27389_, _24759_);
  and (_27391_, _08332_, _05740_);
  nor (_27392_, _27391_, _11982_);
  nand (_27393_, _27392_, _27390_);
  and (_27394_, _08391_, _10606_);
  and (_27395_, _27157_, \oc8051_golden_model_1.PSW [7]);
  or (_27397_, _27395_, _27394_);
  and (_27398_, _27397_, _11982_);
  nor (_27399_, _27398_, _12525_);
  and (_27400_, _27399_, _27393_);
  or (_27401_, _27400_, _27129_);
  nand (_27402_, _27401_, _10825_);
  nor (_27403_, _10825_, _08391_);
  nor (_27404_, _27403_, _10854_);
  nand (_27405_, _27404_, _27402_);
  and (_27406_, _27127_, _10854_);
  nor (_27408_, _27406_, _06298_);
  and (_27409_, _27408_, _27405_);
  and (_27410_, _08798_, _06298_);
  or (_27411_, _27410_, _27409_);
  nand (_27412_, _27411_, _05734_);
  and (_27413_, _08332_, _05732_);
  nor (_27414_, _27413_, _06129_);
  nand (_27415_, _27414_, _27412_);
  and (_27416_, _27210_, _12722_);
  nor (_27417_, _09141_, _12722_);
  or (_27419_, _27417_, _06306_);
  nor (_27420_, _27419_, _27416_);
  nor (_27421_, _27420_, _12541_);
  and (_27422_, _27421_, _27415_);
  or (_27423_, _27422_, _27128_);
  nand (_27424_, _27423_, _10975_);
  nor (_27425_, _10975_, _08391_);
  nor (_27426_, _27425_, _11015_);
  nand (_27427_, _27426_, _27424_);
  and (_27428_, _27127_, _11015_);
  nor (_27430_, _27428_, _06049_);
  and (_27431_, _27430_, _27427_);
  and (_27432_, _08798_, _06049_);
  or (_27433_, _27432_, _27431_);
  nand (_27434_, _27433_, _05748_);
  and (_27435_, _08332_, _05747_);
  nor (_27436_, _27435_, _06126_);
  nand (_27437_, _27436_, _27434_);
  and (_27438_, _09142_, _12722_);
  nor (_27439_, _27170_, _12722_);
  nor (_27441_, _27439_, _27438_);
  and (_27442_, _27441_, _06126_);
  nor (_27443_, _27442_, _12750_);
  nand (_27444_, _27443_, _27437_);
  nor (_27445_, _27127_, _12749_);
  nor (_27446_, _27445_, _06316_);
  and (_27447_, _27446_, _27444_);
  or (_27448_, _27447_, _27125_);
  nand (_27449_, _27448_, _12756_);
  nor (_27450_, _27133_, _12756_);
  nor (_27452_, _27450_, _07458_);
  nand (_27453_, _27452_, _27449_);
  and (_27454_, _08332_, _07458_);
  nor (_27455_, _27454_, _05652_);
  nand (_27456_, _27455_, _27453_);
  and (_27457_, _27441_, _05652_);
  nor (_27458_, _27457_, _12772_);
  nand (_27459_, _27458_, _27456_);
  nor (_27460_, _27127_, _12771_);
  nor (_27461_, _27460_, _06047_);
  and (_27463_, _27461_, _27459_);
  or (_27464_, _27463_, _27124_);
  nand (_27465_, _27464_, _12779_);
  nor (_27466_, _27133_, _12779_);
  nor (_27467_, _27466_, _24749_);
  nand (_27468_, _27467_, _27465_);
  and (_27469_, _24749_, _08332_);
  nor (_27470_, _27469_, _12789_);
  and (_27471_, _27470_, _27468_);
  and (_27472_, _27127_, _12789_);
  or (_27474_, _27472_, _27471_);
  or (_27475_, _27474_, _01340_);
  or (_27476_, _01336_, \oc8051_golden_model_1.PC [7]);
  and (_27477_, _27476_, _42882_);
  and (_43425_, _27477_, _27475_);
  and (_27478_, _11862_, \oc8051_golden_model_1.PC [8]);
  nor (_27479_, _11862_, \oc8051_golden_model_1.PC [8]);
  nor (_27480_, _27479_, _27478_);
  nor (_27481_, _27480_, _12779_);
  nor (_27482_, _09200_, _06016_);
  nor (_27484_, _11982_, _05740_);
  nor (_27485_, _11952_, _08742_);
  and (_27486_, _11952_, _06089_);
  or (_27487_, _27480_, _05675_);
  and (_27488_, _11952_, _06039_);
  nor (_27489_, _06239_, _07272_);
  and (_27490_, _11952_, _06043_);
  and (_27491_, _12205_, _07251_);
  or (_27492_, _27491_, _27480_);
  nand (_27493_, _14066_, _06938_);
  and (_27495_, _27493_, _25758_);
  or (_27496_, _06938_, \oc8051_golden_model_1.PC [8]);
  or (_27497_, _27496_, _07250_);
  nand (_27498_, _27497_, _27495_);
  nand (_27499_, _27498_, _24785_);
  and (_27500_, _27499_, _27492_);
  and (_27501_, _27480_, _06530_);
  or (_27502_, _27501_, _08384_);
  or (_27503_, _27502_, _27500_);
  nor (_27504_, _11955_, _11950_);
  nor (_27506_, _27504_, _11956_);
  and (_27507_, _27506_, _12199_);
  and (_27508_, _12197_, _11952_);
  or (_27509_, _27508_, _08383_);
  or (_27510_, _27509_, _27507_);
  and (_27511_, _27510_, _27503_);
  or (_27512_, _27511_, _06948_);
  not (_27513_, _27480_);
  nand (_27514_, _27513_, _06948_);
  and (_27515_, _27514_, _06954_);
  and (_27517_, _27515_, _27512_);
  and (_27518_, _12117_, _12110_);
  nor (_27519_, _27518_, _12118_);
  or (_27520_, _27519_, _12189_);
  or (_27521_, _12187_, _12112_);
  and (_27522_, _27521_, _06102_);
  and (_27523_, _27522_, _27520_);
  or (_27524_, _27523_, _24805_);
  or (_27525_, _27524_, _27517_);
  or (_27526_, _27480_, _12182_);
  and (_27528_, _27526_, _06044_);
  and (_27529_, _27528_, _27525_);
  or (_27530_, _27529_, _27490_);
  and (_27531_, _27530_, _27489_);
  nand (_27532_, _11952_, _06239_);
  nand (_27533_, _27532_, _12231_);
  or (_27534_, _27533_, _27531_);
  or (_27535_, _27480_, _12231_);
  and (_27536_, _27535_, _06220_);
  and (_27537_, _27536_, _27534_);
  nand (_27539_, _11952_, _06219_);
  nand (_27540_, _27539_, _12239_);
  or (_27541_, _27540_, _27537_);
  or (_27542_, _27480_, _12239_);
  and (_27543_, _27542_, _06040_);
  and (_27544_, _27543_, _27541_);
  or (_27545_, _27544_, _27488_);
  and (_27546_, _27545_, _12244_);
  nand (_27547_, _11952_, _06038_);
  nand (_27548_, _27547_, _12255_);
  or (_27550_, _27548_, _27546_);
  not (_27551_, _27519_);
  nor (_27552_, _27551_, _12289_);
  and (_27553_, _12289_, _12112_);
  or (_27554_, _27553_, _12255_);
  or (_27555_, _27554_, _27552_);
  and (_27556_, _27555_, _12258_);
  and (_27557_, _27556_, _27550_);
  and (_27558_, _27519_, _12174_);
  and (_27559_, _12172_, _12112_);
  or (_27561_, _27559_, _27558_);
  and (_27562_, _27561_, _06104_);
  or (_27563_, _27562_, _06121_);
  or (_27564_, _27563_, _27557_);
  nor (_27565_, _27551_, _12310_);
  and (_27566_, _12310_, _12112_);
  or (_27567_, _27566_, _06509_);
  or (_27568_, _27567_, _27565_);
  and (_27569_, _27568_, _12298_);
  and (_27570_, _27569_, _27564_);
  or (_27572_, _27519_, _12329_);
  nand (_27573_, _12329_, _12113_);
  and (_27574_, _27573_, _06115_);
  and (_27575_, _27574_, _27572_);
  or (_27576_, _27575_, _12012_);
  or (_27577_, _27576_, _27570_);
  nand (_27578_, _27513_, _12012_);
  and (_27579_, _27578_, _06033_);
  and (_27580_, _27579_, _27577_);
  and (_27581_, _11952_, _06032_);
  or (_27583_, _27581_, _07355_);
  or (_27584_, _27583_, _27580_);
  and (_27585_, _27584_, _12344_);
  nor (_27586_, _12344_, _14066_);
  or (_27587_, _27586_, _12355_);
  or (_27588_, _27587_, _27585_);
  or (_27589_, _27480_, _12351_);
  and (_27590_, _27589_, _13765_);
  and (_27591_, _27590_, _27588_);
  and (_27592_, _11952_, _06251_);
  or (_27594_, _27592_, _24866_);
  or (_27595_, _27594_, _27591_);
  and (_27596_, _27595_, _13764_);
  nand (_27597_, _11952_, _06250_);
  nand (_27598_, _27597_, _12362_);
  or (_27599_, _27598_, _27596_);
  or (_27600_, _27480_, _12362_);
  and (_27601_, _27600_, _12366_);
  and (_27602_, _27601_, _27599_);
  nor (_27603_, _14066_, _12366_);
  or (_27605_, _27603_, _05676_);
  or (_27606_, _27605_, _27602_);
  and (_27607_, _27606_, _27487_);
  or (_27608_, _27607_, _06026_);
  nand (_27609_, _14066_, _06026_);
  nor (_27610_, _06110_, _06023_);
  and (_27611_, _27610_, _27609_);
  and (_27612_, _27611_, _27608_);
  and (_27613_, _12112_, _06110_);
  or (_27614_, _27613_, _09818_);
  or (_27616_, _27614_, _27612_);
  nor (_27617_, _11952_, _09817_);
  nor (_27618_, _27617_, _09833_);
  nand (_27619_, _27618_, _27616_);
  nor (_27620_, _12113_, _05669_);
  nor (_27621_, _27620_, _12393_);
  nand (_27622_, _27621_, _27619_);
  nor (_27623_, _27480_, _12389_);
  nor (_27624_, _27623_, _06089_);
  and (_27625_, _27624_, _27622_);
  or (_27627_, _27625_, _27486_);
  nor (_27628_, _12397_, _05719_);
  nand (_27629_, _27628_, _27627_);
  and (_27630_, _27506_, _12397_);
  nor (_27631_, _27630_, _08743_);
  and (_27632_, _27631_, _27629_);
  or (_27633_, _27632_, _27485_);
  nand (_27634_, _27633_, _06020_);
  and (_27635_, _12113_, _06019_);
  nor (_27636_, _27635_, _10661_);
  nand (_27638_, _27636_, _27634_);
  and (_27639_, _11952_, _10661_);
  nor (_27640_, _27639_, _12412_);
  nand (_27641_, _27640_, _27638_);
  nor (_27642_, _12439_, \oc8051_golden_model_1.DPH [0]);
  nor (_27643_, _27642_, _12440_);
  nor (_27644_, _27643_, _12413_);
  nor (_27645_, _27644_, _06088_);
  nand (_27646_, _27645_, _27641_);
  and (_27647_, _11952_, _06088_);
  nor (_27649_, _27647_, _05724_);
  nand (_27650_, _27649_, _27646_);
  nand (_27651_, _27650_, _12454_);
  and (_27652_, _11952_, _11071_);
  and (_27653_, _27506_, _12459_);
  or (_27654_, _27653_, _27652_);
  and (_27655_, _27654_, _12453_);
  nor (_27656_, _27655_, _12006_);
  nand (_27657_, _27656_, _27651_);
  and (_27658_, _27513_, _12006_);
  nor (_27660_, _27658_, _12467_);
  nand (_27661_, _27660_, _27657_);
  nor (_27662_, _12466_, _14066_);
  nor (_27663_, _27662_, _06112_);
  nand (_27664_, _27663_, _27661_);
  and (_27665_, _12113_, _06112_);
  nor (_27666_, _27665_, _06284_);
  nand (_27667_, _27666_, _27664_);
  and (_27668_, _11952_, _06284_);
  nor (_27669_, _27668_, _05727_);
  nand (_27671_, _27669_, _27667_);
  nand (_27672_, _27671_, _12477_);
  nor (_27673_, _27506_, _12459_);
  nor (_27674_, _11952_, _11071_);
  nor (_27675_, _27674_, _12477_);
  not (_27676_, _27675_);
  nor (_27677_, _27676_, _27673_);
  nor (_27678_, _27677_, _12481_);
  nand (_27679_, _27678_, _27672_);
  nor (_27680_, _27480_, _12002_);
  nor (_27682_, _27680_, _10743_);
  nand (_27683_, _27682_, _27679_);
  nor (_27684_, _14066_, _10742_);
  nor (_27685_, _27684_, _06108_);
  and (_27686_, _27685_, _27683_);
  and (_27687_, _12113_, _06108_);
  or (_27688_, _27687_, _27686_);
  nand (_27689_, _27688_, _06278_);
  nor (_27690_, _12497_, _05736_);
  and (_27691_, _14066_, _06277_);
  not (_27693_, _27691_);
  and (_27694_, _27693_, _27690_);
  nand (_27695_, _27694_, _27689_);
  and (_27696_, _11952_, \oc8051_golden_model_1.PSW [7]);
  and (_27697_, _27506_, _10606_);
  or (_27698_, _27697_, _27696_);
  and (_27699_, _27698_, _12497_);
  nor (_27700_, _27699_, _12502_);
  nand (_27701_, _27700_, _27695_);
  nor (_27702_, _27480_, _11993_);
  nor (_27704_, _27702_, _11987_);
  and (_27705_, _27704_, _27701_);
  nor (_27706_, _14066_, _11986_);
  or (_27707_, _27706_, _06130_);
  or (_27708_, _27707_, _27705_);
  and (_27709_, _12113_, _06130_);
  nor (_27710_, _27709_, _06292_);
  and (_27711_, _27710_, _27708_);
  and (_27712_, _11952_, _06292_);
  or (_27713_, _27712_, _27711_);
  nand (_27715_, _27713_, _27484_);
  and (_27716_, _11952_, _10606_);
  and (_27717_, _27506_, \oc8051_golden_model_1.PSW [7]);
  or (_27718_, _27717_, _27716_);
  and (_27719_, _27718_, _11982_);
  nor (_27720_, _27719_, _12525_);
  nand (_27721_, _27720_, _27715_);
  nor (_27722_, _27480_, _12523_);
  nor (_27723_, _27722_, _10826_);
  and (_27724_, _27723_, _27721_);
  nor (_27726_, _14066_, _10825_);
  or (_27727_, _27726_, _10854_);
  or (_27728_, _27727_, _27724_);
  and (_27729_, _27513_, _10854_);
  nor (_27730_, _27729_, _06298_);
  nand (_27731_, _27730_, _27728_);
  and (_27732_, _06931_, _06298_);
  nor (_27733_, _27732_, _05732_);
  nand (_27734_, _27733_, _27731_);
  nand (_27735_, _27734_, _06306_);
  nor (_27737_, _12112_, _12722_);
  and (_27738_, _27551_, _12722_);
  or (_27739_, _27738_, _06306_);
  nor (_27740_, _27739_, _27737_);
  nor (_27741_, _27740_, _12541_);
  nand (_27742_, _27741_, _27735_);
  nor (_27743_, _27480_, _11872_);
  nor (_27744_, _27743_, _10976_);
  nand (_27745_, _27744_, _27742_);
  nor (_27746_, _14066_, _10975_);
  nor (_27748_, _27746_, _11015_);
  nand (_27749_, _27748_, _27745_);
  and (_27750_, _27513_, _11015_);
  nor (_27751_, _27750_, _06049_);
  nand (_27752_, _27751_, _27749_);
  and (_27753_, _06931_, _06049_);
  nor (_27754_, _27753_, _05747_);
  nand (_27755_, _27754_, _27752_);
  nand (_27756_, _27755_, _06704_);
  and (_27757_, _12113_, _12722_);
  nor (_27759_, _27519_, _12722_);
  nor (_27760_, _27759_, _27757_);
  and (_27761_, _27760_, _06126_);
  nor (_27762_, _27761_, _12750_);
  nand (_27763_, _27762_, _27756_);
  nor (_27764_, _27480_, _12749_);
  nor (_27765_, _27764_, _06316_);
  nand (_27766_, _27765_, _27763_);
  and (_27767_, _11952_, _06316_);
  nor (_27768_, _27767_, _25353_);
  nand (_27770_, _27768_, _27766_);
  nor (_27771_, _27480_, _12756_);
  nor (_27772_, _27771_, _06127_);
  and (_27773_, _27772_, _27770_);
  or (_27774_, _27773_, _27482_);
  nor (_27775_, _05752_, _05652_);
  nand (_27776_, _27775_, _27774_);
  and (_27777_, _27760_, _05652_);
  nor (_27778_, _27777_, _12772_);
  nand (_27779_, _27778_, _27776_);
  nor (_27781_, _27480_, _12771_);
  nor (_27782_, _27781_, _06047_);
  nand (_27783_, _27782_, _27779_);
  and (_27784_, _11952_, _06047_);
  nor (_27785_, _27784_, _26405_);
  and (_27786_, _27785_, _27783_);
  or (_27787_, _27786_, _27481_);
  nand (_27788_, _27787_, _12782_);
  nor (_27789_, _12789_, _05751_);
  not (_27790_, _27789_);
  and (_27792_, _06119_, _06016_);
  nor (_27793_, _27792_, _27790_);
  and (_27794_, _27793_, _27788_);
  and (_27795_, _27480_, _12789_);
  or (_27796_, _27795_, _27794_);
  or (_27797_, _27796_, _01340_);
  or (_27798_, _01336_, \oc8051_golden_model_1.PC [8]);
  and (_27799_, _27798_, _42882_);
  and (_43426_, _27799_, _27797_);
  nor (_27800_, _06799_, _09200_);
  nor (_27802_, _27478_, \oc8051_golden_model_1.PC [9]);
  nor (_27803_, _27802_, _11863_);
  nor (_27804_, _27803_, _11872_);
  nor (_27805_, _27803_, _12523_);
  and (_27806_, _12051_, _06130_);
  nor (_27807_, _27803_, _11993_);
  and (_27808_, _12051_, _06108_);
  nor (_27809_, _27803_, _12002_);
  and (_27810_, _12051_, _06112_);
  not (_27811_, _27803_);
  and (_27813_, _27811_, _12006_);
  nor (_27814_, _11900_, _08742_);
  and (_27815_, _11900_, _06089_);
  and (_27816_, _11900_, _06250_);
  nor (_27817_, _27803_, _12351_);
  or (_27818_, _12187_, _12051_);
  nor (_27819_, _12118_, _12114_);
  and (_27820_, _27819_, _12055_);
  nor (_27821_, _27819_, _12055_);
  nor (_27822_, _27821_, _27820_);
  not (_27824_, _27822_);
  or (_27825_, _27824_, _12189_);
  and (_27826_, _27825_, _27818_);
  or (_27827_, _27826_, _06954_);
  nor (_27828_, _11956_, _11953_);
  and (_27829_, _27828_, _11903_);
  nor (_27830_, _27828_, _11903_);
  nor (_27831_, _27830_, _27829_);
  or (_27832_, _27831_, _12197_);
  or (_27833_, _12199_, _14461_);
  and (_27835_, _27833_, _08384_);
  nand (_27836_, _27835_, _27832_);
  and (_27837_, _27803_, _06530_);
  or (_27838_, _27803_, _27491_);
  and (_27839_, _14461_, _06938_);
  nor (_27840_, _27839_, _06530_);
  or (_27841_, _06938_, \oc8051_golden_model_1.PC [9]);
  or (_27842_, _27841_, _07250_);
  nand (_27843_, _27842_, _27840_);
  nand (_27844_, _27843_, _24785_);
  and (_27846_, _27844_, _27838_);
  or (_27847_, _27846_, _08384_);
  nor (_27848_, _27847_, _27837_);
  nor (_27849_, _27848_, _06948_);
  and (_27850_, _27849_, _27836_);
  and (_27851_, _27803_, _06948_);
  or (_27852_, _27851_, _06102_);
  or (_27853_, _27852_, _27850_);
  nand (_27854_, _27853_, _27827_);
  nand (_27855_, _27854_, _12182_);
  nor (_27857_, _27803_, _12182_);
  nor (_27858_, _27857_, _06043_);
  nand (_27859_, _27858_, _27855_);
  and (_27860_, _11900_, _06043_);
  nor (_27861_, _27860_, _07272_);
  nand (_27862_, _27861_, _27859_);
  nand (_27863_, _27862_, _06848_);
  and (_27864_, _11900_, _06239_);
  nor (_27865_, _27864_, _12232_);
  nand (_27866_, _27865_, _27863_);
  nor (_27868_, _27803_, _12231_);
  nor (_27869_, _27868_, _06219_);
  nand (_27870_, _27869_, _27866_);
  and (_27871_, _11900_, _06219_);
  nor (_27872_, _27871_, _12241_);
  nand (_27873_, _27872_, _27870_);
  nor (_27874_, _27803_, _12239_);
  nor (_27875_, _27874_, _06039_);
  nand (_27876_, _27875_, _27873_);
  and (_27877_, _11900_, _06039_);
  nor (_27879_, _27877_, _12243_);
  nand (_27880_, _27879_, _27876_);
  nand (_27881_, _27880_, _07364_);
  and (_27882_, _11900_, _06038_);
  nor (_27883_, _27882_, _12256_);
  and (_27884_, _27883_, _27881_);
  and (_27885_, _12289_, _12051_);
  nor (_27886_, _27822_, _12289_);
  or (_27887_, _27886_, _27885_);
  nor (_27888_, _27887_, _12255_);
  or (_27890_, _27888_, _27884_);
  and (_27891_, _27890_, _13849_);
  and (_27892_, _12172_, _12051_);
  and (_27893_, _27824_, _12174_);
  or (_27894_, _27893_, _27892_);
  nor (_27895_, _27894_, _12258_);
  or (_27896_, _27895_, _27891_);
  or (_27897_, _27896_, _06121_);
  and (_27898_, _12310_, _12051_);
  nor (_27899_, _27822_, _12310_);
  nor (_27901_, _27899_, _27898_);
  or (_27902_, _27901_, _06509_);
  and (_27903_, _27902_, _27897_);
  or (_27904_, _27903_, _06115_);
  nand (_27905_, _12329_, _12051_);
  or (_27906_, _27822_, _12329_);
  and (_27907_, _27906_, _27905_);
  or (_27908_, _27907_, _12298_);
  and (_27909_, _27908_, _27904_);
  or (_27910_, _27909_, _12012_);
  nand (_27912_, _27803_, _12012_);
  and (_27913_, _27912_, _27910_);
  nand (_27914_, _27913_, _06033_);
  and (_27915_, _14461_, _06032_);
  not (_27916_, _27915_);
  and (_27917_, _12344_, _05686_);
  and (_27918_, _27917_, _27916_);
  nand (_27919_, _27918_, _27914_);
  nor (_27920_, _12344_, _14461_);
  nor (_27921_, _27920_, _12355_);
  and (_27923_, _27921_, _27919_);
  nor (_27924_, _27923_, _27817_);
  or (_27925_, _27924_, _06251_);
  nor (_27926_, _06250_, _24866_);
  nand (_27927_, _14461_, _06251_);
  and (_27928_, _27927_, _27926_);
  and (_27929_, _27928_, _27925_);
  or (_27930_, _27929_, _27816_);
  nand (_27931_, _27930_, _12362_);
  nor (_27932_, _27811_, _12362_);
  nor (_27934_, _27932_, _12367_);
  nand (_27935_, _27934_, _27931_);
  nor (_27936_, _11900_, _12366_);
  nor (_27937_, _27936_, _05676_);
  nand (_27938_, _27937_, _27935_);
  nor (_27939_, _27811_, _05675_);
  nor (_27940_, _27939_, _06026_);
  nand (_27941_, _27940_, _27938_);
  not (_27942_, _27610_);
  and (_27943_, _14461_, _06026_);
  nor (_27945_, _27943_, _27942_);
  nand (_27946_, _27945_, _27941_);
  and (_27947_, _12051_, _06110_);
  nor (_27948_, _27947_, _09818_);
  nand (_27949_, _27948_, _27946_);
  nor (_27950_, _11900_, _09817_);
  nor (_27951_, _27950_, _09833_);
  nand (_27952_, _27951_, _27949_);
  nor (_27953_, _12052_, _05669_);
  nor (_27954_, _27953_, _12393_);
  nand (_27956_, _27954_, _27952_);
  nor (_27957_, _27803_, _12389_);
  nor (_27958_, _27957_, _06089_);
  and (_27959_, _27958_, _27956_);
  or (_27960_, _27959_, _27815_);
  nand (_27961_, _27960_, _27628_);
  nor (_27962_, _27831_, _12398_);
  nor (_27963_, _27962_, _08743_);
  and (_27964_, _27963_, _27961_);
  or (_27965_, _27964_, _27814_);
  nand (_27966_, _27965_, _06020_);
  and (_27967_, _12052_, _06019_);
  nor (_27968_, _27967_, _10661_);
  nand (_27969_, _27968_, _27966_);
  and (_27970_, _11900_, _10661_);
  nor (_27971_, _27970_, _12412_);
  nand (_27972_, _27971_, _27969_);
  nor (_27973_, _12440_, \oc8051_golden_model_1.DPH [1]);
  nor (_27974_, _27973_, _12441_);
  nor (_27975_, _27974_, _12413_);
  nor (_27978_, _27975_, _06088_);
  nand (_27979_, _27978_, _27972_);
  and (_27980_, _11900_, _06088_);
  nor (_27981_, _27980_, _05724_);
  nand (_27982_, _27981_, _27979_);
  nand (_27983_, _27982_, _12454_);
  and (_27984_, _11900_, _11071_);
  nor (_27985_, _27831_, _11071_);
  or (_27986_, _27985_, _27984_);
  and (_27987_, _27986_, _12453_);
  nor (_27989_, _27987_, _12006_);
  and (_27990_, _27989_, _27983_);
  or (_27991_, _27990_, _27813_);
  nand (_27992_, _27991_, _12466_);
  nor (_27993_, _12466_, _11900_);
  nor (_27994_, _27993_, _06112_);
  and (_27995_, _27994_, _27992_);
  or (_27996_, _27995_, _27810_);
  nand (_27997_, _27996_, _08756_);
  and (_27998_, _11900_, _06284_);
  nor (_28000_, _27998_, _05727_);
  nand (_28001_, _28000_, _27997_);
  nand (_28002_, _28001_, _12477_);
  and (_28003_, _11900_, _12459_);
  nor (_28004_, _27831_, _12459_);
  or (_28005_, _28004_, _28003_);
  and (_28006_, _28005_, _12476_);
  nor (_28007_, _28006_, _12481_);
  and (_28008_, _28007_, _28002_);
  or (_28009_, _28008_, _27809_);
  nand (_28011_, _28009_, _10742_);
  nor (_28012_, _11900_, _10742_);
  nor (_28013_, _28012_, _06108_);
  and (_28014_, _28013_, _28011_);
  or (_28015_, _28014_, _27808_);
  nand (_28016_, _28015_, _06278_);
  and (_28017_, _11900_, _06277_);
  nor (_28018_, _28017_, _05736_);
  nand (_28019_, _28018_, _28016_);
  nand (_28020_, _28019_, _12498_);
  and (_28022_, _11900_, \oc8051_golden_model_1.PSW [7]);
  nor (_28023_, _27831_, \oc8051_golden_model_1.PSW [7]);
  or (_28024_, _28023_, _28022_);
  and (_28025_, _28024_, _12497_);
  nor (_28026_, _28025_, _12502_);
  and (_28027_, _28026_, _28020_);
  or (_28028_, _28027_, _27807_);
  nand (_28029_, _28028_, _11986_);
  nor (_28030_, _11900_, _11986_);
  nor (_28031_, _28030_, _06130_);
  and (_28033_, _28031_, _28029_);
  or (_28034_, _28033_, _27806_);
  nand (_28035_, _28034_, _08782_);
  and (_28036_, _11900_, _06292_);
  nor (_28037_, _28036_, _05740_);
  nand (_28038_, _28037_, _28035_);
  nand (_28039_, _28038_, _12518_);
  nand (_28040_, _27831_, \oc8051_golden_model_1.PSW [7]);
  or (_28041_, _11900_, \oc8051_golden_model_1.PSW [7]);
  and (_28042_, _28041_, _11982_);
  and (_28044_, _28042_, _28040_);
  nor (_28045_, _28044_, _12525_);
  and (_28046_, _28045_, _28039_);
  or (_28047_, _28046_, _27805_);
  nand (_28048_, _28047_, _10825_);
  nor (_28049_, _11900_, _10825_);
  nor (_28050_, _28049_, _10854_);
  nand (_28051_, _28050_, _28048_);
  and (_28052_, _27803_, _10854_);
  nor (_28053_, _28052_, _06298_);
  nand (_28055_, _28053_, _28051_);
  nor (_28056_, _06129_, _05732_);
  not (_28057_, _28056_);
  and (_28058_, _07132_, _06298_);
  nor (_28059_, _28058_, _28057_);
  nand (_28060_, _28059_, _28055_);
  nor (_28061_, _12051_, _12722_);
  and (_28062_, _27822_, _12722_);
  or (_28063_, _28062_, _06306_);
  nor (_28064_, _28063_, _28061_);
  nor (_28066_, _28064_, _12541_);
  and (_28067_, _28066_, _28060_);
  or (_28068_, _28067_, _27804_);
  nand (_28069_, _28068_, _10975_);
  nor (_28070_, _11900_, _10975_);
  nor (_28071_, _28070_, _11015_);
  nand (_28072_, _28071_, _28069_);
  and (_28073_, _27803_, _11015_);
  nor (_28074_, _28073_, _06049_);
  nand (_28075_, _28074_, _28072_);
  nor (_28077_, _06126_, _05747_);
  not (_28078_, _28077_);
  and (_28079_, _07132_, _06049_);
  nor (_28080_, _28079_, _28078_);
  nand (_28081_, _28080_, _28075_);
  and (_28082_, _12052_, _12722_);
  nor (_28083_, _27824_, _12722_);
  nor (_28084_, _28083_, _28082_);
  and (_28085_, _28084_, _06126_);
  nor (_28086_, _28085_, _12750_);
  nand (_28088_, _28086_, _28081_);
  nor (_28089_, _27803_, _12749_);
  nor (_28090_, _28089_, _06316_);
  nand (_28091_, _28090_, _28088_);
  and (_28092_, _11900_, _06316_);
  nor (_28093_, _28092_, _25353_);
  nand (_28094_, _28093_, _28091_);
  nor (_28095_, _27803_, _12756_);
  nor (_28096_, _28095_, _06127_);
  and (_28097_, _28096_, _28094_);
  or (_28099_, _28097_, _27800_);
  nand (_28100_, _28099_, _27775_);
  and (_28101_, _28084_, _05652_);
  nor (_28102_, _28101_, _12772_);
  nand (_28103_, _28102_, _28100_);
  nor (_28104_, _27803_, _12771_);
  nor (_28105_, _28104_, _06047_);
  nand (_28106_, _28105_, _28103_);
  and (_28107_, _11900_, _06047_);
  nor (_28108_, _28107_, _26405_);
  nand (_28110_, _28108_, _28106_);
  nor (_28111_, _27803_, _12779_);
  nor (_28112_, _28111_, _06119_);
  and (_28113_, _28112_, _28110_);
  nor (_28114_, _06799_, _12782_);
  or (_28115_, _28114_, _28113_);
  and (_28116_, _28115_, _27789_);
  and (_28117_, _27803_, _12789_);
  or (_28118_, _28117_, _28116_);
  or (_28119_, _28118_, _01340_);
  or (_28121_, _01336_, \oc8051_golden_model_1.PC [9]);
  and (_28122_, _28121_, _42882_);
  and (_43427_, _28122_, _28119_);
  nor (_28123_, _11863_, \oc8051_golden_model_1.PC [10]);
  nor (_28124_, _28123_, _11864_);
  and (_28125_, _28124_, _12393_);
  or (_28126_, _12344_, _11887_);
  or (_28127_, _28124_, _12231_);
  nor (_28128_, _12122_, _12119_);
  not (_28129_, _28128_);
  and (_28131_, _28129_, _12047_);
  nor (_28132_, _28129_, _12047_);
  nor (_28133_, _28132_, _28131_);
  and (_28134_, _28133_, _12187_);
  and (_28135_, _12189_, _12043_);
  or (_28136_, _28135_, _06954_);
  or (_28137_, _28136_, _28134_);
  nor (_28138_, _11960_, _11957_);
  not (_28139_, _28138_);
  and (_28140_, _28139_, _11896_);
  nor (_28142_, _28139_, _11896_);
  nor (_28143_, _28142_, _28140_);
  or (_28144_, _28143_, _12197_);
  or (_28145_, _12199_, _11887_);
  and (_28146_, _28145_, _28144_);
  or (_28147_, _28146_, _08383_);
  and (_28148_, _11887_, _06938_);
  nand (_28149_, _06939_, \oc8051_golden_model_1.PC [10]);
  nor (_28150_, _28149_, _07250_);
  or (_28151_, _28150_, _28148_);
  and (_28153_, _28151_, _25758_);
  or (_28154_, _28153_, _06943_);
  and (_28155_, _28154_, _12205_);
  not (_28156_, _12215_);
  and (_28157_, _28124_, _28156_);
  or (_28158_, _28157_, _08384_);
  or (_28159_, _28158_, _28155_);
  and (_28160_, _28159_, _06949_);
  and (_28161_, _28160_, _28147_);
  and (_28162_, _28124_, _06948_);
  or (_28164_, _28162_, _06102_);
  or (_28165_, _28164_, _28161_);
  and (_28166_, _28165_, _28137_);
  or (_28167_, _28166_, _24805_);
  or (_28168_, _28124_, _12182_);
  and (_28169_, _28168_, _06044_);
  and (_28170_, _28169_, _28167_);
  or (_28171_, _28170_, _07272_);
  and (_28172_, _28171_, _06848_);
  nor (_28173_, _14664_, _06244_);
  or (_28175_, _28173_, _12232_);
  or (_28176_, _28175_, _28172_);
  and (_28177_, _28176_, _28127_);
  or (_28178_, _28177_, _06219_);
  nand (_28179_, _14664_, _06219_);
  and (_28180_, _28179_, _12239_);
  and (_28181_, _28180_, _28178_);
  and (_28182_, _28124_, _12241_);
  or (_28183_, _28182_, _28181_);
  and (_28184_, _28183_, _06040_);
  and (_28186_, _11887_, _06039_);
  or (_28187_, _28186_, _12243_);
  or (_28188_, _28187_, _28184_);
  and (_28189_, _28188_, _07364_);
  nand (_28190_, _11887_, _06038_);
  nand (_28191_, _28190_, _12255_);
  or (_28192_, _28191_, _28189_);
  and (_28193_, _28133_, _13828_);
  and (_28194_, _12289_, _12043_);
  or (_28195_, _28194_, _12255_);
  or (_28197_, _28195_, _28193_);
  and (_28198_, _28197_, _28192_);
  or (_28199_, _28198_, _06104_);
  and (_28200_, _28133_, _12174_);
  and (_28201_, _12172_, _12043_);
  or (_28202_, _28201_, _12258_);
  or (_28203_, _28202_, _28200_);
  and (_28204_, _28203_, _28199_);
  or (_28205_, _28204_, _06121_);
  and (_28206_, _28133_, _12312_);
  and (_28208_, _12310_, _12043_);
  or (_28209_, _28208_, _06509_);
  or (_28210_, _28209_, _28206_);
  and (_28211_, _28210_, _12298_);
  and (_28212_, _28211_, _28205_);
  or (_28213_, _28133_, _12329_);
  nand (_28214_, _12329_, _12044_);
  and (_28215_, _28214_, _06115_);
  and (_28216_, _28215_, _28213_);
  or (_28217_, _28216_, _12012_);
  or (_28219_, _28217_, _28212_);
  or (_28220_, _28124_, _12013_);
  and (_28221_, _28220_, _06033_);
  and (_28222_, _28221_, _28219_);
  and (_28223_, _11887_, _06032_);
  nor (_28224_, _28223_, _28222_);
  nand (_28225_, _28224_, _27917_);
  and (_28226_, _28225_, _28126_);
  or (_28227_, _28226_, _12355_);
  or (_28228_, _28124_, _12351_);
  and (_28230_, _28228_, _13765_);
  and (_28231_, _28230_, _28227_);
  or (_28232_, _28231_, _24866_);
  and (_28233_, _28232_, _13764_);
  nor (_28234_, _14664_, _06252_);
  or (_28235_, _28234_, _12368_);
  or (_28236_, _28235_, _28233_);
  or (_28237_, _28124_, _12362_);
  and (_28238_, _28237_, _12366_);
  and (_28239_, _28238_, _28236_);
  nor (_28241_, _14664_, _12366_);
  or (_28242_, _28241_, _05676_);
  or (_28243_, _28242_, _28239_);
  or (_28244_, _28124_, _05675_);
  and (_28245_, _28244_, _06027_);
  and (_28246_, _28245_, _28243_);
  nand (_28247_, _11887_, _06026_);
  nand (_28248_, _28247_, _27610_);
  or (_28249_, _28248_, _28246_);
  nand (_28250_, _12044_, _06110_);
  and (_28252_, _28250_, _09817_);
  and (_28253_, _28252_, _28249_);
  nor (_28254_, _14664_, _09817_);
  or (_28255_, _28254_, _09833_);
  or (_28256_, _28255_, _28253_);
  or (_28257_, _12043_, _05669_);
  and (_28258_, _28257_, _12389_);
  and (_28259_, _28258_, _28256_);
  or (_28260_, _28259_, _28125_);
  and (_28261_, _28260_, _25023_);
  nand (_28263_, _11887_, _06089_);
  nand (_28264_, _28263_, _27628_);
  or (_28265_, _28264_, _28261_);
  or (_28266_, _28143_, _12398_);
  and (_28267_, _28266_, _08742_);
  and (_28268_, _28267_, _28265_);
  nor (_28269_, _14664_, _08742_);
  or (_28270_, _28269_, _06019_);
  or (_28271_, _28270_, _28268_);
  nand (_28272_, _12044_, _06019_);
  and (_28273_, _28272_, _10662_);
  and (_28274_, _28273_, _28271_);
  and (_28275_, _11887_, _10661_);
  or (_28276_, _28275_, _12412_);
  or (_28277_, _28276_, _28274_);
  nor (_28278_, _12441_, \oc8051_golden_model_1.DPH [2]);
  nor (_28279_, _28278_, _12442_);
  or (_28280_, _28279_, _12413_);
  and (_28281_, _28280_, _06636_);
  and (_28282_, _28281_, _28277_);
  and (_28285_, _11887_, _06088_);
  or (_28286_, _28285_, _28282_);
  nand (_28287_, _07187_, _05569_);
  and (_28288_, _28287_, _28286_);
  or (_28289_, _28143_, _11071_);
  or (_28290_, _11887_, _12459_);
  and (_28291_, _28290_, _12453_);
  and (_28292_, _28291_, _28289_);
  or (_28293_, _28292_, _12006_);
  or (_28294_, _28293_, _28288_);
  or (_28296_, _28124_, _12007_);
  and (_28297_, _28296_, _12466_);
  and (_28298_, _28297_, _28294_);
  nor (_28299_, _12466_, _14664_);
  or (_28300_, _28299_, _06112_);
  or (_28301_, _28300_, _28298_);
  nand (_28302_, _12044_, _06112_);
  and (_28303_, _28302_, _28301_);
  or (_28304_, _28303_, _06284_);
  nand (_28305_, _14664_, _06284_);
  nor (_28307_, _12476_, _05727_);
  and (_28308_, _28307_, _28305_);
  and (_28309_, _28308_, _28304_);
  or (_28310_, _28143_, _12459_);
  or (_28311_, _11887_, _11071_);
  and (_28312_, _28311_, _12476_);
  and (_28313_, _28312_, _28310_);
  or (_28314_, _28313_, _12481_);
  or (_28315_, _28314_, _28309_);
  or (_28316_, _28124_, _12002_);
  and (_28318_, _28316_, _10742_);
  and (_28319_, _28318_, _28315_);
  nor (_28320_, _14664_, _10742_);
  or (_28321_, _28320_, _06108_);
  or (_28322_, _28321_, _28319_);
  nand (_28323_, _12044_, _06108_);
  and (_28324_, _28323_, _28322_);
  or (_28325_, _28324_, _06277_);
  nand (_28326_, _14664_, _06277_);
  and (_28327_, _28326_, _27690_);
  and (_28329_, _28327_, _28325_);
  or (_28330_, _28143_, \oc8051_golden_model_1.PSW [7]);
  or (_28331_, _11887_, _10606_);
  and (_28332_, _28331_, _12497_);
  and (_28333_, _28332_, _28330_);
  or (_28334_, _28333_, _12502_);
  or (_28335_, _28334_, _28329_);
  or (_28336_, _28124_, _11993_);
  and (_28337_, _28336_, _11986_);
  and (_28338_, _28337_, _28335_);
  nor (_28340_, _14664_, _11986_);
  or (_28341_, _28340_, _06130_);
  or (_28342_, _28341_, _28338_);
  nand (_28343_, _12044_, _06130_);
  and (_28344_, _28343_, _28342_);
  or (_28345_, _28344_, _06292_);
  nand (_28346_, _14664_, _06292_);
  and (_28347_, _28346_, _27484_);
  and (_28348_, _28347_, _28345_);
  or (_28349_, _28143_, _10606_);
  or (_28351_, _11887_, \oc8051_golden_model_1.PSW [7]);
  and (_28352_, _28351_, _11982_);
  and (_28353_, _28352_, _28349_);
  or (_28354_, _28353_, _12525_);
  or (_28355_, _28354_, _28348_);
  or (_28356_, _28124_, _12523_);
  and (_28357_, _28356_, _10825_);
  and (_28358_, _28357_, _28355_);
  nor (_28359_, _14664_, _10825_);
  or (_28360_, _28359_, _10854_);
  or (_28362_, _28360_, _28358_);
  or (_28363_, _28124_, _10855_);
  and (_28364_, _28363_, _28362_);
  or (_28365_, _28364_, _06298_);
  nand (_28366_, _07530_, _06298_);
  and (_28367_, _28366_, _28056_);
  and (_28368_, _28367_, _28365_);
  or (_28369_, _28133_, _12723_);
  or (_28370_, _12043_, _12722_);
  and (_28371_, _28370_, _06129_);
  and (_28373_, _28371_, _28369_);
  or (_28374_, _28373_, _12541_);
  or (_28375_, _28374_, _28368_);
  or (_28376_, _28124_, _11872_);
  and (_28377_, _28376_, _10975_);
  and (_28378_, _28377_, _28375_);
  nor (_28379_, _14664_, _10975_);
  or (_28380_, _28379_, _11015_);
  or (_28381_, _28380_, _28378_);
  or (_28382_, _28124_, _11016_);
  and (_28384_, _28382_, _28381_);
  or (_28385_, _28384_, _06049_);
  nand (_28386_, _07530_, _06049_);
  and (_28387_, _28386_, _28077_);
  and (_28388_, _28387_, _28385_);
  or (_28389_, _28133_, _12722_);
  nand (_28390_, _12044_, _12722_);
  and (_28391_, _28390_, _28389_);
  and (_28392_, _28391_, _06126_);
  or (_28393_, _28392_, _12750_);
  or (_28395_, _28393_, _28388_);
  or (_28396_, _28124_, _12749_);
  and (_28397_, _28396_, _28395_);
  or (_28398_, _28397_, _06316_);
  nand (_28399_, _14664_, _06316_);
  and (_28400_, _28399_, _12756_);
  and (_28401_, _28400_, _28398_);
  and (_28402_, _28124_, _25353_);
  or (_28403_, _28402_, _06127_);
  or (_28404_, _28403_, _28401_);
  nand (_28406_, _06403_, _06127_);
  and (_28407_, _28406_, _27775_);
  and (_28408_, _28407_, _28404_);
  and (_28409_, _28391_, _05652_);
  or (_28410_, _28409_, _12772_);
  or (_28411_, _28410_, _28408_);
  or (_28412_, _28124_, _12771_);
  and (_28413_, _28412_, _28411_);
  or (_28414_, _28413_, _06047_);
  nand (_28415_, _14664_, _06047_);
  and (_28417_, _28415_, _12779_);
  and (_28418_, _28417_, _28414_);
  and (_28419_, _28124_, _26405_);
  or (_28420_, _28419_, _06119_);
  or (_28421_, _28420_, _28418_);
  nand (_28422_, _06403_, _06119_);
  and (_28423_, _28422_, _27789_);
  and (_28424_, _28423_, _28421_);
  and (_28425_, _28124_, _12789_);
  or (_28426_, _28425_, _28424_);
  or (_28428_, _28426_, _01340_);
  or (_28429_, _01336_, \oc8051_golden_model_1.PC [10]);
  and (_28430_, _28429_, _42882_);
  and (_43428_, _28430_, _28428_);
  nor (_28431_, _11864_, \oc8051_golden_model_1.PC [11]);
  nor (_28432_, _28431_, _11865_);
  or (_28433_, _28432_, _11872_);
  or (_28434_, _28432_, _12523_);
  or (_28435_, _28432_, _11993_);
  or (_28436_, _28432_, _12007_);
  nor (_28438_, _12037_, _05669_);
  nor (_28439_, _28131_, _12045_);
  and (_28440_, _28439_, _12040_);
  nor (_28441_, _28439_, _12040_);
  or (_28442_, _28441_, _28440_);
  or (_28443_, _28442_, _12172_);
  or (_28444_, _12174_, _12036_);
  and (_28445_, _28444_, _06104_);
  and (_28446_, _28445_, _28443_);
  and (_28447_, _11891_, _06219_);
  or (_28449_, _12179_, _11891_);
  or (_28450_, _12187_, _12036_);
  or (_28451_, _28442_, _12189_);
  and (_28452_, _28451_, _06102_);
  and (_28453_, _28452_, _28450_);
  nor (_28454_, _28140_, _11888_);
  nor (_28455_, _28454_, _11894_);
  and (_28456_, _28454_, _11894_);
  or (_28457_, _28456_, _28455_);
  and (_28458_, _28457_, _12199_);
  and (_28460_, _12197_, _11891_);
  or (_28461_, _28460_, _08383_);
  or (_28462_, _28461_, _28458_);
  or (_28463_, _28432_, _12215_);
  or (_28464_, _11891_, _07233_);
  or (_28465_, _11891_, _06939_);
  or (_28466_, _06938_, \oc8051_golden_model_1.PC [11]);
  or (_28467_, _28466_, _07250_);
  and (_28468_, _28467_, _28465_);
  nand (_28469_, _24785_, _25758_);
  or (_28471_, _28469_, _28468_);
  and (_28472_, _28471_, _28464_);
  and (_28473_, _28472_, _28463_);
  or (_28474_, _28473_, _08384_);
  and (_28475_, _28474_, _12219_);
  and (_28476_, _28475_, _28462_);
  or (_28477_, _28476_, _28453_);
  and (_28478_, _28477_, _12182_);
  and (_28479_, _28432_, _12226_);
  or (_28480_, _28479_, _12224_);
  or (_28482_, _28480_, _28478_);
  and (_28483_, _28482_, _28449_);
  or (_28484_, _28483_, _12232_);
  or (_28485_, _28432_, _12231_);
  and (_28486_, _28485_, _06220_);
  and (_28487_, _28486_, _28484_);
  or (_28488_, _28487_, _28447_);
  and (_28489_, _28488_, _12239_);
  and (_28490_, _28432_, _12241_);
  or (_28491_, _28490_, _12246_);
  or (_28493_, _28491_, _28489_);
  or (_28494_, _12245_, _11891_);
  and (_28495_, _28494_, _28493_);
  or (_28496_, _28495_, _12256_);
  or (_28497_, _28442_, _12289_);
  nand (_28498_, _12289_, _12037_);
  and (_28499_, _28498_, _28497_);
  or (_28500_, _28499_, _12255_);
  and (_28501_, _28500_, _12258_);
  and (_28502_, _28501_, _28496_);
  or (_28504_, _28502_, _06121_);
  or (_28505_, _28504_, _28446_);
  and (_28506_, _12310_, _12036_);
  and (_28507_, _28442_, _12312_);
  or (_28508_, _28507_, _06509_);
  or (_28509_, _28508_, _28506_);
  and (_28510_, _28509_, _12298_);
  and (_28511_, _28510_, _28505_);
  or (_28512_, _28442_, _12329_);
  nand (_28513_, _12329_, _12037_);
  and (_28515_, _28513_, _06115_);
  and (_28516_, _28515_, _28512_);
  or (_28517_, _28516_, _28511_);
  and (_28518_, _28517_, _12013_);
  nand (_28519_, _28432_, _12012_);
  nand (_28520_, _28519_, _12345_);
  or (_28521_, _28520_, _28518_);
  or (_28522_, _12345_, _11891_);
  and (_28523_, _28522_, _12351_);
  and (_28524_, _28523_, _28521_);
  and (_28526_, _28432_, _12355_);
  or (_28527_, _28526_, _12358_);
  or (_28528_, _28527_, _28524_);
  or (_28529_, _12357_, _11891_);
  and (_28530_, _28529_, _12362_);
  and (_28531_, _28530_, _28528_);
  and (_28532_, _28432_, _12368_);
  or (_28533_, _28532_, _12367_);
  or (_28534_, _28533_, _28531_);
  or (_28535_, _11891_, _12366_);
  and (_28537_, _28535_, _05675_);
  and (_28538_, _28537_, _28534_);
  nand (_28539_, _28432_, _05676_);
  nand (_28540_, _28539_, _12376_);
  or (_28541_, _28540_, _28538_);
  or (_28542_, _12376_, _11891_);
  and (_28543_, _28542_, _06111_);
  and (_28544_, _28543_, _28541_);
  nand (_28545_, _12036_, _06110_);
  nand (_28546_, _28545_, _09817_);
  or (_28548_, _28546_, _28544_);
  or (_28549_, _11891_, _09817_);
  and (_28550_, _28549_, _05669_);
  and (_28551_, _28550_, _28548_);
  or (_28552_, _28551_, _28438_);
  and (_28553_, _28552_, _12389_);
  and (_28554_, _28432_, _12393_);
  or (_28555_, _28554_, _12392_);
  or (_28556_, _28555_, _28553_);
  or (_28557_, _12391_, _11891_);
  and (_28559_, _28557_, _12398_);
  and (_28560_, _28559_, _28556_);
  and (_28561_, _28457_, _12397_);
  or (_28562_, _28561_, _08743_);
  or (_28563_, _28562_, _28560_);
  or (_28564_, _11891_, _08742_);
  and (_28565_, _28564_, _06020_);
  and (_28566_, _28565_, _28563_);
  and (_28567_, _12036_, _06019_);
  or (_28568_, _28567_, _10661_);
  or (_28570_, _28568_, _28566_);
  or (_28571_, _11891_, _10662_);
  and (_28572_, _28571_, _12413_);
  and (_28573_, _28572_, _28570_);
  or (_28574_, _12442_, \oc8051_golden_model_1.DPH [3]);
  nor (_28575_, _12443_, _12413_);
  and (_28576_, _28575_, _28574_);
  or (_28577_, _28576_, _12416_);
  or (_28578_, _28577_, _28573_);
  or (_28579_, _12415_, _11891_);
  and (_28581_, _28579_, _12454_);
  and (_28582_, _28581_, _28578_);
  or (_28583_, _28457_, _11071_);
  or (_28584_, _11891_, _12459_);
  and (_28585_, _28584_, _12453_);
  and (_28586_, _28585_, _28583_);
  or (_28587_, _28586_, _12006_);
  or (_28588_, _28587_, _28582_);
  and (_28589_, _28588_, _28436_);
  or (_28590_, _28589_, _12467_);
  or (_28592_, _12466_, _11891_);
  and (_28593_, _28592_, _08751_);
  and (_28594_, _28593_, _28590_);
  nand (_28595_, _12036_, _06112_);
  nand (_28596_, _28595_, _12473_);
  or (_28597_, _28596_, _28594_);
  or (_28598_, _12473_, _11891_);
  and (_28599_, _28598_, _12477_);
  and (_28600_, _28599_, _28597_);
  or (_28601_, _28457_, _12459_);
  or (_28603_, _11891_, _11071_);
  and (_28604_, _28603_, _12476_);
  and (_28605_, _28604_, _28601_);
  or (_28606_, _28605_, _28600_);
  and (_28607_, _28606_, _12002_);
  and (_28608_, _28432_, _12481_);
  or (_28609_, _28608_, _10743_);
  or (_28610_, _28609_, _28607_);
  or (_28611_, _11891_, _10742_);
  and (_28612_, _28611_, _07032_);
  and (_28614_, _28612_, _28610_);
  nand (_28615_, _12036_, _06108_);
  nand (_28616_, _28615_, _12494_);
  or (_28617_, _28616_, _28614_);
  or (_28618_, _12494_, _11891_);
  and (_28619_, _28618_, _12498_);
  and (_28620_, _28619_, _28617_);
  or (_28621_, _28457_, \oc8051_golden_model_1.PSW [7]);
  or (_28622_, _11891_, _10606_);
  and (_28623_, _28622_, _12497_);
  and (_28624_, _28623_, _28621_);
  or (_28625_, _28624_, _12502_);
  or (_28626_, _28625_, _28620_);
  and (_28627_, _28626_, _28435_);
  or (_28628_, _28627_, _11987_);
  or (_28629_, _11891_, _11986_);
  and (_28630_, _28629_, _08777_);
  and (_28631_, _28630_, _28628_);
  nand (_28632_, _12036_, _06130_);
  nand (_28633_, _28632_, _12515_);
  or (_28636_, _28633_, _28631_);
  or (_28637_, _12515_, _11891_);
  and (_28638_, _28637_, _12518_);
  and (_28639_, _28638_, _28636_);
  or (_28640_, _28457_, _10606_);
  or (_28641_, _11891_, \oc8051_golden_model_1.PSW [7]);
  and (_28642_, _28641_, _11982_);
  and (_28643_, _28642_, _28640_);
  or (_28644_, _28643_, _12525_);
  or (_28645_, _28644_, _28639_);
  and (_28647_, _28645_, _28434_);
  or (_28648_, _28647_, _10826_);
  or (_28649_, _11891_, _10825_);
  and (_28650_, _28649_, _10855_);
  and (_28651_, _28650_, _28648_);
  and (_28652_, _28432_, _10854_);
  or (_28653_, _28652_, _06298_);
  or (_28654_, _28653_, _28651_);
  nand (_28655_, _07353_, _06298_);
  and (_28656_, _28655_, _28654_);
  or (_28658_, _28656_, _05732_);
  or (_28659_, _11891_, _05734_);
  and (_28660_, _28659_, _06306_);
  and (_28661_, _28660_, _28658_);
  or (_28662_, _28442_, _12723_);
  or (_28663_, _12036_, _12722_);
  and (_28664_, _28663_, _06129_);
  and (_28665_, _28664_, _28662_);
  or (_28666_, _28665_, _12541_);
  or (_28667_, _28666_, _28661_);
  and (_28669_, _28667_, _28433_);
  or (_28670_, _28669_, _10976_);
  or (_28671_, _11891_, _10975_);
  and (_28672_, _28671_, _11016_);
  and (_28673_, _28672_, _28670_);
  and (_28674_, _28432_, _11015_);
  or (_28675_, _28674_, _06049_);
  or (_28676_, _28675_, _28673_);
  nand (_28677_, _07353_, _06049_);
  and (_28678_, _28677_, _28676_);
  or (_28680_, _28678_, _05747_);
  or (_28681_, _11891_, _05748_);
  and (_28682_, _28681_, _06704_);
  and (_28683_, _28682_, _28680_);
  or (_28684_, _28442_, _12722_);
  nand (_28685_, _12037_, _12722_);
  and (_28686_, _28685_, _28684_);
  and (_28687_, _28686_, _06126_);
  or (_28688_, _28687_, _12750_);
  or (_28689_, _28688_, _28683_);
  or (_28691_, _28432_, _12749_);
  and (_28692_, _28691_, _06718_);
  and (_28693_, _28692_, _28689_);
  nand (_28694_, _11891_, _06316_);
  nand (_28695_, _28694_, _12756_);
  or (_28696_, _28695_, _28693_);
  or (_28697_, _28432_, _12756_);
  and (_28698_, _28697_, _09200_);
  and (_28699_, _28698_, _28696_);
  nor (_28700_, _09200_, _05983_);
  or (_28702_, _28700_, _05752_);
  or (_28703_, _28702_, _28699_);
  or (_28704_, _11891_, _12766_);
  and (_28705_, _28704_, _05653_);
  and (_28706_, _28705_, _28703_);
  and (_28707_, _28686_, _05652_);
  or (_28708_, _28707_, _12772_);
  or (_28709_, _28708_, _28706_);
  or (_28710_, _28432_, _12771_);
  and (_28711_, _28710_, _06048_);
  and (_28713_, _28711_, _28709_);
  nand (_28714_, _11891_, _06047_);
  nand (_28715_, _28714_, _12779_);
  or (_28716_, _28715_, _28713_);
  or (_28717_, _28432_, _12779_);
  and (_28718_, _28717_, _12782_);
  and (_28719_, _28718_, _28716_);
  nor (_28720_, _12782_, _05983_);
  or (_28721_, _28720_, _05751_);
  or (_28722_, _28721_, _28719_);
  or (_28724_, _11891_, _12791_);
  and (_28725_, _28724_, _12790_);
  and (_28726_, _28725_, _28722_);
  and (_28727_, _28432_, _12789_);
  or (_28728_, _28727_, _28726_);
  or (_28729_, _28728_, _01340_);
  or (_28730_, _01336_, \oc8051_golden_model_1.PC [11]);
  and (_28731_, _28730_, _42882_);
  and (_43429_, _28731_, _28729_);
  and (_28732_, _15062_, _05752_);
  and (_28734_, _11884_, _10606_);
  and (_28735_, _11967_, _11964_);
  nor (_28736_, _28735_, _11968_);
  and (_28737_, _28736_, \oc8051_golden_model_1.PSW [7]);
  or (_28738_, _28737_, _28734_);
  and (_28739_, _28738_, _11982_);
  nor (_28740_, _11884_, _08742_);
  nor (_28741_, _12033_, _05669_);
  and (_28742_, _12129_, _12126_);
  nor (_28743_, _28742_, _12130_);
  and (_28745_, _28743_, _12174_);
  and (_28746_, _12172_, _12032_);
  nor (_28747_, _28746_, _28745_);
  nor (_28748_, _28747_, _12258_);
  nand (_28749_, _12289_, _12033_);
  or (_28750_, _28743_, _12289_);
  and (_28751_, _28750_, _12256_);
  and (_28752_, _28751_, _28749_);
  and (_28753_, _11862_, _09202_);
  and (_28754_, _28753_, \oc8051_golden_model_1.PC [11]);
  and (_28756_, _28754_, \oc8051_golden_model_1.PC [12]);
  nor (_28757_, _28754_, \oc8051_golden_model_1.PC [12]);
  nor (_28758_, _28757_, _28756_);
  nor (_28759_, _28758_, _12225_);
  or (_28760_, _12187_, _12033_);
  not (_28761_, _28743_);
  or (_28762_, _28761_, _12189_);
  and (_28763_, _28762_, _06102_);
  and (_28764_, _28763_, _28760_);
  nor (_28765_, _12199_, _11884_);
  or (_28767_, _28736_, _12197_);
  nand (_28768_, _28767_, _08384_);
  or (_28769_, _28768_, _28765_);
  nor (_28770_, _28758_, _12215_);
  nor (_28771_, _12206_, _11884_);
  or (_28772_, _06938_, \oc8051_golden_model_1.PC [12]);
  or (_28773_, _28772_, _12208_);
  nor (_28774_, _28773_, _07250_);
  or (_28775_, _28774_, _28771_);
  and (_28776_, _28775_, _12205_);
  or (_28778_, _28776_, _08384_);
  or (_28779_, _28778_, _28770_);
  and (_28780_, _28779_, _12219_);
  and (_28781_, _28780_, _28769_);
  or (_28782_, _28781_, _28764_);
  and (_28783_, _28782_, _12182_);
  or (_28784_, _28783_, _28759_);
  nand (_28785_, _28784_, _12179_);
  nor (_28786_, _12179_, _11884_);
  nor (_28787_, _28786_, _12232_);
  nand (_28789_, _28787_, _28785_);
  not (_28790_, _28758_);
  nor (_28791_, _28790_, _12231_);
  nor (_28792_, _28791_, _06219_);
  nand (_28793_, _28792_, _28789_);
  and (_28794_, _15062_, _06219_);
  nor (_28795_, _28794_, _12241_);
  nand (_28796_, _28795_, _28793_);
  nor (_28797_, _28790_, _12239_);
  nor (_28798_, _28797_, _12246_);
  nand (_28800_, _28798_, _28796_);
  nor (_28801_, _12245_, _11884_);
  not (_28802_, _28801_);
  and (_28803_, _28802_, _12255_);
  and (_28804_, _28803_, _28800_);
  or (_28805_, _28804_, _28752_);
  and (_28806_, _28805_, _12258_);
  or (_28807_, _28806_, _28748_);
  and (_28808_, _28807_, _06509_);
  and (_28809_, _12310_, _12032_);
  nor (_28811_, _28761_, _12310_);
  nor (_28812_, _28811_, _28809_);
  nor (_28813_, _28812_, _06509_);
  or (_28814_, _28813_, _28808_);
  nand (_28815_, _28814_, _12298_);
  nand (_28816_, _12329_, _12032_);
  nand (_28817_, _28743_, _26881_);
  and (_28818_, _28817_, _28816_);
  or (_28819_, _28818_, _12298_);
  nand (_28820_, _28819_, _28815_);
  nand (_28822_, _28820_, _12013_);
  and (_28823_, _28758_, _12012_);
  not (_28824_, _28823_);
  and (_28825_, _28824_, _12345_);
  nand (_28826_, _28825_, _28822_);
  nor (_28827_, _12345_, _11884_);
  nor (_28828_, _28827_, _12355_);
  nand (_28829_, _28828_, _28826_);
  nor (_28830_, _28790_, _12351_);
  nor (_28831_, _28830_, _12358_);
  nand (_28833_, _28831_, _28829_);
  nor (_28834_, _12357_, _11884_);
  nor (_28835_, _28834_, _12368_);
  nand (_28836_, _28835_, _28833_);
  or (_28837_, _28790_, _12362_);
  and (_28838_, _28837_, _12366_);
  nand (_28839_, _28838_, _28836_);
  nor (_28840_, _11884_, _12366_);
  nor (_28841_, _28840_, _05676_);
  nand (_28842_, _28841_, _28839_);
  nor (_28844_, _28790_, _05675_);
  not (_28845_, _28844_);
  and (_28846_, _28845_, _12376_);
  nand (_28847_, _28846_, _28842_);
  nor (_28848_, _12376_, _11884_);
  nor (_28849_, _28848_, _06110_);
  nand (_28850_, _28849_, _28847_);
  and (_28851_, _12032_, _06110_);
  nor (_28852_, _28851_, _09818_);
  nand (_28853_, _28852_, _28850_);
  nor (_28855_, _11884_, _09817_);
  nor (_28856_, _28855_, _09833_);
  and (_28857_, _28856_, _28853_);
  or (_28858_, _28857_, _28741_);
  nand (_28859_, _28858_, _12389_);
  nor (_28860_, _28790_, _12389_);
  nor (_28861_, _28860_, _12392_);
  nand (_28862_, _28861_, _28859_);
  nor (_28863_, _12391_, _11884_);
  nor (_28864_, _28863_, _12397_);
  nand (_28866_, _28864_, _28862_);
  and (_28867_, _28736_, _12397_);
  nor (_28868_, _28867_, _08743_);
  and (_28869_, _28868_, _28866_);
  or (_28870_, _28869_, _28740_);
  nand (_28871_, _28870_, _06020_);
  and (_28872_, _12033_, _06019_);
  nor (_28873_, _28872_, _10661_);
  and (_28874_, _28873_, _28871_);
  and (_28875_, _11884_, _10661_);
  or (_28877_, _28875_, _28874_);
  nand (_28878_, _28877_, _12413_);
  nor (_28879_, _12443_, \oc8051_golden_model_1.DPH [4]);
  nor (_28880_, _28879_, _12444_);
  and (_28881_, _28880_, _12412_);
  nor (_28882_, _28881_, _12416_);
  nand (_28883_, _28882_, _28878_);
  nor (_28884_, _12415_, _11884_);
  nor (_28885_, _28884_, _12453_);
  and (_28886_, _28885_, _28883_);
  and (_28888_, _11884_, _11071_);
  and (_28889_, _28736_, _12459_);
  or (_28890_, _28889_, _28888_);
  and (_28891_, _28890_, _12453_);
  or (_28892_, _28891_, _28886_);
  nand (_28893_, _28892_, _12007_);
  and (_28894_, _28758_, _12006_);
  nor (_28895_, _28894_, _12467_);
  nand (_28896_, _28895_, _28893_);
  nor (_28897_, _12466_, _11884_);
  nor (_28899_, _28897_, _06112_);
  nand (_28900_, _28899_, _28896_);
  not (_28901_, _12473_);
  and (_28902_, _12032_, _06112_);
  nor (_28903_, _28902_, _28901_);
  nand (_28904_, _28903_, _28900_);
  nor (_28905_, _12473_, _11884_);
  nor (_28906_, _28905_, _12476_);
  and (_28907_, _28906_, _28904_);
  and (_28908_, _11884_, _12459_);
  and (_28910_, _28736_, _11071_);
  or (_28911_, _28910_, _28908_);
  and (_28912_, _28911_, _12476_);
  or (_28913_, _28912_, _28907_);
  nand (_28914_, _28913_, _12002_);
  nor (_28915_, _28790_, _12002_);
  nor (_28916_, _28915_, _10743_);
  nand (_28917_, _28916_, _28914_);
  nor (_28918_, _11884_, _10742_);
  nor (_28919_, _28918_, _06108_);
  nand (_28921_, _28919_, _28917_);
  not (_28922_, _12494_);
  and (_28923_, _12032_, _06108_);
  nor (_28924_, _28923_, _28922_);
  nand (_28925_, _28924_, _28921_);
  nor (_28926_, _12494_, _11884_);
  nor (_28927_, _28926_, _12497_);
  and (_28928_, _28927_, _28925_);
  and (_28929_, _11884_, \oc8051_golden_model_1.PSW [7]);
  and (_28930_, _28736_, _10606_);
  or (_28932_, _28930_, _28929_);
  and (_28933_, _28932_, _12497_);
  or (_28934_, _28933_, _28928_);
  nand (_28935_, _28934_, _11993_);
  nor (_28936_, _28790_, _11993_);
  nor (_28937_, _28936_, _11987_);
  nand (_28938_, _28937_, _28935_);
  nor (_28939_, _11884_, _11986_);
  nor (_28940_, _28939_, _06130_);
  nand (_28941_, _28940_, _28938_);
  not (_28943_, _12515_);
  and (_28944_, _12032_, _06130_);
  nor (_28945_, _28944_, _28943_);
  nand (_28946_, _28945_, _28941_);
  nor (_28947_, _12515_, _11884_);
  nor (_28948_, _28947_, _11982_);
  and (_28949_, _28948_, _28946_);
  or (_28950_, _28949_, _28739_);
  nand (_28951_, _28950_, _12523_);
  nor (_28952_, _28790_, _12523_);
  nor (_28954_, _28952_, _10826_);
  nand (_28955_, _28954_, _28951_);
  nor (_28956_, _11884_, _10825_);
  nor (_28957_, _28956_, _10854_);
  nand (_28958_, _28957_, _28955_);
  and (_28959_, _28758_, _10854_);
  nor (_28960_, _28959_, _06298_);
  and (_28961_, _28960_, _28958_);
  and (_28962_, _08270_, _06298_);
  or (_28963_, _28962_, _28961_);
  nand (_28965_, _28963_, _05734_);
  and (_28966_, _15062_, _05732_);
  nor (_28967_, _28966_, _06129_);
  and (_28968_, _28967_, _28965_);
  and (_28969_, _28743_, _12722_);
  nor (_28970_, _12033_, _12722_);
  nor (_28971_, _28970_, _28969_);
  nor (_28972_, _28971_, _06306_);
  or (_28973_, _28972_, _28968_);
  nand (_28974_, _28973_, _11872_);
  nor (_28976_, _28790_, _11872_);
  nor (_28977_, _28976_, _10976_);
  nand (_28978_, _28977_, _28974_);
  nor (_28979_, _11884_, _10975_);
  nor (_28980_, _28979_, _11015_);
  nand (_28981_, _28980_, _28978_);
  and (_28982_, _28758_, _11015_);
  nor (_28983_, _28982_, _06049_);
  nand (_28984_, _28983_, _28981_);
  and (_28985_, _08270_, _06049_);
  nor (_28987_, _28985_, _05747_);
  and (_28988_, _28987_, _28984_);
  and (_28989_, _11884_, _05747_);
  or (_28990_, _28989_, _06126_);
  or (_28991_, _28990_, _28988_);
  nor (_28992_, _28743_, _12722_);
  and (_28993_, _12033_, _12722_);
  nor (_28994_, _28993_, _28992_);
  nor (_28995_, _28994_, _06704_);
  nor (_28996_, _28995_, _12750_);
  nand (_28997_, _28996_, _28991_);
  nor (_28998_, _28790_, _12749_);
  nor (_28999_, _28998_, _06316_);
  nand (_29000_, _28999_, _28997_);
  and (_29001_, _15062_, _06316_);
  nor (_29002_, _29001_, _25353_);
  and (_29003_, _29002_, _29000_);
  nor (_29004_, _28790_, _12756_);
  or (_29005_, _29004_, _06127_);
  nor (_29006_, _29005_, _29003_);
  and (_29009_, _06758_, _06127_);
  or (_29010_, _29009_, _29006_);
  and (_29011_, _29010_, _12766_);
  or (_29012_, _29011_, _28732_);
  nand (_29013_, _29012_, _05653_);
  nor (_29014_, _28994_, _05653_);
  nor (_29015_, _29014_, _12772_);
  nand (_29016_, _29015_, _29013_);
  nor (_29017_, _28790_, _12771_);
  nor (_29018_, _29017_, _06047_);
  nand (_29020_, _29018_, _29016_);
  and (_29021_, _15062_, _06047_);
  nor (_29022_, _29021_, _26405_);
  nand (_29023_, _29022_, _29020_);
  nor (_29024_, _28790_, _12779_);
  nor (_29025_, _29024_, _06119_);
  nand (_29026_, _29025_, _29023_);
  and (_29027_, _06758_, _06119_);
  nor (_29028_, _29027_, _05751_);
  nand (_29029_, _29028_, _29026_);
  and (_29031_, _11884_, _05751_);
  nor (_29032_, _29031_, _12789_);
  and (_29033_, _29032_, _29029_);
  and (_29034_, _28790_, _12789_);
  nor (_29035_, _29034_, _29033_);
  or (_29036_, _29035_, _01340_);
  or (_29037_, _01336_, \oc8051_golden_model_1.PC [12]);
  and (_29038_, _29037_, _42882_);
  and (_43430_, _29038_, _29036_);
  and (_29039_, _28756_, \oc8051_golden_model_1.PC [13]);
  nor (_29041_, _28756_, \oc8051_golden_model_1.PC [13]);
  nor (_29042_, _29041_, _29039_);
  or (_29043_, _29042_, _11872_);
  or (_29044_, _29042_, _12523_);
  or (_29045_, _29042_, _11993_);
  or (_29046_, _11882_, _11881_);
  not (_29047_, _29046_);
  nor (_29048_, _29047_, _11969_);
  and (_29049_, _29047_, _11969_);
  or (_29050_, _29049_, _29048_);
  or (_29052_, _29050_, _11071_);
  or (_29053_, _11880_, _12459_);
  and (_29054_, _29053_, _12453_);
  and (_29055_, _29054_, _29052_);
  or (_29056_, _11880_, _08742_);
  nor (_29057_, _12028_, _05669_);
  or (_29058_, _12030_, _12029_);
  not (_29059_, _29058_);
  nor (_29060_, _29059_, _12131_);
  and (_29061_, _29059_, _12131_);
  or (_29063_, _29061_, _29060_);
  or (_29064_, _29063_, _12172_);
  nor (_29065_, _12174_, _12027_);
  nor (_29066_, _29065_, _12258_);
  and (_29067_, _29066_, _29064_);
  and (_29068_, _11880_, _06219_);
  or (_29069_, _12179_, _11880_);
  or (_29070_, _12187_, _12027_);
  or (_29071_, _29063_, _12189_);
  and (_29072_, _29071_, _06102_);
  and (_29074_, _29072_, _29070_);
  and (_29075_, _29050_, _12199_);
  and (_29076_, _12197_, _11880_);
  or (_29077_, _29076_, _08383_);
  or (_29078_, _29077_, _29075_);
  or (_29079_, _29042_, _12215_);
  or (_29080_, _12206_, _11880_);
  or (_29081_, _06530_, \oc8051_golden_model_1.PC [13]);
  or (_29082_, _29081_, _06938_);
  nor (_29083_, _29082_, _07250_);
  nand (_29085_, _29083_, _24785_);
  and (_29086_, _29085_, _29080_);
  and (_29087_, _29086_, _29079_);
  or (_29088_, _29087_, _08384_);
  and (_29089_, _29088_, _12219_);
  and (_29090_, _29089_, _29078_);
  or (_29091_, _29090_, _29074_);
  and (_29092_, _29091_, _12182_);
  not (_29093_, _29042_);
  nor (_29094_, _29093_, _12225_);
  or (_29096_, _29094_, _12224_);
  or (_29097_, _29096_, _29092_);
  and (_29098_, _29097_, _29069_);
  or (_29099_, _29098_, _12232_);
  or (_29100_, _29042_, _12231_);
  and (_29101_, _29100_, _06220_);
  and (_29102_, _29101_, _29099_);
  or (_29103_, _29102_, _29068_);
  and (_29104_, _29103_, _12239_);
  or (_29105_, _29093_, _12239_);
  nand (_29107_, _29105_, _12245_);
  or (_29108_, _29107_, _29104_);
  or (_29109_, _12245_, _11880_);
  and (_29110_, _29109_, _29108_);
  or (_29111_, _29110_, _12256_);
  or (_29112_, _29063_, _12289_);
  nand (_29113_, _12289_, _12028_);
  and (_29114_, _29113_, _29112_);
  or (_29115_, _29114_, _12255_);
  and (_29116_, _29115_, _12258_);
  and (_29118_, _29116_, _29111_);
  or (_29119_, _29118_, _06121_);
  or (_29120_, _29119_, _29067_);
  and (_29121_, _12310_, _12027_);
  and (_29122_, _29063_, _12312_);
  or (_29123_, _29122_, _06509_);
  or (_29124_, _29123_, _29121_);
  and (_29125_, _29124_, _12298_);
  and (_29126_, _29125_, _29120_);
  or (_29127_, _29063_, _12329_);
  nand (_29129_, _12329_, _12028_);
  and (_29130_, _29129_, _06115_);
  and (_29131_, _29130_, _29127_);
  or (_29132_, _29131_, _29126_);
  and (_29133_, _29132_, _12013_);
  nand (_29134_, _29042_, _12012_);
  nand (_29135_, _29134_, _12345_);
  or (_29136_, _29135_, _29133_);
  or (_29137_, _12345_, _11880_);
  and (_29138_, _29137_, _12351_);
  and (_29140_, _29138_, _29136_);
  nor (_29141_, _29093_, _12351_);
  or (_29142_, _29141_, _12358_);
  or (_29143_, _29142_, _29140_);
  or (_29144_, _12357_, _11880_);
  and (_29145_, _29144_, _12362_);
  and (_29146_, _29145_, _29143_);
  or (_29147_, _29093_, _12362_);
  nand (_29148_, _29147_, _12366_);
  or (_29149_, _29148_, _29146_);
  or (_29151_, _11880_, _12366_);
  and (_29152_, _29151_, _05675_);
  and (_29153_, _29152_, _29149_);
  or (_29154_, _29093_, _05675_);
  nand (_29155_, _29154_, _12376_);
  or (_29156_, _29155_, _29153_);
  or (_29157_, _12376_, _11880_);
  and (_29158_, _29157_, _06111_);
  and (_29159_, _29158_, _29156_);
  nand (_29160_, _12027_, _06110_);
  nand (_29162_, _29160_, _09817_);
  or (_29163_, _29162_, _29159_);
  or (_29164_, _11880_, _09817_);
  and (_29165_, _29164_, _05669_);
  and (_29166_, _29165_, _29163_);
  or (_29167_, _29166_, _29057_);
  and (_29168_, _29167_, _12389_);
  nor (_29169_, _29093_, _12389_);
  or (_29170_, _29169_, _12392_);
  or (_29171_, _29170_, _29168_);
  or (_29173_, _12391_, _11880_);
  and (_29174_, _29173_, _12398_);
  and (_29175_, _29174_, _29171_);
  and (_29176_, _29050_, _12397_);
  or (_29177_, _29176_, _08743_);
  or (_29178_, _29177_, _29175_);
  and (_29179_, _29178_, _29056_);
  or (_29180_, _29179_, _06019_);
  nand (_29181_, _12028_, _06019_);
  and (_29182_, _29181_, _10662_);
  and (_29184_, _29182_, _29180_);
  and (_29185_, _11880_, _10661_);
  or (_29186_, _29185_, _29184_);
  and (_29187_, _29186_, _12413_);
  or (_29188_, _12444_, \oc8051_golden_model_1.DPH [5]);
  nor (_29189_, _12445_, _12413_);
  and (_29190_, _29189_, _29188_);
  or (_29191_, _29190_, _12416_);
  or (_29192_, _29191_, _29187_);
  or (_29193_, _12415_, _11880_);
  and (_29195_, _29193_, _12454_);
  and (_29196_, _29195_, _29192_);
  or (_29197_, _29196_, _29055_);
  and (_29198_, _29197_, _12007_);
  and (_29199_, _29042_, _12006_);
  or (_29200_, _29199_, _12467_);
  or (_29201_, _29200_, _29198_);
  or (_29202_, _12466_, _11880_);
  and (_29203_, _29202_, _08751_);
  and (_29204_, _29203_, _29201_);
  nand (_29206_, _12027_, _06112_);
  nand (_29207_, _29206_, _12473_);
  or (_29208_, _29207_, _29204_);
  or (_29209_, _12473_, _11880_);
  and (_29210_, _29209_, _12477_);
  and (_29211_, _29210_, _29208_);
  or (_29212_, _29050_, _12459_);
  or (_29213_, _11880_, _11071_);
  and (_29214_, _29213_, _12476_);
  and (_29215_, _29214_, _29212_);
  or (_29217_, _29215_, _29211_);
  and (_29218_, _29217_, _12002_);
  nor (_29219_, _29093_, _12002_);
  or (_29220_, _29219_, _10743_);
  or (_29221_, _29220_, _29218_);
  or (_29222_, _11880_, _10742_);
  and (_29223_, _29222_, _07032_);
  and (_29224_, _29223_, _29221_);
  nand (_29225_, _12027_, _06108_);
  nand (_29226_, _29225_, _12494_);
  or (_29228_, _29226_, _29224_);
  or (_29229_, _12494_, _11880_);
  and (_29230_, _29229_, _12498_);
  and (_29231_, _29230_, _29228_);
  or (_29232_, _29050_, \oc8051_golden_model_1.PSW [7]);
  or (_29233_, _11880_, _10606_);
  and (_29234_, _29233_, _12497_);
  and (_29235_, _29234_, _29232_);
  or (_29236_, _29235_, _12502_);
  or (_29237_, _29236_, _29231_);
  and (_29239_, _29237_, _29045_);
  or (_29240_, _29239_, _11987_);
  or (_29241_, _11880_, _11986_);
  and (_29242_, _29241_, _08777_);
  and (_29243_, _29242_, _29240_);
  nand (_29244_, _12027_, _06130_);
  nand (_29245_, _29244_, _12515_);
  or (_29246_, _29245_, _29243_);
  or (_29247_, _12515_, _11880_);
  and (_29248_, _29247_, _12518_);
  and (_29250_, _29248_, _29246_);
  or (_29251_, _29050_, _10606_);
  or (_29252_, _11880_, \oc8051_golden_model_1.PSW [7]);
  and (_29253_, _29252_, _11982_);
  and (_29254_, _29253_, _29251_);
  or (_29255_, _29254_, _12525_);
  or (_29256_, _29255_, _29250_);
  and (_29257_, _29256_, _29044_);
  or (_29258_, _29257_, _10826_);
  or (_29259_, _11880_, _10825_);
  and (_29261_, _29259_, _10855_);
  and (_29262_, _29261_, _29258_);
  and (_29263_, _29042_, _10854_);
  or (_29264_, _29263_, _06298_);
  or (_29265_, _29264_, _29262_);
  nand (_29266_, _07977_, _06298_);
  and (_29267_, _29266_, _29265_);
  or (_29268_, _29267_, _05732_);
  nand (_29269_, _15259_, _05732_);
  and (_29270_, _29269_, _06306_);
  and (_29272_, _29270_, _29268_);
  or (_29273_, _29063_, _12723_);
  or (_29274_, _12027_, _12722_);
  and (_29275_, _29274_, _06129_);
  and (_29276_, _29275_, _29273_);
  or (_29277_, _29276_, _12541_);
  or (_29278_, _29277_, _29272_);
  and (_29279_, _29278_, _29043_);
  or (_29280_, _29279_, _10976_);
  or (_29281_, _11880_, _10975_);
  and (_29283_, _29281_, _11016_);
  and (_29284_, _29283_, _29280_);
  and (_29285_, _29042_, _11015_);
  or (_29286_, _29285_, _06049_);
  or (_29287_, _29286_, _29284_);
  nand (_29288_, _07977_, _06049_);
  and (_29289_, _29288_, _29287_);
  or (_29290_, _29289_, _05747_);
  nand (_29291_, _15259_, _05747_);
  and (_29292_, _29291_, _06704_);
  and (_29294_, _29292_, _29290_);
  or (_29295_, _29063_, _12722_);
  nand (_29296_, _12028_, _12722_);
  and (_29297_, _29296_, _29295_);
  and (_29298_, _29297_, _06126_);
  or (_29299_, _29298_, _12750_);
  or (_29300_, _29299_, _29294_);
  or (_29301_, _29042_, _12749_);
  and (_29302_, _29301_, _06718_);
  and (_29303_, _29302_, _29300_);
  nand (_29305_, _11880_, _06316_);
  nand (_29306_, _29305_, _12756_);
  or (_29307_, _29306_, _29303_);
  or (_29308_, _29042_, _12756_);
  and (_29309_, _29308_, _09200_);
  and (_29310_, _29309_, _29307_);
  nor (_29311_, _06359_, _09200_);
  or (_29312_, _29311_, _05752_);
  or (_29313_, _29312_, _29310_);
  nand (_29314_, _15259_, _05752_);
  and (_29316_, _29314_, _05653_);
  and (_29317_, _29316_, _29313_);
  and (_29318_, _29297_, _05652_);
  or (_29319_, _29318_, _12772_);
  or (_29320_, _29319_, _29317_);
  or (_29321_, _29042_, _12771_);
  and (_29322_, _29321_, _06048_);
  and (_29323_, _29322_, _29320_);
  nand (_29324_, _11880_, _06047_);
  nand (_29325_, _29324_, _12779_);
  or (_29327_, _29325_, _29323_);
  or (_29328_, _29042_, _12779_);
  and (_29329_, _29328_, _12782_);
  and (_29330_, _29329_, _29327_);
  nor (_29331_, _06359_, _12782_);
  or (_29332_, _29331_, _05751_);
  or (_29333_, _29332_, _29330_);
  nand (_29334_, _15259_, _05751_);
  and (_29335_, _29334_, _12790_);
  and (_29336_, _29335_, _29333_);
  and (_29338_, _29042_, _12789_);
  or (_29339_, _29338_, _29336_);
  or (_29340_, _29339_, _01340_);
  or (_29341_, _01336_, \oc8051_golden_model_1.PC [13]);
  and (_29342_, _29341_, _42882_);
  and (_43431_, _29342_, _29340_);
  and (_29343_, _15457_, _06047_);
  nor (_29344_, _29039_, \oc8051_golden_model_1.PC [14]);
  nor (_29345_, _29344_, _11868_);
  not (_29346_, _29345_);
  nand (_29348_, _29346_, _11015_);
  nor (_29349_, _12515_, _15457_);
  nor (_29350_, _12494_, _15457_);
  nor (_29351_, _12473_, _15457_);
  or (_29352_, _29345_, _12231_);
  and (_29353_, _29345_, _06948_);
  and (_29354_, _12197_, _11875_);
  nor (_29355_, _11972_, _11878_);
  nor (_29356_, _29355_, _11973_);
  and (_29357_, _29356_, _12199_);
  or (_29359_, _29357_, _29354_);
  or (_29360_, _29359_, _08383_);
  or (_29361_, _29345_, _12205_);
  nand (_29362_, _12205_, _15457_);
  and (_29363_, _29362_, _29361_);
  or (_29364_, _29363_, _24785_);
  nor (_29365_, _29346_, _12215_);
  nand (_29366_, _15457_, _06938_);
  and (_29367_, _29366_, _25758_);
  and (_29368_, _07251_, \oc8051_golden_model_1.PC [14]);
  or (_29370_, _29368_, _06938_);
  and (_29371_, _29370_, _29367_);
  or (_29372_, _29371_, _06943_);
  or (_29373_, _29372_, _29365_);
  and (_29374_, _29373_, _29364_);
  or (_29375_, _29374_, _08384_);
  and (_29376_, _29375_, _06949_);
  and (_29377_, _29376_, _29360_);
  or (_29378_, _29377_, _29353_);
  or (_29379_, _29378_, _06102_);
  or (_29381_, _12187_, _12020_);
  and (_29382_, _12133_, _12025_);
  nor (_29383_, _29382_, _12134_);
  or (_29384_, _29383_, _12189_);
  and (_29385_, _29384_, _29381_);
  or (_29386_, _29385_, _06954_);
  and (_29387_, _29386_, _29379_);
  or (_29388_, _29387_, _24805_);
  or (_29389_, _29345_, _12182_);
  and (_29390_, _29389_, _12179_);
  and (_29392_, _29390_, _29388_);
  nor (_29393_, _12179_, _15457_);
  or (_29394_, _29393_, _12232_);
  or (_29395_, _29394_, _29392_);
  and (_29396_, _29395_, _29352_);
  or (_29397_, _29396_, _06219_);
  nand (_29398_, _15457_, _06219_);
  and (_29399_, _29398_, _12239_);
  and (_29400_, _29399_, _29397_);
  nor (_29401_, _29346_, _12239_);
  or (_29403_, _29401_, _29400_);
  and (_29404_, _29403_, _12245_);
  or (_29405_, _12245_, _15457_);
  nand (_29406_, _29405_, _12255_);
  or (_29407_, _29406_, _29404_);
  and (_29408_, _12289_, _12020_);
  not (_29409_, _29383_);
  nor (_29410_, _29409_, _12289_);
  or (_29411_, _29410_, _29408_);
  or (_29412_, _29411_, _12255_);
  and (_29414_, _29412_, _12258_);
  and (_29415_, _29414_, _29407_);
  nand (_29416_, _29409_, _12174_);
  or (_29417_, _12174_, _12020_);
  and (_29418_, _29417_, _06104_);
  and (_29419_, _29418_, _29416_);
  or (_29420_, _29419_, _06121_);
  or (_29421_, _29420_, _29415_);
  and (_29422_, _12310_, _12020_);
  nor (_29423_, _29409_, _12310_);
  or (_29425_, _29423_, _06509_);
  or (_29426_, _29425_, _29422_);
  and (_29427_, _29426_, _12298_);
  and (_29428_, _29427_, _29421_);
  or (_29429_, _29383_, _12329_);
  nand (_29430_, _12329_, _12021_);
  and (_29431_, _29430_, _06115_);
  and (_29432_, _29431_, _29429_);
  or (_29433_, _29432_, _12012_);
  or (_29434_, _29433_, _29428_);
  or (_29436_, _29345_, _12013_);
  and (_29437_, _29436_, _12345_);
  and (_29438_, _29437_, _29434_);
  nor (_29439_, _12345_, _15457_);
  or (_29440_, _29439_, _12355_);
  or (_29441_, _29440_, _29438_);
  or (_29442_, _29345_, _12351_);
  and (_29443_, _29442_, _12357_);
  and (_29444_, _29443_, _29441_);
  nor (_29445_, _12357_, _15457_);
  or (_29447_, _29445_, _12368_);
  or (_29448_, _29447_, _29444_);
  or (_29449_, _29345_, _12362_);
  and (_29450_, _29449_, _12366_);
  and (_29451_, _29450_, _29448_);
  nor (_29452_, _15457_, _12366_);
  or (_29453_, _29452_, _05676_);
  or (_29454_, _29453_, _29451_);
  or (_29455_, _29345_, _05675_);
  and (_29456_, _29455_, _12376_);
  and (_29458_, _29456_, _29454_);
  nor (_29459_, _12376_, _15457_);
  or (_29460_, _29459_, _06110_);
  or (_29461_, _29460_, _29458_);
  nand (_29462_, _12021_, _06110_);
  and (_29463_, _29462_, _09817_);
  and (_29464_, _29463_, _29461_);
  nor (_29465_, _15457_, _09817_);
  or (_29466_, _29465_, _09833_);
  or (_29467_, _29466_, _29464_);
  or (_29469_, _12020_, _05669_);
  and (_29470_, _29469_, _12389_);
  and (_29471_, _29470_, _29467_);
  nor (_29472_, _29346_, _12389_);
  or (_29473_, _29472_, _12392_);
  or (_29474_, _29473_, _29471_);
  or (_29475_, _12391_, _11875_);
  and (_29476_, _29475_, _12398_);
  and (_29477_, _29476_, _29474_);
  and (_29478_, _29356_, _12397_);
  or (_29480_, _29478_, _08743_);
  or (_29481_, _29480_, _29477_);
  or (_29482_, _11875_, _08742_);
  and (_29483_, _29482_, _29481_);
  or (_29484_, _29483_, _06019_);
  nand (_29485_, _12021_, _06019_);
  and (_29486_, _29485_, _10662_);
  and (_29487_, _29486_, _29484_);
  and (_29488_, _11875_, _10661_);
  or (_29489_, _29488_, _12412_);
  or (_29491_, _29489_, _29487_);
  nor (_29492_, _12445_, \oc8051_golden_model_1.DPH [6]);
  nor (_29493_, _29492_, _12446_);
  or (_29494_, _29493_, _12413_);
  and (_29495_, _29494_, _12415_);
  and (_29496_, _29495_, _29491_);
  nor (_29497_, _12415_, _15457_);
  or (_29498_, _29497_, _29496_);
  and (_29499_, _29498_, _12454_);
  or (_29500_, _29356_, _11071_);
  or (_29502_, _11875_, _12459_);
  and (_29503_, _29502_, _12453_);
  and (_29504_, _29503_, _29500_);
  or (_29505_, _29504_, _12006_);
  or (_29506_, _29505_, _29499_);
  nand (_29507_, _29346_, _12006_);
  and (_29508_, _29507_, _12466_);
  and (_29509_, _29508_, _29506_);
  nor (_29510_, _12466_, _15457_);
  or (_29511_, _29510_, _06112_);
  or (_29513_, _29511_, _29509_);
  nand (_29514_, _12021_, _06112_);
  and (_29515_, _29514_, _12473_);
  and (_29516_, _29515_, _29513_);
  or (_29517_, _29516_, _29351_);
  and (_29518_, _29517_, _12477_);
  or (_29519_, _29356_, _12459_);
  or (_29520_, _11875_, _11071_);
  and (_29521_, _29520_, _12476_);
  and (_29522_, _29521_, _29519_);
  or (_29523_, _29522_, _12481_);
  or (_29524_, _29523_, _29518_);
  or (_29525_, _29345_, _12002_);
  and (_29526_, _29525_, _10742_);
  and (_29527_, _29526_, _29524_);
  nor (_29528_, _15457_, _10742_);
  or (_29529_, _29528_, _06108_);
  or (_29530_, _29529_, _29527_);
  nand (_29531_, _12021_, _06108_);
  and (_29532_, _29531_, _12494_);
  and (_29535_, _29532_, _29530_);
  or (_29536_, _29535_, _29350_);
  and (_29537_, _29536_, _12498_);
  or (_29538_, _29356_, \oc8051_golden_model_1.PSW [7]);
  or (_29539_, _11875_, _10606_);
  and (_29540_, _29539_, _12497_);
  and (_29541_, _29540_, _29538_);
  or (_29542_, _29541_, _12502_);
  or (_29543_, _29542_, _29537_);
  or (_29544_, _29345_, _11993_);
  and (_29546_, _29544_, _11986_);
  and (_29547_, _29546_, _29543_);
  nor (_29548_, _15457_, _11986_);
  or (_29549_, _29548_, _06130_);
  or (_29550_, _29549_, _29547_);
  nand (_29551_, _12021_, _06130_);
  and (_29552_, _29551_, _12515_);
  and (_29553_, _29552_, _29550_);
  or (_29554_, _29553_, _29349_);
  and (_29555_, _29554_, _12518_);
  or (_29557_, _29356_, _10606_);
  or (_29558_, _11875_, \oc8051_golden_model_1.PSW [7]);
  and (_29559_, _29558_, _11982_);
  and (_29560_, _29559_, _29557_);
  or (_29561_, _29560_, _12525_);
  or (_29562_, _29561_, _29555_);
  or (_29563_, _29345_, _12523_);
  and (_29564_, _29563_, _10825_);
  and (_29565_, _29564_, _29562_);
  nor (_29566_, _15457_, _10825_);
  or (_29568_, _29566_, _10854_);
  or (_29569_, _29568_, _29565_);
  nand (_29570_, _29346_, _10854_);
  and (_29571_, _29570_, _13619_);
  and (_29572_, _29571_, _29569_);
  nor (_29573_, _07883_, _13619_);
  or (_29574_, _29573_, _05732_);
  or (_29575_, _29574_, _29572_);
  nand (_29576_, _15457_, _05732_);
  and (_29577_, _29576_, _06306_);
  and (_29579_, _29577_, _29575_);
  or (_29580_, _12020_, _12722_);
  nand (_29581_, _29409_, _12722_);
  and (_29582_, _29581_, _06129_);
  and (_29583_, _29582_, _29580_);
  or (_29584_, _29583_, _12541_);
  or (_29585_, _29584_, _29579_);
  or (_29586_, _29345_, _11872_);
  and (_29587_, _29586_, _10975_);
  and (_29588_, _29587_, _29585_);
  nor (_29590_, _15457_, _10975_);
  or (_29591_, _29590_, _11015_);
  or (_29592_, _29591_, _29588_);
  and (_29593_, _29592_, _29348_);
  or (_29594_, _29593_, _06049_);
  nand (_29595_, _07883_, _06049_);
  and (_29596_, _29595_, _05748_);
  and (_29597_, _29596_, _29594_);
  and (_29598_, _11875_, _05747_);
  or (_29599_, _29598_, _06126_);
  or (_29601_, _29599_, _29597_);
  and (_29602_, _12021_, _12722_);
  nor (_29603_, _29383_, _12722_);
  nor (_29604_, _29603_, _29602_);
  or (_29605_, _29604_, _06704_);
  and (_29606_, _29605_, _29601_);
  nor (_29607_, _29606_, _12750_);
  nor (_29608_, _29345_, _12749_);
  nor (_29609_, _29608_, _29607_);
  nor (_29610_, _29609_, _06316_);
  nand (_29612_, _15457_, _06316_);
  and (_29613_, _29612_, _12756_);
  not (_29614_, _29613_);
  nor (_29615_, _29614_, _29610_);
  nor (_29616_, _29346_, _12756_);
  nor (_29617_, _29616_, _06127_);
  not (_29618_, _29617_);
  nor (_29619_, _29618_, _29615_);
  and (_29620_, _06127_, _06084_);
  or (_29621_, _29620_, _05752_);
  nor (_29623_, _29621_, _29619_);
  and (_29624_, _11875_, _05752_);
  or (_29625_, _29624_, _05652_);
  nor (_29626_, _29625_, _29623_);
  nor (_29627_, _29604_, _05653_);
  nor (_29628_, _29627_, _12772_);
  not (_29629_, _29628_);
  nor (_29630_, _29629_, _29626_);
  nor (_29631_, _29346_, _12771_);
  nor (_29632_, _29631_, _06047_);
  not (_29634_, _29632_);
  nor (_29635_, _29634_, _29630_);
  or (_29636_, _29635_, _26405_);
  nor (_29637_, _29636_, _29343_);
  nor (_29638_, _29346_, _12779_);
  or (_29639_, _29638_, _29637_);
  and (_29640_, _29639_, _12782_);
  nor (_29641_, _12782_, _06084_);
  or (_29642_, _29641_, _29640_);
  and (_29643_, _29642_, _12791_);
  and (_29645_, _11875_, _05751_);
  or (_29646_, _29645_, _29643_);
  and (_29647_, _29646_, _12790_);
  and (_29648_, _29345_, _12789_);
  or (_29649_, _29648_, _29647_);
  or (_29650_, _29649_, _01340_);
  or (_29651_, _01336_, \oc8051_golden_model_1.PC [14]);
  and (_29652_, _29651_, _42882_);
  and (_43432_, _29652_, _29650_);
  nor (_29653_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_29655_, _29653_, _00000_);
  and (_29656_, _12800_, \oc8051_golden_model_1.P2 [0]);
  and (_29657_, _07686_, _08672_);
  or (_29658_, _29657_, _29656_);
  or (_29659_, _29658_, _06020_);
  and (_29660_, _09120_, _07686_);
  or (_29661_, _29656_, _07012_);
  or (_29662_, _29661_, _29660_);
  nor (_29663_, _08127_, _12800_);
  or (_29664_, _29663_, _29656_);
  or (_29666_, _29664_, _06954_);
  and (_29667_, _07686_, \oc8051_golden_model_1.ACC [0]);
  or (_29668_, _29667_, _29656_);
  and (_29669_, _29668_, _06938_);
  and (_29670_, _06939_, \oc8051_golden_model_1.P2 [0]);
  or (_29671_, _29670_, _06102_);
  or (_29672_, _29671_, _29669_);
  and (_29673_, _29672_, _06044_);
  and (_29674_, _29673_, _29666_);
  and (_29675_, _12819_, \oc8051_golden_model_1.P2 [0]);
  and (_29677_, _14102_, _08349_);
  or (_29678_, _29677_, _29675_);
  and (_29679_, _29678_, _06043_);
  or (_29680_, _29679_, _29674_);
  and (_29681_, _29680_, _06848_);
  and (_29682_, _07686_, _06931_);
  or (_29683_, _29682_, _29656_);
  and (_29684_, _29683_, _06239_);
  or (_29685_, _29684_, _06219_);
  or (_29686_, _29685_, _29681_);
  or (_29688_, _29668_, _06220_);
  and (_29689_, _29688_, _06040_);
  and (_29690_, _29689_, _29686_);
  and (_29691_, _29656_, _06039_);
  or (_29692_, _29691_, _06032_);
  or (_29693_, _29692_, _29690_);
  or (_29694_, _29664_, _06033_);
  and (_29695_, _29694_, _06027_);
  and (_29696_, _29695_, _29693_);
  or (_29697_, _29675_, _14131_);
  and (_29699_, _29697_, _06026_);
  and (_29700_, _29699_, _29678_);
  or (_29701_, _29700_, _09818_);
  or (_29702_, _29701_, _29696_);
  or (_29703_, _29683_, _09827_);
  and (_29704_, _29703_, _05669_);
  and (_29705_, _29704_, _29702_);
  and (_29706_, _29705_, _29662_);
  and (_29707_, _14186_, _07686_);
  or (_29708_, _29707_, _29656_);
  and (_29710_, _29708_, _09833_);
  or (_29711_, _29710_, _06019_);
  or (_29712_, _29711_, _29706_);
  and (_29713_, _29712_, _29659_);
  or (_29714_, _29713_, _06112_);
  and (_29715_, _14086_, _07686_);
  or (_29716_, _29656_, _08751_);
  or (_29717_, _29716_, _29715_);
  and (_29718_, _29717_, _08756_);
  and (_29719_, _29718_, _29714_);
  nor (_29721_, _12302_, _12800_);
  or (_29722_, _29721_, _29656_);
  nand (_29723_, _10995_, _07686_);
  and (_29724_, _29723_, _06284_);
  and (_29725_, _29724_, _29722_);
  or (_29726_, _29725_, _29719_);
  and (_29727_, _29726_, _07032_);
  nand (_29728_, _29658_, _06108_);
  nor (_29729_, _29728_, _29663_);
  or (_29730_, _29729_, _06277_);
  or (_29732_, _29730_, _29727_);
  nor (_29733_, _29656_, _06278_);
  nand (_29734_, _29733_, _29723_);
  and (_29735_, _29734_, _29732_);
  or (_29736_, _29735_, _06130_);
  and (_29737_, _14083_, _07686_);
  or (_29738_, _29656_, _08777_);
  or (_29739_, _29738_, _29737_);
  and (_29740_, _29739_, _08782_);
  and (_29741_, _29740_, _29736_);
  and (_29743_, _29722_, _06292_);
  or (_29744_, _29743_, _06316_);
  or (_29745_, _29744_, _29741_);
  or (_29746_, _29664_, _06718_);
  and (_29747_, _29746_, _29745_);
  or (_29748_, _29747_, _05652_);
  or (_29749_, _29656_, _05653_);
  and (_29750_, _29749_, _29748_);
  or (_29751_, _29750_, _06047_);
  or (_29752_, _29664_, _06048_);
  and (_29754_, _29752_, _01336_);
  and (_29755_, _29754_, _29751_);
  or (_43434_, _29755_, _29655_);
  nor (_29756_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_29757_, _29756_, _00000_);
  and (_29758_, _12800_, \oc8051_golden_model_1.P2 [1]);
  nor (_29759_, _10993_, _12800_);
  or (_29760_, _29759_, _29758_);
  or (_29761_, _29760_, _08782_);
  nor (_29762_, _12800_, _07132_);
  or (_29764_, _29762_, _29758_);
  or (_29765_, _29764_, _06848_);
  or (_29766_, _07686_, \oc8051_golden_model_1.P2 [1]);
  and (_29767_, _14284_, _07686_);
  not (_29768_, _29767_);
  and (_29769_, _29768_, _29766_);
  or (_29770_, _29769_, _06954_);
  and (_29771_, _07686_, \oc8051_golden_model_1.ACC [1]);
  or (_29772_, _29771_, _29758_);
  and (_29773_, _29772_, _06938_);
  and (_29775_, _06939_, \oc8051_golden_model_1.P2 [1]);
  or (_29776_, _29775_, _06102_);
  or (_29777_, _29776_, _29773_);
  and (_29778_, _29777_, _06044_);
  and (_29779_, _29778_, _29770_);
  and (_29780_, _12819_, \oc8051_golden_model_1.P2 [1]);
  and (_29781_, _14266_, _08349_);
  or (_29782_, _29781_, _29780_);
  and (_29783_, _29782_, _06043_);
  or (_29784_, _29783_, _06239_);
  or (_29786_, _29784_, _29779_);
  and (_29787_, _29786_, _29765_);
  or (_29788_, _29787_, _06219_);
  or (_29789_, _29772_, _06220_);
  and (_29790_, _29789_, _06040_);
  and (_29791_, _29790_, _29788_);
  and (_29792_, _14273_, _08349_);
  or (_29793_, _29792_, _29780_);
  and (_29794_, _29793_, _06039_);
  or (_29795_, _29794_, _06032_);
  or (_29796_, _29795_, _29791_);
  and (_29797_, _29781_, _14302_);
  or (_29798_, _29780_, _06033_);
  or (_29799_, _29798_, _29797_);
  and (_29800_, _29799_, _06027_);
  and (_29801_, _29800_, _29796_);
  or (_29802_, _29780_, _14267_);
  and (_29803_, _29802_, _06026_);
  and (_29804_, _29803_, _29782_);
  or (_29805_, _29804_, _09818_);
  or (_29808_, _29805_, _29801_);
  and (_29809_, _09075_, _07686_);
  or (_29810_, _29758_, _07012_);
  or (_29811_, _29810_, _29809_);
  or (_29812_, _29764_, _09827_);
  and (_29813_, _29812_, _05669_);
  and (_29814_, _29813_, _29811_);
  and (_29815_, _29814_, _29808_);
  and (_29816_, _14367_, _07686_);
  or (_29817_, _29816_, _29758_);
  and (_29819_, _29817_, _09833_);
  or (_29820_, _29819_, _29815_);
  and (_29821_, _29820_, _06020_);
  nand (_29822_, _07686_, _06832_);
  and (_29823_, _29766_, _06019_);
  and (_29824_, _29823_, _29822_);
  or (_29825_, _29824_, _29821_);
  and (_29826_, _29825_, _08751_);
  or (_29827_, _14263_, _12800_);
  and (_29828_, _29766_, _06112_);
  and (_29830_, _29828_, _29827_);
  or (_29831_, _29830_, _06284_);
  or (_29832_, _29831_, _29826_);
  nand (_29833_, _10992_, _07686_);
  and (_29834_, _29833_, _29760_);
  or (_29835_, _29834_, _08756_);
  and (_29836_, _29835_, _07032_);
  and (_29837_, _29836_, _29832_);
  or (_29838_, _14261_, _12800_);
  and (_29839_, _29766_, _06108_);
  and (_29841_, _29839_, _29838_);
  or (_29842_, _29841_, _06277_);
  or (_29843_, _29842_, _29837_);
  nor (_29844_, _29758_, _06278_);
  nand (_29845_, _29844_, _29833_);
  and (_29846_, _29845_, _08777_);
  and (_29847_, _29846_, _29843_);
  or (_29848_, _29822_, _08078_);
  and (_29849_, _29766_, _06130_);
  and (_29850_, _29849_, _29848_);
  or (_29852_, _29850_, _06292_);
  or (_29853_, _29852_, _29847_);
  and (_29854_, _29853_, _29761_);
  or (_29855_, _29854_, _06316_);
  or (_29856_, _29769_, _06718_);
  and (_29857_, _29856_, _05653_);
  and (_29858_, _29857_, _29855_);
  and (_29859_, _29793_, _05652_);
  or (_29860_, _29859_, _06047_);
  or (_29861_, _29860_, _29858_);
  or (_29863_, _29758_, _06048_);
  or (_29864_, _29863_, _29767_);
  and (_29865_, _29864_, _01336_);
  and (_29866_, _29865_, _29861_);
  or (_43435_, _29866_, _29757_);
  nor (_29867_, \oc8051_golden_model_1.P2 [2], rst);
  nor (_29868_, _29867_, _00000_);
  and (_29869_, _12800_, \oc8051_golden_model_1.P2 [2]);
  or (_29870_, _29869_, _08177_);
  and (_29871_, _07686_, _08730_);
  or (_29873_, _29871_, _29869_);
  and (_29874_, _29873_, _06108_);
  and (_29875_, _29874_, _29870_);
  or (_29876_, _29873_, _06020_);
  nor (_29877_, _12800_, _07530_);
  or (_29878_, _29877_, _29869_);
  or (_29879_, _29878_, _06848_);
  and (_29880_, _14493_, _07686_);
  or (_29881_, _29880_, _29869_);
  or (_29882_, _29881_, _06954_);
  and (_29884_, _07686_, \oc8051_golden_model_1.ACC [2]);
  or (_29885_, _29884_, _29869_);
  and (_29886_, _29885_, _06938_);
  and (_29887_, _06939_, \oc8051_golden_model_1.P2 [2]);
  or (_29888_, _29887_, _06102_);
  or (_29889_, _29888_, _29886_);
  and (_29890_, _29889_, _06044_);
  and (_29891_, _29890_, _29882_);
  and (_29892_, _12819_, \oc8051_golden_model_1.P2 [2]);
  and (_29893_, _14497_, _08349_);
  or (_29895_, _29893_, _29892_);
  and (_29896_, _29895_, _06043_);
  or (_29897_, _29896_, _06239_);
  or (_29898_, _29897_, _29891_);
  and (_29899_, _29898_, _29879_);
  or (_29900_, _29899_, _06219_);
  or (_29901_, _29885_, _06220_);
  and (_29902_, _29901_, _06040_);
  and (_29903_, _29902_, _29900_);
  and (_29904_, _14479_, _08349_);
  or (_29906_, _29904_, _29892_);
  and (_29907_, _29906_, _06039_);
  or (_29908_, _29907_, _06032_);
  or (_29909_, _29908_, _29903_);
  and (_29910_, _29893_, _14512_);
  or (_29911_, _29892_, _06033_);
  or (_29912_, _29911_, _29910_);
  and (_29913_, _29912_, _06027_);
  and (_29914_, _29913_, _29909_);
  or (_29915_, _29892_, _14525_);
  and (_29917_, _29915_, _06026_);
  and (_29918_, _29917_, _29895_);
  or (_29919_, _29918_, _09818_);
  or (_29920_, _29919_, _29914_);
  and (_29921_, _09182_, _07686_);
  or (_29922_, _29869_, _07012_);
  or (_29923_, _29922_, _29921_);
  or (_29924_, _29878_, _09827_);
  and (_29925_, _29924_, _05669_);
  and (_29926_, _29925_, _29923_);
  and (_29928_, _29926_, _29920_);
  and (_29929_, _14580_, _07686_);
  or (_29930_, _29929_, _29869_);
  and (_29931_, _29930_, _09833_);
  or (_29932_, _29931_, _06019_);
  or (_29933_, _29932_, _29928_);
  and (_29934_, _29933_, _29876_);
  or (_29935_, _29934_, _06112_);
  and (_29936_, _14596_, _07686_);
  or (_29937_, _29936_, _29869_);
  or (_29939_, _29937_, _08751_);
  and (_29940_, _29939_, _08756_);
  and (_29941_, _29940_, _29935_);
  and (_29942_, _10991_, _07686_);
  or (_29943_, _29942_, _29869_);
  and (_29944_, _29943_, _06284_);
  or (_29945_, _29944_, _29941_);
  and (_29946_, _29945_, _07032_);
  or (_29947_, _29946_, _29875_);
  and (_29948_, _29947_, _06278_);
  and (_29950_, _29885_, _06277_);
  and (_29951_, _29950_, _29870_);
  or (_29952_, _29951_, _06130_);
  or (_29953_, _29952_, _29948_);
  and (_29954_, _14593_, _07686_);
  or (_29955_, _29869_, _08777_);
  or (_29956_, _29955_, _29954_);
  and (_29957_, _29956_, _08782_);
  and (_29958_, _29957_, _29953_);
  nor (_29959_, _10990_, _12800_);
  or (_29961_, _29959_, _29869_);
  and (_29962_, _29961_, _06292_);
  or (_29963_, _29962_, _06316_);
  or (_29964_, _29963_, _29958_);
  or (_29965_, _29881_, _06718_);
  and (_29966_, _29965_, _05653_);
  and (_29967_, _29966_, _29964_);
  and (_29968_, _29906_, _05652_);
  or (_29969_, _29968_, _06047_);
  or (_29970_, _29969_, _29967_);
  and (_29972_, _14657_, _07686_);
  or (_29973_, _29869_, _06048_);
  or (_29974_, _29973_, _29972_);
  and (_29975_, _29974_, _01336_);
  and (_29976_, _29975_, _29970_);
  or (_43436_, _29976_, _29868_);
  and (_29977_, _12800_, \oc8051_golden_model_1.P2 [3]);
  and (_29978_, _07686_, _08662_);
  or (_29979_, _29978_, _29977_);
  or (_29980_, _29979_, _06020_);
  and (_29982_, _14672_, _07686_);
  or (_29983_, _29982_, _29977_);
  or (_29984_, _29983_, _06954_);
  and (_29985_, _07686_, \oc8051_golden_model_1.ACC [3]);
  or (_29986_, _29985_, _29977_);
  and (_29987_, _29986_, _06938_);
  and (_29988_, _06939_, \oc8051_golden_model_1.P2 [3]);
  or (_29989_, _29988_, _06102_);
  or (_29990_, _29989_, _29987_);
  and (_29991_, _29990_, _06044_);
  and (_29993_, _29991_, _29984_);
  and (_29994_, _12819_, \oc8051_golden_model_1.P2 [3]);
  and (_29995_, _14683_, _08349_);
  or (_29996_, _29995_, _29994_);
  and (_29997_, _29996_, _06043_);
  or (_29998_, _29997_, _06239_);
  or (_29999_, _29998_, _29993_);
  nor (_30000_, _12800_, _07353_);
  or (_30001_, _30000_, _29977_);
  or (_30002_, _30001_, _06848_);
  and (_30004_, _30002_, _29999_);
  or (_30005_, _30004_, _06219_);
  or (_30006_, _29986_, _06220_);
  and (_30007_, _30006_, _06040_);
  and (_30008_, _30007_, _30005_);
  and (_30009_, _14681_, _08349_);
  or (_30010_, _30009_, _29994_);
  and (_30011_, _30010_, _06039_);
  or (_30012_, _30011_, _06032_);
  or (_30013_, _30012_, _30008_);
  or (_30015_, _29994_, _14708_);
  and (_30016_, _30015_, _29996_);
  or (_30017_, _30016_, _06033_);
  and (_30018_, _30017_, _06027_);
  and (_30019_, _30018_, _30013_);
  and (_30020_, _14724_, _08349_);
  or (_30021_, _30020_, _29994_);
  and (_30022_, _30021_, _06026_);
  or (_30023_, _30022_, _09818_);
  or (_30024_, _30023_, _30019_);
  and (_30026_, _09181_, _07686_);
  or (_30027_, _29977_, _07012_);
  or (_30028_, _30027_, _30026_);
  or (_30029_, _30001_, _09827_);
  and (_30030_, _30029_, _05669_);
  and (_30031_, _30030_, _30028_);
  and (_30032_, _30031_, _30024_);
  and (_30033_, _14778_, _07686_);
  or (_30034_, _30033_, _29977_);
  and (_30035_, _30034_, _09833_);
  or (_30037_, _30035_, _06019_);
  or (_30038_, _30037_, _30032_);
  and (_30039_, _30038_, _29980_);
  or (_30040_, _30039_, _06112_);
  and (_30041_, _14793_, _07686_);
  or (_30042_, _29977_, _08751_);
  or (_30043_, _30042_, _30041_);
  and (_30044_, _30043_, _08756_);
  and (_30045_, _30044_, _30040_);
  and (_30046_, _12299_, _07686_);
  or (_30048_, _30046_, _29977_);
  and (_30049_, _30048_, _06284_);
  or (_30050_, _30049_, _30045_);
  and (_30051_, _30050_, _07032_);
  or (_30052_, _29977_, _08029_);
  and (_30053_, _29979_, _06108_);
  and (_30054_, _30053_, _30052_);
  or (_30055_, _30054_, _30051_);
  and (_30056_, _30055_, _06278_);
  and (_30057_, _29986_, _06277_);
  and (_30059_, _30057_, _30052_);
  or (_30060_, _30059_, _06130_);
  or (_30061_, _30060_, _30056_);
  and (_30062_, _14792_, _07686_);
  or (_30063_, _29977_, _08777_);
  or (_30064_, _30063_, _30062_);
  and (_30065_, _30064_, _08782_);
  and (_30066_, _30065_, _30061_);
  nor (_30067_, _10988_, _12800_);
  or (_30068_, _30067_, _29977_);
  and (_30070_, _30068_, _06292_);
  or (_30071_, _30070_, _06316_);
  or (_30072_, _30071_, _30066_);
  or (_30073_, _29983_, _06718_);
  and (_30074_, _30073_, _05653_);
  and (_30075_, _30074_, _30072_);
  and (_30076_, _30010_, _05652_);
  or (_30077_, _30076_, _06047_);
  or (_30078_, _30077_, _30075_);
  and (_30079_, _14849_, _07686_);
  or (_30081_, _29977_, _06048_);
  or (_30082_, _30081_, _30079_);
  and (_30083_, _30082_, _01336_);
  and (_30084_, _30083_, _30078_);
  nor (_30085_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_30086_, _30085_, _00000_);
  or (_43437_, _30086_, _30084_);
  and (_30087_, _12800_, \oc8051_golden_model_1.P2 [4]);
  and (_30088_, _08665_, _07686_);
  or (_30089_, _30088_, _30087_);
  or (_30091_, _30089_, _06020_);
  and (_30092_, _14887_, _07686_);
  or (_30093_, _30092_, _30087_);
  or (_30094_, _30093_, _06954_);
  and (_30095_, _07686_, \oc8051_golden_model_1.ACC [4]);
  or (_30096_, _30095_, _30087_);
  and (_30097_, _30096_, _06938_);
  and (_30098_, _06939_, \oc8051_golden_model_1.P2 [4]);
  or (_30099_, _30098_, _06102_);
  or (_30100_, _30099_, _30097_);
  and (_30102_, _30100_, _06044_);
  and (_30103_, _30102_, _30094_);
  and (_30104_, _12819_, \oc8051_golden_model_1.P2 [4]);
  and (_30105_, _14878_, _08349_);
  or (_30106_, _30105_, _30104_);
  and (_30107_, _30106_, _06043_);
  or (_30108_, _30107_, _06239_);
  or (_30109_, _30108_, _30103_);
  nor (_30110_, _08270_, _12800_);
  or (_30111_, _30110_, _30087_);
  or (_30113_, _30111_, _06848_);
  and (_30114_, _30113_, _30109_);
  or (_30115_, _30114_, _06219_);
  or (_30116_, _30096_, _06220_);
  and (_30117_, _30116_, _06040_);
  and (_30118_, _30117_, _30115_);
  and (_30119_, _14882_, _08349_);
  or (_30120_, _30119_, _30104_);
  and (_30121_, _30120_, _06039_);
  or (_30122_, _30121_, _06032_);
  or (_30124_, _30122_, _30118_);
  or (_30125_, _30104_, _14914_);
  and (_30126_, _30125_, _30106_);
  or (_30127_, _30126_, _06033_);
  and (_30128_, _30127_, _06027_);
  and (_30129_, _30128_, _30124_);
  or (_30130_, _30104_, _14879_);
  and (_30131_, _30130_, _06026_);
  and (_30132_, _30131_, _30106_);
  or (_30133_, _30132_, _09818_);
  or (_30135_, _30133_, _30129_);
  and (_30136_, _09180_, _07686_);
  or (_30137_, _30087_, _07012_);
  or (_30138_, _30137_, _30136_);
  or (_30139_, _30111_, _09827_);
  and (_30140_, _30139_, _05669_);
  and (_30141_, _30140_, _30138_);
  and (_30142_, _30141_, _30135_);
  and (_30143_, _14983_, _07686_);
  or (_30144_, _30143_, _30087_);
  and (_30146_, _30144_, _09833_);
  or (_30147_, _30146_, _06019_);
  or (_30148_, _30147_, _30142_);
  and (_30149_, _30148_, _30091_);
  or (_30150_, _30149_, _06112_);
  and (_30151_, _14876_, _07686_);
  or (_30152_, _30087_, _08751_);
  or (_30153_, _30152_, _30151_);
  and (_30154_, _30153_, _08756_);
  and (_30155_, _30154_, _30150_);
  and (_30157_, _10986_, _07686_);
  or (_30158_, _30157_, _30087_);
  and (_30159_, _30158_, _06284_);
  or (_30160_, _30159_, _30155_);
  and (_30161_, _30160_, _07032_);
  or (_30162_, _30087_, _08273_);
  and (_30163_, _30089_, _06108_);
  and (_30164_, _30163_, _30162_);
  or (_30165_, _30164_, _30161_);
  and (_30166_, _30165_, _06278_);
  and (_30168_, _30096_, _06277_);
  and (_30169_, _30168_, _30162_);
  or (_30170_, _30169_, _06130_);
  or (_30171_, _30170_, _30166_);
  and (_30172_, _14873_, _07686_);
  or (_30173_, _30087_, _08777_);
  or (_30174_, _30173_, _30172_);
  and (_30175_, _30174_, _08782_);
  and (_30176_, _30175_, _30171_);
  nor (_30177_, _10985_, _12800_);
  or (_30179_, _30177_, _30087_);
  and (_30180_, _30179_, _06292_);
  or (_30181_, _30180_, _06316_);
  or (_30182_, _30181_, _30176_);
  or (_30183_, _30093_, _06718_);
  and (_30184_, _30183_, _05653_);
  and (_30185_, _30184_, _30182_);
  and (_30186_, _30120_, _05652_);
  or (_30187_, _30186_, _06047_);
  or (_30188_, _30187_, _30185_);
  and (_30190_, _15055_, _07686_);
  or (_30191_, _30087_, _06048_);
  or (_30192_, _30191_, _30190_);
  and (_30193_, _30192_, _01336_);
  and (_30194_, _30193_, _30188_);
  nor (_30195_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_30196_, _30195_, _00000_);
  or (_43438_, _30196_, _30194_);
  and (_30197_, _12800_, \oc8051_golden_model_1.P2 [5]);
  and (_30198_, _08652_, _07686_);
  or (_30200_, _30198_, _30197_);
  or (_30201_, _30200_, _06020_);
  and (_30202_, _15093_, _07686_);
  or (_30203_, _30202_, _30197_);
  or (_30204_, _30203_, _06954_);
  and (_30205_, _07686_, \oc8051_golden_model_1.ACC [5]);
  or (_30206_, _30205_, _30197_);
  and (_30207_, _30206_, _06938_);
  and (_30208_, _06939_, \oc8051_golden_model_1.P2 [5]);
  or (_30209_, _30208_, _06102_);
  or (_30211_, _30209_, _30207_);
  and (_30212_, _30211_, _06044_);
  and (_30213_, _30212_, _30204_);
  and (_30214_, _12819_, \oc8051_golden_model_1.P2 [5]);
  and (_30215_, _15073_, _08349_);
  or (_30216_, _30215_, _30214_);
  and (_30217_, _30216_, _06043_);
  or (_30218_, _30217_, _06239_);
  or (_30219_, _30218_, _30213_);
  nor (_30220_, _07977_, _12800_);
  or (_30222_, _30220_, _30197_);
  or (_30223_, _30222_, _06848_);
  and (_30224_, _30223_, _30219_);
  or (_30225_, _30224_, _06219_);
  or (_30226_, _30206_, _06220_);
  and (_30227_, _30226_, _06040_);
  and (_30228_, _30227_, _30225_);
  and (_30229_, _15077_, _08349_);
  or (_30230_, _30229_, _30214_);
  and (_30231_, _30230_, _06039_);
  or (_30233_, _30231_, _06032_);
  or (_30234_, _30233_, _30228_);
  or (_30235_, _30214_, _15110_);
  and (_30236_, _30235_, _30216_);
  or (_30237_, _30236_, _06033_);
  and (_30238_, _30237_, _06027_);
  and (_30239_, _30238_, _30234_);
  or (_30240_, _30214_, _15074_);
  and (_30241_, _30240_, _06026_);
  and (_30242_, _30241_, _30216_);
  or (_30244_, _30242_, _09818_);
  or (_30245_, _30244_, _30239_);
  and (_30246_, _09179_, _07686_);
  or (_30247_, _30197_, _07012_);
  or (_30248_, _30247_, _30246_);
  or (_30249_, _30222_, _09827_);
  and (_30250_, _30249_, _05669_);
  and (_30251_, _30250_, _30248_);
  and (_30252_, _30251_, _30245_);
  and (_30253_, _15179_, _07686_);
  or (_30255_, _30253_, _30197_);
  and (_30256_, _30255_, _09833_);
  or (_30257_, _30256_, _06019_);
  or (_30258_, _30257_, _30252_);
  and (_30259_, _30258_, _30201_);
  or (_30260_, _30259_, _06112_);
  and (_30261_, _15195_, _07686_);
  or (_30262_, _30197_, _08751_);
  or (_30263_, _30262_, _30261_);
  and (_30264_, _30263_, _08756_);
  and (_30266_, _30264_, _30260_);
  and (_30267_, _12306_, _07686_);
  or (_30268_, _30267_, _30197_);
  and (_30269_, _30268_, _06284_);
  or (_30270_, _30269_, _30266_);
  and (_30271_, _30270_, _07032_);
  or (_30272_, _30197_, _07980_);
  and (_30273_, _30200_, _06108_);
  and (_30274_, _30273_, _30272_);
  or (_30275_, _30274_, _30271_);
  and (_30277_, _30275_, _06278_);
  and (_30278_, _30206_, _06277_);
  and (_30279_, _30278_, _30272_);
  or (_30280_, _30279_, _06130_);
  or (_30281_, _30280_, _30277_);
  and (_30282_, _15194_, _07686_);
  or (_30283_, _30197_, _08777_);
  or (_30284_, _30283_, _30282_);
  and (_30285_, _30284_, _08782_);
  and (_30286_, _30285_, _30281_);
  nor (_30288_, _10982_, _12800_);
  or (_30289_, _30288_, _30197_);
  and (_30290_, _30289_, _06292_);
  or (_30291_, _30290_, _06316_);
  or (_30292_, _30291_, _30286_);
  or (_30293_, _30203_, _06718_);
  and (_30294_, _30293_, _05653_);
  and (_30295_, _30294_, _30292_);
  and (_30296_, _30230_, _05652_);
  or (_30297_, _30296_, _06047_);
  or (_30299_, _30297_, _30295_);
  and (_30300_, _15253_, _07686_);
  or (_30301_, _30197_, _06048_);
  or (_30302_, _30301_, _30300_);
  and (_30303_, _30302_, _01336_);
  and (_30304_, _30303_, _30299_);
  nor (_30305_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_30306_, _30305_, _00000_);
  or (_43440_, _30306_, _30304_);
  nor (_30307_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_30309_, _30307_, _00000_);
  and (_30310_, _12800_, \oc8051_golden_model_1.P2 [6]);
  and (_30311_, _15389_, _07686_);
  or (_30312_, _30311_, _30310_);
  or (_30313_, _30312_, _06020_);
  and (_30314_, _15293_, _07686_);
  or (_30315_, _30314_, _30310_);
  or (_30316_, _30315_, _06954_);
  and (_30317_, _07686_, \oc8051_golden_model_1.ACC [6]);
  or (_30318_, _30317_, _30310_);
  and (_30320_, _30318_, _06938_);
  and (_30321_, _06939_, \oc8051_golden_model_1.P2 [6]);
  or (_30322_, _30321_, _06102_);
  or (_30323_, _30322_, _30320_);
  and (_30324_, _30323_, _06044_);
  and (_30325_, _30324_, _30316_);
  and (_30326_, _12819_, \oc8051_golden_model_1.P2 [6]);
  and (_30327_, _15280_, _08349_);
  or (_30328_, _30327_, _30326_);
  and (_30329_, _30328_, _06043_);
  or (_30331_, _30329_, _06239_);
  or (_30332_, _30331_, _30325_);
  nor (_30333_, _07883_, _12800_);
  or (_30334_, _30333_, _30310_);
  or (_30335_, _30334_, _06848_);
  and (_30336_, _30335_, _30332_);
  or (_30337_, _30336_, _06219_);
  or (_30338_, _30318_, _06220_);
  and (_30339_, _30338_, _06040_);
  and (_30340_, _30339_, _30337_);
  and (_30342_, _15278_, _08349_);
  or (_30343_, _30342_, _30326_);
  and (_30344_, _30343_, _06039_);
  or (_30345_, _30344_, _06032_);
  or (_30346_, _30345_, _30340_);
  or (_30347_, _30326_, _15310_);
  and (_30348_, _30347_, _30328_);
  or (_30349_, _30348_, _06033_);
  and (_30350_, _30349_, _06027_);
  and (_30351_, _30350_, _30346_);
  or (_30353_, _30326_, _15326_);
  and (_30354_, _30353_, _06026_);
  and (_30355_, _30354_, _30328_);
  or (_30356_, _30355_, _09818_);
  or (_30357_, _30356_, _30351_);
  and (_30358_, _09178_, _07686_);
  or (_30359_, _30310_, _07012_);
  or (_30360_, _30359_, _30358_);
  or (_30361_, _30334_, _09827_);
  and (_30362_, _30361_, _05669_);
  and (_30364_, _30362_, _30360_);
  and (_30365_, _30364_, _30357_);
  and (_30366_, _15382_, _07686_);
  or (_30367_, _30366_, _30310_);
  and (_30368_, _30367_, _09833_);
  or (_30369_, _30368_, _06019_);
  or (_30370_, _30369_, _30365_);
  and (_30371_, _30370_, _30313_);
  or (_30372_, _30371_, _06112_);
  and (_30373_, _15399_, _07686_);
  or (_30375_, _30373_, _30310_);
  or (_30376_, _30375_, _08751_);
  and (_30377_, _30376_, _08756_);
  and (_30378_, _30377_, _30372_);
  and (_30379_, _10980_, _07686_);
  or (_30380_, _30379_, _30310_);
  and (_30381_, _30380_, _06284_);
  or (_30382_, _30381_, _30378_);
  and (_30383_, _30382_, _07032_);
  or (_30384_, _30310_, _07886_);
  and (_30386_, _30312_, _06108_);
  and (_30387_, _30386_, _30384_);
  or (_30388_, _30387_, _30383_);
  and (_30389_, _30388_, _06278_);
  and (_30390_, _30318_, _06277_);
  and (_30391_, _30390_, _30384_);
  or (_30392_, _30391_, _06130_);
  or (_30393_, _30392_, _30389_);
  and (_30394_, _15396_, _07686_);
  or (_30395_, _30310_, _08777_);
  or (_30397_, _30395_, _30394_);
  and (_30398_, _30397_, _08782_);
  and (_30399_, _30398_, _30393_);
  nor (_30400_, _10979_, _12800_);
  or (_30401_, _30400_, _30310_);
  and (_30402_, _30401_, _06292_);
  or (_30403_, _30402_, _06316_);
  or (_30404_, _30403_, _30399_);
  or (_30405_, _30315_, _06718_);
  and (_30406_, _30405_, _05653_);
  and (_30408_, _30406_, _30404_);
  and (_30409_, _30343_, _05652_);
  or (_30410_, _30409_, _06047_);
  or (_30411_, _30410_, _30408_);
  and (_30412_, _15451_, _07686_);
  or (_30413_, _30310_, _06048_);
  or (_30414_, _30413_, _30412_);
  and (_30415_, _30414_, _01336_);
  and (_30416_, _30415_, _30411_);
  or (_43441_, _30416_, _30309_);
  nand (_30417_, _10995_, _07692_);
  and (_30418_, _12902_, \oc8051_golden_model_1.P3 [0]);
  nor (_30419_, _30418_, _06278_);
  nand (_30420_, _30419_, _30417_);
  and (_30421_, _07692_, _08672_);
  or (_30422_, _30421_, _30418_);
  or (_30423_, _30422_, _06020_);
  and (_30424_, _09120_, _07692_);
  or (_30425_, _30418_, _07012_);
  or (_30426_, _30425_, _30424_);
  nor (_30429_, _08127_, _12902_);
  or (_30430_, _30429_, _30418_);
  or (_30431_, _30430_, _06954_);
  and (_30432_, _07692_, \oc8051_golden_model_1.ACC [0]);
  or (_30433_, _30432_, _30418_);
  and (_30434_, _30433_, _06938_);
  and (_30435_, _06939_, \oc8051_golden_model_1.P3 [0]);
  or (_30436_, _30435_, _06102_);
  or (_30437_, _30436_, _30434_);
  and (_30438_, _30437_, _06044_);
  and (_30440_, _30438_, _30431_);
  and (_30441_, _12921_, \oc8051_golden_model_1.P3 [0]);
  and (_30442_, _14102_, _08353_);
  or (_30443_, _30442_, _30441_);
  and (_30444_, _30443_, _06043_);
  or (_30445_, _30444_, _30440_);
  and (_30446_, _30445_, _06848_);
  and (_30447_, _07692_, _06931_);
  or (_30448_, _30447_, _30418_);
  and (_30449_, _30448_, _06239_);
  or (_30451_, _30449_, _06219_);
  or (_30452_, _30451_, _30446_);
  or (_30453_, _30433_, _06220_);
  and (_30454_, _30453_, _06040_);
  and (_30455_, _30454_, _30452_);
  and (_30456_, _30418_, _06039_);
  or (_30457_, _30456_, _06032_);
  or (_30458_, _30457_, _30455_);
  or (_30459_, _30430_, _06033_);
  and (_30460_, _30459_, _06027_);
  and (_30462_, _30460_, _30458_);
  or (_30463_, _30441_, _14131_);
  and (_30464_, _30463_, _06026_);
  and (_30465_, _30464_, _30443_);
  or (_30466_, _30465_, _09818_);
  or (_30467_, _30466_, _30462_);
  or (_30468_, _30448_, _09827_);
  and (_30469_, _30468_, _05669_);
  and (_30470_, _30469_, _30467_);
  and (_30471_, _30470_, _30426_);
  and (_30473_, _14186_, _07692_);
  or (_30474_, _30473_, _30418_);
  and (_30475_, _30474_, _09833_);
  or (_30476_, _30475_, _06019_);
  or (_30477_, _30476_, _30471_);
  and (_30478_, _30477_, _30423_);
  or (_30479_, _30478_, _06112_);
  and (_30480_, _14086_, _07692_);
  or (_30481_, _30418_, _08751_);
  or (_30482_, _30481_, _30480_);
  and (_30484_, _30482_, _08756_);
  and (_30485_, _30484_, _30479_);
  nor (_30486_, _12302_, _12902_);
  or (_30487_, _30486_, _30418_);
  and (_30488_, _30417_, _06284_);
  and (_30489_, _30488_, _30487_);
  or (_30490_, _30489_, _30485_);
  and (_30491_, _30490_, _07032_);
  nand (_30492_, _30422_, _06108_);
  nor (_30493_, _30492_, _30429_);
  or (_30495_, _30493_, _06277_);
  or (_30496_, _30495_, _30491_);
  and (_30497_, _30496_, _30420_);
  or (_30498_, _30497_, _06130_);
  and (_30499_, _14083_, _07692_);
  or (_30500_, _30418_, _08777_);
  or (_30501_, _30500_, _30499_);
  and (_30502_, _30501_, _08782_);
  and (_30503_, _30502_, _30498_);
  and (_30504_, _30487_, _06292_);
  or (_30506_, _30504_, _06316_);
  or (_30507_, _30506_, _30503_);
  or (_30508_, _30430_, _06718_);
  and (_30509_, _30508_, _30507_);
  or (_30510_, _30509_, _05652_);
  or (_30511_, _30418_, _05653_);
  and (_30512_, _30511_, _30510_);
  or (_30513_, _30512_, _06047_);
  or (_30514_, _30430_, _06048_);
  and (_30515_, _30514_, _01336_);
  and (_30517_, _30515_, _30513_);
  nor (_30518_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_30519_, _30518_, _00000_);
  or (_43442_, _30519_, _30517_);
  and (_30520_, _12902_, \oc8051_golden_model_1.P3 [1]);
  nor (_30521_, _10993_, _12902_);
  or (_30522_, _30521_, _30520_);
  or (_30523_, _30522_, _08782_);
  nor (_30524_, _12902_, _07132_);
  or (_30525_, _30524_, _30520_);
  or (_30527_, _30525_, _06848_);
  or (_30528_, _07692_, \oc8051_golden_model_1.P3 [1]);
  and (_30529_, _14284_, _07692_);
  not (_30530_, _30529_);
  and (_30531_, _30530_, _30528_);
  or (_30532_, _30531_, _06954_);
  and (_30533_, _07692_, \oc8051_golden_model_1.ACC [1]);
  or (_30534_, _30533_, _30520_);
  and (_30535_, _30534_, _06938_);
  and (_30536_, _06939_, \oc8051_golden_model_1.P3 [1]);
  or (_30538_, _30536_, _06102_);
  or (_30539_, _30538_, _30535_);
  and (_30540_, _30539_, _06044_);
  and (_30541_, _30540_, _30532_);
  and (_30542_, _12921_, \oc8051_golden_model_1.P3 [1]);
  and (_30543_, _14266_, _08353_);
  or (_30544_, _30543_, _30542_);
  and (_30545_, _30544_, _06043_);
  or (_30546_, _30545_, _06239_);
  or (_30547_, _30546_, _30541_);
  and (_30549_, _30547_, _30527_);
  or (_30550_, _30549_, _06219_);
  or (_30551_, _30534_, _06220_);
  and (_30552_, _30551_, _06040_);
  and (_30553_, _30552_, _30550_);
  and (_30554_, _14273_, _08353_);
  or (_30555_, _30554_, _30542_);
  and (_30556_, _30555_, _06039_);
  or (_30557_, _30556_, _06032_);
  or (_30558_, _30557_, _30553_);
  and (_30560_, _30543_, _14302_);
  or (_30561_, _30542_, _06033_);
  or (_30562_, _30561_, _30560_);
  and (_30563_, _30562_, _06027_);
  and (_30564_, _30563_, _30558_);
  or (_30565_, _30542_, _14267_);
  and (_30566_, _30565_, _06026_);
  and (_30567_, _30566_, _30544_);
  or (_30568_, _30567_, _09818_);
  or (_30569_, _30568_, _30564_);
  and (_30571_, _09075_, _07692_);
  or (_30572_, _30520_, _07012_);
  or (_30573_, _30572_, _30571_);
  or (_30574_, _30525_, _09827_);
  and (_30575_, _30574_, _05669_);
  and (_30576_, _30575_, _30573_);
  and (_30577_, _30576_, _30569_);
  and (_30578_, _14367_, _07692_);
  or (_30579_, _30578_, _30520_);
  and (_30580_, _30579_, _09833_);
  or (_30582_, _30580_, _30577_);
  and (_30583_, _30582_, _06020_);
  nand (_30584_, _07692_, _06832_);
  and (_30585_, _30528_, _06019_);
  and (_30586_, _30585_, _30584_);
  or (_30587_, _30586_, _30583_);
  and (_30588_, _30587_, _08751_);
  or (_30589_, _14263_, _12902_);
  and (_30590_, _30528_, _06112_);
  and (_30591_, _30590_, _30589_);
  or (_30593_, _30591_, _06284_);
  or (_30594_, _30593_, _30588_);
  nand (_30595_, _10992_, _07692_);
  and (_30596_, _30595_, _30522_);
  or (_30597_, _30596_, _08756_);
  and (_30598_, _30597_, _07032_);
  and (_30599_, _30598_, _30594_);
  or (_30600_, _14261_, _12902_);
  and (_30601_, _30528_, _06108_);
  and (_30602_, _30601_, _30600_);
  or (_30604_, _30602_, _06277_);
  or (_30605_, _30604_, _30599_);
  nor (_30606_, _30520_, _06278_);
  nand (_30607_, _30606_, _30595_);
  and (_30608_, _30607_, _08777_);
  and (_30609_, _30608_, _30605_);
  or (_30610_, _30584_, _08078_);
  and (_30611_, _30528_, _06130_);
  and (_30612_, _30611_, _30610_);
  or (_30613_, _30612_, _06292_);
  or (_30615_, _30613_, _30609_);
  and (_30616_, _30615_, _30523_);
  or (_30617_, _30616_, _06316_);
  or (_30618_, _30531_, _06718_);
  and (_30619_, _30618_, _05653_);
  and (_30620_, _30619_, _30617_);
  and (_30621_, _30555_, _05652_);
  or (_30622_, _30621_, _06047_);
  or (_30623_, _30622_, _30620_);
  or (_30624_, _30520_, _06048_);
  or (_30626_, _30624_, _30529_);
  and (_30627_, _30626_, _01336_);
  and (_30628_, _30627_, _30623_);
  nor (_30629_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_30630_, _30629_, _00000_);
  or (_43444_, _30630_, _30628_);
  nor (_30631_, \oc8051_golden_model_1.P3 [2], rst);
  nor (_30632_, _30631_, _00000_);
  and (_30633_, _12902_, \oc8051_golden_model_1.P3 [2]);
  and (_30634_, _07692_, _08730_);
  or (_30636_, _30634_, _30633_);
  or (_30637_, _30636_, _06020_);
  nor (_30638_, _12902_, _07530_);
  or (_30639_, _30638_, _30633_);
  and (_30640_, _30639_, _06239_);
  and (_30641_, _12921_, \oc8051_golden_model_1.P3 [2]);
  and (_30642_, _14497_, _08353_);
  or (_30643_, _30642_, _30641_);
  or (_30644_, _30643_, _06044_);
  and (_30645_, _14493_, _07692_);
  or (_30647_, _30645_, _30633_);
  and (_30648_, _30647_, _06102_);
  and (_30649_, _06939_, \oc8051_golden_model_1.P3 [2]);
  and (_30650_, _07692_, \oc8051_golden_model_1.ACC [2]);
  or (_30651_, _30650_, _30633_);
  and (_30652_, _30651_, _06938_);
  or (_30653_, _30652_, _30649_);
  and (_30654_, _30653_, _06954_);
  or (_30655_, _30654_, _06043_);
  or (_30656_, _30655_, _30648_);
  and (_30658_, _30656_, _30644_);
  and (_30659_, _30658_, _06848_);
  or (_30660_, _30659_, _30640_);
  or (_30661_, _30660_, _06219_);
  or (_30662_, _30651_, _06220_);
  and (_30663_, _30662_, _06040_);
  and (_30664_, _30663_, _30661_);
  and (_30665_, _14479_, _08353_);
  or (_30666_, _30665_, _30641_);
  and (_30667_, _30666_, _06039_);
  or (_30669_, _30667_, _06032_);
  or (_30670_, _30669_, _30664_);
  or (_30671_, _30641_, _14512_);
  and (_30672_, _30671_, _30643_);
  or (_30673_, _30672_, _06033_);
  and (_30674_, _30673_, _06027_);
  and (_30675_, _30674_, _30670_);
  or (_30676_, _30641_, _14525_);
  and (_30677_, _30676_, _06026_);
  and (_30678_, _30677_, _30643_);
  or (_30680_, _30678_, _09818_);
  or (_30681_, _30680_, _30675_);
  and (_30682_, _09182_, _07692_);
  or (_30683_, _30633_, _07012_);
  or (_30684_, _30683_, _30682_);
  or (_30685_, _30639_, _09827_);
  and (_30686_, _30685_, _05669_);
  and (_30687_, _30686_, _30684_);
  and (_30688_, _30687_, _30681_);
  and (_30689_, _14580_, _07692_);
  or (_30691_, _30689_, _30633_);
  and (_30692_, _30691_, _09833_);
  or (_30693_, _30692_, _06019_);
  or (_30694_, _30693_, _30688_);
  and (_30695_, _30694_, _30637_);
  or (_30696_, _30695_, _06112_);
  and (_30697_, _14596_, _07692_);
  or (_30698_, _30633_, _08751_);
  or (_30699_, _30698_, _30697_);
  and (_30700_, _30699_, _08756_);
  and (_30702_, _30700_, _30696_);
  and (_30703_, _10991_, _07692_);
  or (_30704_, _30703_, _30633_);
  and (_30705_, _30704_, _06284_);
  or (_30706_, _30705_, _30702_);
  and (_30707_, _30706_, _07032_);
  or (_30708_, _30633_, _08177_);
  and (_30709_, _30636_, _06108_);
  and (_30710_, _30709_, _30708_);
  or (_30711_, _30710_, _30707_);
  and (_30713_, _30711_, _06278_);
  and (_30714_, _30651_, _06277_);
  and (_30715_, _30714_, _30708_);
  or (_30716_, _30715_, _06130_);
  or (_30717_, _30716_, _30713_);
  and (_30718_, _14593_, _07692_);
  or (_30719_, _30633_, _08777_);
  or (_30720_, _30719_, _30718_);
  and (_30721_, _30720_, _08782_);
  and (_30722_, _30721_, _30717_);
  nor (_30724_, _10990_, _12902_);
  or (_30725_, _30724_, _30633_);
  and (_30726_, _30725_, _06292_);
  or (_30727_, _30726_, _06316_);
  or (_30728_, _30727_, _30722_);
  or (_30729_, _30647_, _06718_);
  and (_30730_, _30729_, _05653_);
  and (_30731_, _30730_, _30728_);
  and (_30732_, _30666_, _05652_);
  or (_30733_, _30732_, _06047_);
  or (_30735_, _30733_, _30731_);
  and (_30736_, _14657_, _07692_);
  or (_30737_, _30633_, _06048_);
  or (_30738_, _30737_, _30736_);
  and (_30739_, _30738_, _01336_);
  and (_30740_, _30739_, _30735_);
  or (_43445_, _30740_, _30632_);
  nor (_30741_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_30742_, _30741_, _00000_);
  and (_30743_, _12902_, \oc8051_golden_model_1.P3 [3]);
  and (_30745_, _07692_, _08662_);
  or (_30746_, _30745_, _30743_);
  or (_30747_, _30746_, _06020_);
  and (_30748_, _14672_, _07692_);
  or (_30749_, _30748_, _30743_);
  or (_30750_, _30749_, _06954_);
  and (_30751_, _07692_, \oc8051_golden_model_1.ACC [3]);
  or (_30752_, _30751_, _30743_);
  and (_30753_, _30752_, _06938_);
  and (_30754_, _06939_, \oc8051_golden_model_1.P3 [3]);
  or (_30756_, _30754_, _06102_);
  or (_30757_, _30756_, _30753_);
  and (_30758_, _30757_, _06044_);
  and (_30759_, _30758_, _30750_);
  and (_30760_, _12921_, \oc8051_golden_model_1.P3 [3]);
  and (_30761_, _14683_, _08353_);
  or (_30762_, _30761_, _30760_);
  and (_30763_, _30762_, _06043_);
  or (_30764_, _30763_, _06239_);
  or (_30765_, _30764_, _30759_);
  nor (_30767_, _12902_, _07353_);
  or (_30768_, _30767_, _30743_);
  or (_30769_, _30768_, _06848_);
  and (_30770_, _30769_, _30765_);
  or (_30771_, _30770_, _06219_);
  or (_30772_, _30752_, _06220_);
  and (_30773_, _30772_, _06040_);
  and (_30774_, _30773_, _30771_);
  and (_30775_, _14681_, _08353_);
  or (_30776_, _30775_, _30760_);
  and (_30778_, _30776_, _06039_);
  or (_30779_, _30778_, _06032_);
  or (_30780_, _30779_, _30774_);
  or (_30781_, _30760_, _14708_);
  and (_30782_, _30781_, _30762_);
  or (_30783_, _30782_, _06033_);
  and (_30784_, _30783_, _06027_);
  and (_30785_, _30784_, _30780_);
  and (_30786_, _14724_, _08353_);
  or (_30787_, _30786_, _30760_);
  and (_30789_, _30787_, _06026_);
  or (_30790_, _30789_, _09818_);
  or (_30791_, _30790_, _30785_);
  and (_30792_, _09181_, _07692_);
  or (_30793_, _30743_, _07012_);
  or (_30794_, _30793_, _30792_);
  or (_30795_, _30768_, _09827_);
  and (_30796_, _30795_, _05669_);
  and (_30797_, _30796_, _30794_);
  and (_30798_, _30797_, _30791_);
  and (_30800_, _14778_, _07692_);
  or (_30801_, _30800_, _30743_);
  and (_30802_, _30801_, _09833_);
  or (_30803_, _30802_, _06019_);
  or (_30804_, _30803_, _30798_);
  and (_30805_, _30804_, _30747_);
  or (_30806_, _30805_, _06112_);
  and (_30807_, _14793_, _07692_);
  or (_30808_, _30743_, _08751_);
  or (_30809_, _30808_, _30807_);
  and (_30811_, _30809_, _08756_);
  and (_30812_, _30811_, _30806_);
  and (_30813_, _12299_, _07692_);
  or (_30814_, _30813_, _30743_);
  and (_30815_, _30814_, _06284_);
  or (_30816_, _30815_, _30812_);
  and (_30817_, _30816_, _07032_);
  or (_30818_, _30743_, _08029_);
  and (_30819_, _30746_, _06108_);
  and (_30820_, _30819_, _30818_);
  or (_30822_, _30820_, _30817_);
  and (_30823_, _30822_, _06278_);
  and (_30824_, _30752_, _06277_);
  and (_30825_, _30824_, _30818_);
  or (_30826_, _30825_, _06130_);
  or (_30827_, _30826_, _30823_);
  and (_30828_, _14792_, _07692_);
  or (_30829_, _30743_, _08777_);
  or (_30830_, _30829_, _30828_);
  and (_30831_, _30830_, _08782_);
  and (_30833_, _30831_, _30827_);
  nor (_30834_, _10988_, _12902_);
  or (_30835_, _30834_, _30743_);
  and (_30836_, _30835_, _06292_);
  or (_30837_, _30836_, _06316_);
  or (_30838_, _30837_, _30833_);
  or (_30839_, _30749_, _06718_);
  and (_30840_, _30839_, _05653_);
  and (_30841_, _30840_, _30838_);
  and (_30842_, _30776_, _05652_);
  or (_30844_, _30842_, _06047_);
  or (_30845_, _30844_, _30841_);
  and (_30846_, _14849_, _07692_);
  or (_30847_, _30743_, _06048_);
  or (_30848_, _30847_, _30846_);
  and (_30849_, _30848_, _01336_);
  and (_30850_, _30849_, _30845_);
  or (_43446_, _30850_, _30742_);
  and (_30851_, _12902_, \oc8051_golden_model_1.P3 [4]);
  and (_30852_, _08665_, _07692_);
  or (_30854_, _30852_, _30851_);
  or (_30855_, _30854_, _06020_);
  and (_30856_, _14887_, _07692_);
  or (_30857_, _30856_, _30851_);
  or (_30858_, _30857_, _06954_);
  and (_30859_, _07692_, \oc8051_golden_model_1.ACC [4]);
  or (_30860_, _30859_, _30851_);
  and (_30861_, _30860_, _06938_);
  and (_30862_, _06939_, \oc8051_golden_model_1.P3 [4]);
  or (_30863_, _30862_, _06102_);
  or (_30865_, _30863_, _30861_);
  and (_30866_, _30865_, _06044_);
  and (_30867_, _30866_, _30858_);
  and (_30868_, _12921_, \oc8051_golden_model_1.P3 [4]);
  and (_30869_, _14878_, _08353_);
  or (_30870_, _30869_, _30868_);
  and (_30871_, _30870_, _06043_);
  or (_30872_, _30871_, _06239_);
  or (_30873_, _30872_, _30867_);
  nor (_30874_, _08270_, _12902_);
  or (_30876_, _30874_, _30851_);
  or (_30877_, _30876_, _06848_);
  and (_30878_, _30877_, _30873_);
  or (_30879_, _30878_, _06219_);
  or (_30880_, _30860_, _06220_);
  and (_30881_, _30880_, _06040_);
  and (_30882_, _30881_, _30879_);
  and (_30883_, _14882_, _08353_);
  or (_30884_, _30883_, _30868_);
  and (_30885_, _30884_, _06039_);
  or (_30887_, _30885_, _06032_);
  or (_30888_, _30887_, _30882_);
  or (_30889_, _30868_, _14914_);
  and (_30890_, _30889_, _30870_);
  or (_30891_, _30890_, _06033_);
  and (_30892_, _30891_, _06027_);
  and (_30893_, _30892_, _30888_);
  or (_30894_, _30868_, _14879_);
  and (_30895_, _30894_, _06026_);
  and (_30896_, _30895_, _30870_);
  or (_30898_, _30896_, _09818_);
  or (_30899_, _30898_, _30893_);
  and (_30900_, _09180_, _07692_);
  or (_30901_, _30851_, _07012_);
  or (_30902_, _30901_, _30900_);
  or (_30903_, _30876_, _09827_);
  and (_30904_, _30903_, _05669_);
  and (_30905_, _30904_, _30902_);
  and (_30906_, _30905_, _30899_);
  and (_30907_, _14983_, _07692_);
  or (_30909_, _30907_, _30851_);
  and (_30910_, _30909_, _09833_);
  or (_30911_, _30910_, _06019_);
  or (_30912_, _30911_, _30906_);
  and (_30913_, _30912_, _30855_);
  or (_30914_, _30913_, _06112_);
  and (_30915_, _14876_, _07692_);
  or (_30916_, _30915_, _30851_);
  or (_30917_, _30916_, _08751_);
  and (_30918_, _30917_, _08756_);
  and (_30920_, _30918_, _30914_);
  and (_30921_, _10986_, _07692_);
  or (_30922_, _30921_, _30851_);
  and (_30923_, _30922_, _06284_);
  or (_30924_, _30923_, _30920_);
  and (_30925_, _30924_, _07032_);
  or (_30926_, _30851_, _08273_);
  and (_30927_, _30854_, _06108_);
  and (_30928_, _30927_, _30926_);
  or (_30929_, _30928_, _30925_);
  and (_30931_, _30929_, _06278_);
  and (_30932_, _30860_, _06277_);
  and (_30933_, _30932_, _30926_);
  or (_30934_, _30933_, _06130_);
  or (_30935_, _30934_, _30931_);
  and (_30936_, _14873_, _07692_);
  or (_30937_, _30851_, _08777_);
  or (_30938_, _30937_, _30936_);
  and (_30939_, _30938_, _08782_);
  and (_30940_, _30939_, _30935_);
  nor (_30942_, _10985_, _12902_);
  or (_30943_, _30942_, _30851_);
  and (_30944_, _30943_, _06292_);
  or (_30945_, _30944_, _06316_);
  or (_30946_, _30945_, _30940_);
  or (_30947_, _30857_, _06718_);
  and (_30948_, _30947_, _05653_);
  and (_30949_, _30948_, _30946_);
  and (_30950_, _30884_, _05652_);
  or (_30951_, _30950_, _06047_);
  or (_30953_, _30951_, _30949_);
  and (_30954_, _15055_, _07692_);
  or (_30955_, _30851_, _06048_);
  or (_30956_, _30955_, _30954_);
  and (_30957_, _30956_, _01336_);
  and (_30958_, _30957_, _30953_);
  nor (_30959_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_30960_, _30959_, _00000_);
  or (_43447_, _30960_, _30958_);
  nor (_30961_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_30963_, _30961_, _00000_);
  and (_30964_, _12902_, \oc8051_golden_model_1.P3 [5]);
  and (_30965_, _08652_, _07692_);
  or (_30966_, _30965_, _30964_);
  or (_30967_, _30966_, _06020_);
  and (_30968_, _15093_, _07692_);
  or (_30969_, _30968_, _30964_);
  or (_30970_, _30969_, _06954_);
  and (_30971_, _07692_, \oc8051_golden_model_1.ACC [5]);
  or (_30972_, _30971_, _30964_);
  and (_30974_, _30972_, _06938_);
  and (_30975_, _06939_, \oc8051_golden_model_1.P3 [5]);
  or (_30976_, _30975_, _06102_);
  or (_30977_, _30976_, _30974_);
  and (_30978_, _30977_, _06044_);
  and (_30979_, _30978_, _30970_);
  and (_30980_, _12921_, \oc8051_golden_model_1.P3 [5]);
  and (_30981_, _15073_, _08353_);
  or (_30982_, _30981_, _30980_);
  and (_30983_, _30982_, _06043_);
  or (_30985_, _30983_, _06239_);
  or (_30986_, _30985_, _30979_);
  nor (_30987_, _07977_, _12902_);
  or (_30988_, _30987_, _30964_);
  or (_30989_, _30988_, _06848_);
  and (_30990_, _30989_, _30986_);
  or (_30991_, _30990_, _06219_);
  or (_30992_, _30972_, _06220_);
  and (_30993_, _30992_, _06040_);
  and (_30994_, _30993_, _30991_);
  and (_30996_, _15077_, _08353_);
  or (_30997_, _30996_, _30980_);
  and (_30998_, _30997_, _06039_);
  or (_30999_, _30998_, _06032_);
  or (_31000_, _30999_, _30994_);
  or (_31001_, _30980_, _15110_);
  and (_31002_, _31001_, _30982_);
  or (_31003_, _31002_, _06033_);
  and (_31004_, _31003_, _06027_);
  and (_31005_, _31004_, _31000_);
  or (_31007_, _30980_, _15074_);
  and (_31008_, _31007_, _06026_);
  and (_31009_, _31008_, _30982_);
  or (_31010_, _31009_, _09818_);
  or (_31011_, _31010_, _31005_);
  and (_31012_, _09179_, _07692_);
  or (_31013_, _30964_, _07012_);
  or (_31014_, _31013_, _31012_);
  or (_31015_, _30988_, _09827_);
  and (_31016_, _31015_, _05669_);
  and (_31018_, _31016_, _31014_);
  and (_31019_, _31018_, _31011_);
  and (_31020_, _15179_, _07692_);
  or (_31021_, _31020_, _30964_);
  and (_31022_, _31021_, _09833_);
  or (_31023_, _31022_, _06019_);
  or (_31024_, _31023_, _31019_);
  and (_31025_, _31024_, _30967_);
  or (_31026_, _31025_, _06112_);
  and (_31027_, _15195_, _07692_);
  or (_31029_, _30964_, _08751_);
  or (_31030_, _31029_, _31027_);
  and (_31031_, _31030_, _08756_);
  and (_31032_, _31031_, _31026_);
  and (_31033_, _12306_, _07692_);
  or (_31034_, _31033_, _30964_);
  and (_31035_, _31034_, _06284_);
  or (_31036_, _31035_, _31032_);
  and (_31037_, _31036_, _07032_);
  or (_31038_, _30964_, _07980_);
  and (_31040_, _30966_, _06108_);
  and (_31041_, _31040_, _31038_);
  or (_31042_, _31041_, _31037_);
  and (_31043_, _31042_, _06278_);
  and (_31044_, _30972_, _06277_);
  and (_31045_, _31044_, _31038_);
  or (_31046_, _31045_, _06130_);
  or (_31047_, _31046_, _31043_);
  and (_31048_, _15194_, _07692_);
  or (_31049_, _30964_, _08777_);
  or (_31051_, _31049_, _31048_);
  and (_31052_, _31051_, _08782_);
  and (_31053_, _31052_, _31047_);
  nor (_31054_, _10982_, _12902_);
  or (_31055_, _31054_, _30964_);
  and (_31056_, _31055_, _06292_);
  or (_31057_, _31056_, _06316_);
  or (_31058_, _31057_, _31053_);
  or (_31059_, _30969_, _06718_);
  and (_31060_, _31059_, _05653_);
  and (_31062_, _31060_, _31058_);
  and (_31063_, _30997_, _05652_);
  or (_31064_, _31063_, _06047_);
  or (_31065_, _31064_, _31062_);
  and (_31066_, _15253_, _07692_);
  or (_31067_, _30964_, _06048_);
  or (_31068_, _31067_, _31066_);
  and (_31069_, _31068_, _01336_);
  and (_31070_, _31069_, _31065_);
  or (_43448_, _31070_, _30963_);
  and (_31072_, _12902_, \oc8051_golden_model_1.P3 [6]);
  and (_31073_, _15389_, _07692_);
  or (_31074_, _31073_, _31072_);
  or (_31075_, _31074_, _06020_);
  and (_31076_, _15293_, _07692_);
  or (_31077_, _31076_, _31072_);
  or (_31078_, _31077_, _06954_);
  and (_31079_, _07692_, \oc8051_golden_model_1.ACC [6]);
  or (_31080_, _31079_, _31072_);
  and (_31081_, _31080_, _06938_);
  and (_31083_, _06939_, \oc8051_golden_model_1.P3 [6]);
  or (_31084_, _31083_, _06102_);
  or (_31085_, _31084_, _31081_);
  and (_31086_, _31085_, _06044_);
  and (_31087_, _31086_, _31078_);
  and (_31088_, _12921_, \oc8051_golden_model_1.P3 [6]);
  and (_31089_, _15280_, _08353_);
  or (_31090_, _31089_, _31088_);
  and (_31091_, _31090_, _06043_);
  or (_31092_, _31091_, _06239_);
  or (_31094_, _31092_, _31087_);
  nor (_31095_, _07883_, _12902_);
  or (_31096_, _31095_, _31072_);
  or (_31097_, _31096_, _06848_);
  and (_31098_, _31097_, _31094_);
  or (_31099_, _31098_, _06219_);
  or (_31100_, _31080_, _06220_);
  and (_31101_, _31100_, _06040_);
  and (_31102_, _31101_, _31099_);
  and (_31103_, _15278_, _08353_);
  or (_31105_, _31103_, _31088_);
  and (_31106_, _31105_, _06039_);
  or (_31107_, _31106_, _06032_);
  or (_31108_, _31107_, _31102_);
  or (_31109_, _31088_, _15310_);
  and (_31110_, _31109_, _31090_);
  or (_31111_, _31110_, _06033_);
  and (_31112_, _31111_, _06027_);
  and (_31113_, _31112_, _31108_);
  or (_31114_, _31088_, _15326_);
  and (_31116_, _31114_, _06026_);
  and (_31117_, _31116_, _31090_);
  or (_31118_, _31117_, _09818_);
  or (_31119_, _31118_, _31113_);
  and (_31120_, _09178_, _07692_);
  or (_31121_, _31072_, _07012_);
  or (_31122_, _31121_, _31120_);
  or (_31123_, _31096_, _09827_);
  and (_31124_, _31123_, _05669_);
  and (_31125_, _31124_, _31122_);
  and (_31127_, _31125_, _31119_);
  and (_31128_, _15382_, _07692_);
  or (_31129_, _31128_, _31072_);
  and (_31130_, _31129_, _09833_);
  or (_31131_, _31130_, _06019_);
  or (_31132_, _31131_, _31127_);
  and (_31133_, _31132_, _31075_);
  or (_31134_, _31133_, _06112_);
  and (_31135_, _15399_, _07692_);
  or (_31136_, _31072_, _08751_);
  or (_31139_, _31136_, _31135_);
  and (_31140_, _31139_, _08756_);
  and (_31141_, _31140_, _31134_);
  and (_31142_, _10980_, _07692_);
  or (_31143_, _31142_, _31072_);
  and (_31144_, _31143_, _06284_);
  or (_31145_, _31144_, _31141_);
  and (_31146_, _31145_, _07032_);
  or (_31147_, _31072_, _07886_);
  and (_31148_, _31074_, _06108_);
  and (_31150_, _31148_, _31147_);
  or (_31151_, _31150_, _31146_);
  and (_31152_, _31151_, _06278_);
  and (_31153_, _31080_, _06277_);
  and (_31154_, _31153_, _31147_);
  or (_31155_, _31154_, _06130_);
  or (_31156_, _31155_, _31152_);
  and (_31157_, _15396_, _07692_);
  or (_31158_, _31072_, _08777_);
  or (_31159_, _31158_, _31157_);
  and (_31162_, _31159_, _08782_);
  and (_31163_, _31162_, _31156_);
  nor (_31164_, _10979_, _12902_);
  or (_31165_, _31164_, _31072_);
  and (_31166_, _31165_, _06292_);
  or (_31167_, _31166_, _06316_);
  or (_31168_, _31167_, _31163_);
  or (_31169_, _31077_, _06718_);
  and (_31170_, _31169_, _05653_);
  and (_31171_, _31170_, _31168_);
  and (_31173_, _31105_, _05652_);
  or (_31174_, _31173_, _06047_);
  or (_31175_, _31174_, _31171_);
  and (_31176_, _15451_, _07692_);
  or (_31177_, _31072_, _06048_);
  or (_31178_, _31177_, _31176_);
  and (_31179_, _31178_, _01336_);
  and (_31180_, _31179_, _31175_);
  nor (_31181_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_31182_, _31181_, _00000_);
  or (_43449_, _31182_, _31180_);
  nor (_31185_, \oc8051_golden_model_1.P0 [0], rst);
  nor (_31186_, _31185_, _00000_);
  nand (_31187_, _10995_, _07730_);
  not (_31188_, \oc8051_golden_model_1.P0 [0]);
  nor (_31189_, _07730_, _31188_);
  nor (_31190_, _31189_, _06278_);
  nand (_31191_, _31190_, _31187_);
  and (_31192_, _07730_, _08672_);
  or (_31193_, _31192_, _31189_);
  or (_31195_, _31193_, _06020_);
  and (_31196_, _09120_, _07730_);
  or (_31197_, _31189_, _07012_);
  or (_31198_, _31197_, _31196_);
  nor (_31199_, _08127_, _13006_);
  or (_31200_, _31199_, _31189_);
  or (_31201_, _31200_, _06954_);
  and (_31202_, _07730_, \oc8051_golden_model_1.ACC [0]);
  or (_31203_, _31202_, _31189_);
  and (_31204_, _31203_, _06938_);
  nor (_31207_, _06938_, _31188_);
  or (_31208_, _31207_, _06102_);
  or (_31209_, _31208_, _31204_);
  and (_31210_, _31209_, _06044_);
  and (_31211_, _31210_, _31201_);
  nor (_31212_, _07638_, _31188_);
  and (_31213_, _14102_, _07638_);
  or (_31214_, _31213_, _31212_);
  and (_31215_, _31214_, _06043_);
  or (_31216_, _31215_, _31211_);
  and (_31218_, _31216_, _06848_);
  and (_31219_, _07730_, _06931_);
  or (_31220_, _31219_, _31189_);
  and (_31221_, _31220_, _06239_);
  or (_31222_, _31221_, _06219_);
  or (_31223_, _31222_, _31218_);
  or (_31224_, _31203_, _06220_);
  and (_31225_, _31224_, _06040_);
  and (_31226_, _31225_, _31223_);
  and (_31227_, _31189_, _06039_);
  or (_31229_, _31227_, _06032_);
  or (_31230_, _31229_, _31226_);
  or (_31231_, _31200_, _06033_);
  and (_31232_, _31231_, _06027_);
  and (_31233_, _31232_, _31230_);
  or (_31234_, _31212_, _14131_);
  and (_31235_, _31234_, _06026_);
  and (_31236_, _31235_, _31214_);
  or (_31237_, _31236_, _09818_);
  or (_31238_, _31237_, _31233_);
  or (_31240_, _31220_, _09827_);
  and (_31241_, _31240_, _05669_);
  and (_31242_, _31241_, _31238_);
  and (_31243_, _31242_, _31198_);
  and (_31244_, _14186_, _07730_);
  or (_31245_, _31244_, _31189_);
  and (_31246_, _31245_, _09833_);
  or (_31247_, _31246_, _06019_);
  or (_31248_, _31247_, _31243_);
  and (_31249_, _31248_, _31195_);
  or (_31250_, _31249_, _06112_);
  and (_31251_, _14086_, _07730_);
  or (_31252_, _31251_, _31189_);
  or (_31253_, _31252_, _08751_);
  and (_31254_, _31253_, _08756_);
  and (_31255_, _31254_, _31250_);
  nor (_31256_, _12302_, _13006_);
  or (_31257_, _31256_, _31189_);
  and (_31258_, _31187_, _06284_);
  and (_31259_, _31258_, _31257_);
  or (_31262_, _31259_, _31255_);
  and (_31263_, _31262_, _07032_);
  nand (_31264_, _31193_, _06108_);
  nor (_31265_, _31264_, _31199_);
  or (_31266_, _31265_, _06277_);
  or (_31267_, _31266_, _31263_);
  and (_31268_, _31267_, _31191_);
  or (_31269_, _31268_, _06130_);
  and (_31270_, _14083_, _07730_);
  or (_31271_, _31189_, _08777_);
  or (_31272_, _31271_, _31270_);
  and (_31273_, _31272_, _08782_);
  and (_31274_, _31273_, _31269_);
  and (_31275_, _31257_, _06292_);
  or (_31276_, _31275_, _06316_);
  or (_31277_, _31276_, _31274_);
  or (_31278_, _31200_, _06718_);
  and (_31279_, _31278_, _31277_);
  or (_31280_, _31279_, _05652_);
  or (_31281_, _31189_, _05653_);
  and (_31284_, _31281_, _31280_);
  or (_31285_, _31284_, _06047_);
  or (_31286_, _31200_, _06048_);
  and (_31287_, _31286_, _01336_);
  and (_31288_, _31287_, _31285_);
  or (_43451_, _31288_, _31186_);
  nor (_31289_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_31290_, _31289_, _00000_);
  and (_31291_, _13006_, \oc8051_golden_model_1.P0 [1]);
  nor (_31292_, _10993_, _13006_);
  or (_31293_, _31292_, _31291_);
  or (_31294_, _31293_, _08782_);
  or (_31295_, _14367_, _13006_);
  or (_31296_, _07730_, \oc8051_golden_model_1.P0 [1]);
  and (_31297_, _31296_, _09833_);
  and (_31298_, _31297_, _31295_);
  nor (_31299_, _13006_, _07132_);
  or (_31300_, _31299_, _31291_);
  or (_31301_, _31300_, _06848_);
  and (_31302_, _14284_, _07730_);
  not (_31305_, _31302_);
  and (_31306_, _31305_, _31296_);
  or (_31307_, _31306_, _06954_);
  and (_31308_, _07730_, \oc8051_golden_model_1.ACC [1]);
  or (_31309_, _31308_, _31291_);
  and (_31310_, _31309_, _06938_);
  and (_31311_, _06939_, \oc8051_golden_model_1.P0 [1]);
  or (_31312_, _31311_, _06102_);
  or (_31313_, _31312_, _31310_);
  and (_31314_, _31313_, _06044_);
  and (_31315_, _31314_, _31307_);
  and (_31316_, _13025_, \oc8051_golden_model_1.P0 [1]);
  and (_31317_, _14266_, _07638_);
  or (_31318_, _31317_, _31316_);
  and (_31319_, _31318_, _06043_);
  or (_31320_, _31319_, _06239_);
  or (_31321_, _31320_, _31315_);
  and (_31322_, _31321_, _31301_);
  or (_31323_, _31322_, _06219_);
  or (_31324_, _31309_, _06220_);
  and (_31327_, _31324_, _06040_);
  and (_31328_, _31327_, _31323_);
  and (_31329_, _14273_, _07638_);
  or (_31330_, _31329_, _31316_);
  and (_31331_, _31330_, _06039_);
  or (_31332_, _31331_, _06032_);
  or (_31333_, _31332_, _31328_);
  and (_31334_, _31317_, _14302_);
  or (_31335_, _31316_, _06033_);
  or (_31336_, _31335_, _31334_);
  and (_31337_, _31336_, _06027_);
  and (_31338_, _31337_, _31333_);
  or (_31339_, _31316_, _14267_);
  and (_31340_, _31339_, _06026_);
  and (_31341_, _31340_, _31318_);
  or (_31342_, _31341_, _09818_);
  or (_31343_, _31342_, _31338_);
  and (_31344_, _09075_, _07730_);
  or (_31345_, _31344_, _31291_);
  or (_31346_, _31345_, _07012_);
  or (_31349_, _31300_, _09827_);
  and (_31350_, _31349_, _05669_);
  and (_31351_, _31350_, _31346_);
  and (_31352_, _31351_, _31343_);
  or (_31353_, _31352_, _31298_);
  and (_31354_, _31353_, _06020_);
  nand (_31355_, _07730_, _06832_);
  and (_31356_, _31296_, _06019_);
  and (_31357_, _31356_, _31355_);
  or (_31358_, _31357_, _31354_);
  and (_31359_, _31358_, _08751_);
  or (_31360_, _14263_, _13006_);
  and (_31361_, _31296_, _06112_);
  and (_31362_, _31361_, _31360_);
  or (_31363_, _31362_, _06284_);
  or (_31364_, _31363_, _31359_);
  and (_31365_, _10994_, _07730_);
  or (_31366_, _31365_, _31291_);
  or (_31367_, _31366_, _08756_);
  and (_31368_, _31367_, _07032_);
  and (_31371_, _31368_, _31364_);
  or (_31372_, _14261_, _13006_);
  and (_31373_, _31296_, _06108_);
  and (_31374_, _31373_, _31372_);
  or (_31375_, _31374_, _06277_);
  or (_31376_, _31375_, _31371_);
  and (_31377_, _31308_, _08078_);
  or (_31378_, _31291_, _06278_);
  or (_31379_, _31378_, _31377_);
  and (_31380_, _31379_, _08777_);
  and (_31381_, _31380_, _31376_);
  or (_31382_, _31355_, _08078_);
  and (_31383_, _31296_, _06130_);
  and (_31384_, _31383_, _31382_);
  or (_31385_, _31384_, _06292_);
  or (_31386_, _31385_, _31381_);
  and (_31387_, _31386_, _31294_);
  or (_31388_, _31387_, _06316_);
  or (_31389_, _31306_, _06718_);
  and (_31390_, _31389_, _05653_);
  and (_31393_, _31390_, _31388_);
  and (_31394_, _31330_, _05652_);
  or (_31395_, _31394_, _06047_);
  or (_31396_, _31395_, _31393_);
  or (_31397_, _31291_, _06048_);
  or (_31398_, _31397_, _31302_);
  and (_31399_, _31398_, _01336_);
  and (_31400_, _31399_, _31396_);
  or (_43452_, _31400_, _31290_);
  nor (_31401_, \oc8051_golden_model_1.P0 [2], rst);
  nor (_31402_, _31401_, _00000_);
  and (_31403_, _13006_, \oc8051_golden_model_1.P0 [2]);
  or (_31404_, _31403_, _08177_);
  and (_31405_, _07730_, _08730_);
  or (_31406_, _31405_, _31403_);
  and (_31407_, _31406_, _06108_);
  and (_31408_, _31407_, _31404_);
  or (_31409_, _31406_, _06020_);
  nor (_31410_, _13006_, _07530_);
  or (_31411_, _31410_, _31403_);
  or (_31413_, _31411_, _06848_);
  and (_31414_, _14493_, _07730_);
  or (_31415_, _31414_, _31403_);
  or (_31416_, _31415_, _06954_);
  and (_31417_, _07730_, \oc8051_golden_model_1.ACC [2]);
  or (_31418_, _31417_, _31403_);
  and (_31419_, _31418_, _06938_);
  and (_31420_, _06939_, \oc8051_golden_model_1.P0 [2]);
  or (_31421_, _31420_, _06102_);
  or (_31422_, _31421_, _31419_);
  and (_31423_, _31422_, _06044_);
  and (_31424_, _31423_, _31416_);
  and (_31425_, _13025_, \oc8051_golden_model_1.P0 [2]);
  and (_31426_, _14497_, _07638_);
  or (_31427_, _31426_, _31425_);
  and (_31428_, _31427_, _06043_);
  or (_31429_, _31428_, _06239_);
  or (_31430_, _31429_, _31424_);
  and (_31431_, _31430_, _31413_);
  or (_31432_, _31431_, _06219_);
  or (_31435_, _31418_, _06220_);
  and (_31436_, _31435_, _06040_);
  and (_31437_, _31436_, _31432_);
  and (_31438_, _14479_, _07638_);
  or (_31439_, _31438_, _31425_);
  and (_31440_, _31439_, _06039_);
  or (_31441_, _31440_, _06032_);
  or (_31442_, _31441_, _31437_);
  and (_31443_, _31426_, _14512_);
  or (_31444_, _31425_, _06033_);
  or (_31445_, _31444_, _31443_);
  and (_31446_, _31445_, _06027_);
  and (_31447_, _31446_, _31442_);
  or (_31448_, _31425_, _14525_);
  and (_31449_, _31448_, _06026_);
  and (_31450_, _31449_, _31427_);
  or (_31451_, _31450_, _09818_);
  or (_31452_, _31451_, _31447_);
  and (_31453_, _09182_, _07730_);
  or (_31454_, _31403_, _07012_);
  or (_31457_, _31454_, _31453_);
  or (_31458_, _31411_, _09827_);
  and (_31459_, _31458_, _05669_);
  and (_31460_, _31459_, _31457_);
  and (_31461_, _31460_, _31452_);
  and (_31462_, _14580_, _07730_);
  or (_31463_, _31462_, _31403_);
  and (_31464_, _31463_, _09833_);
  or (_31465_, _31464_, _06019_);
  or (_31466_, _31465_, _31461_);
  and (_31467_, _31466_, _31409_);
  or (_31468_, _31467_, _06112_);
  and (_31469_, _14596_, _07730_);
  or (_31470_, _31403_, _08751_);
  or (_31471_, _31470_, _31469_);
  and (_31472_, _31471_, _08756_);
  and (_31473_, _31472_, _31468_);
  and (_31474_, _10991_, _07730_);
  or (_31475_, _31474_, _31403_);
  and (_31476_, _31475_, _06284_);
  or (_31479_, _31476_, _31473_);
  and (_31480_, _31479_, _07032_);
  or (_31481_, _31480_, _31408_);
  and (_31482_, _31481_, _06278_);
  and (_31483_, _31418_, _06277_);
  and (_31484_, _31483_, _31404_);
  or (_31485_, _31484_, _06130_);
  or (_31486_, _31485_, _31482_);
  and (_31487_, _14593_, _07730_);
  or (_31488_, _31403_, _08777_);
  or (_31489_, _31488_, _31487_);
  and (_31490_, _31489_, _08782_);
  and (_31491_, _31490_, _31486_);
  nor (_31492_, _10990_, _13006_);
  or (_31493_, _31492_, _31403_);
  and (_31494_, _31493_, _06292_);
  or (_31495_, _31494_, _06316_);
  or (_31496_, _31495_, _31491_);
  or (_31497_, _31415_, _06718_);
  and (_31498_, _31497_, _05653_);
  and (_31501_, _31498_, _31496_);
  and (_31502_, _31439_, _05652_);
  or (_31503_, _31502_, _06047_);
  or (_31504_, _31503_, _31501_);
  and (_31505_, _14657_, _07730_);
  or (_31506_, _31403_, _06048_);
  or (_31507_, _31506_, _31505_);
  and (_31508_, _31507_, _01336_);
  and (_31509_, _31508_, _31504_);
  or (_43453_, _31509_, _31402_);
  and (_31510_, _13006_, \oc8051_golden_model_1.P0 [3]);
  and (_31511_, _07730_, _08662_);
  or (_31512_, _31511_, _31510_);
  or (_31513_, _31512_, _06020_);
  and (_31514_, _14672_, _07730_);
  or (_31515_, _31514_, _31510_);
  or (_31516_, _31515_, _06954_);
  and (_31517_, _07730_, \oc8051_golden_model_1.ACC [3]);
  or (_31518_, _31517_, _31510_);
  and (_31519_, _31518_, _06938_);
  and (_31522_, _06939_, \oc8051_golden_model_1.P0 [3]);
  or (_31523_, _31522_, _06102_);
  or (_31524_, _31523_, _31519_);
  and (_31525_, _31524_, _06044_);
  and (_31526_, _31525_, _31516_);
  and (_31527_, _13025_, \oc8051_golden_model_1.P0 [3]);
  and (_31528_, _14683_, _07638_);
  or (_31529_, _31528_, _31527_);
  and (_31530_, _31529_, _06043_);
  or (_31531_, _31530_, _06239_);
  or (_31532_, _31531_, _31526_);
  nor (_31533_, _13006_, _07353_);
  or (_31534_, _31533_, _31510_);
  or (_31535_, _31534_, _06848_);
  and (_31536_, _31535_, _31532_);
  or (_31537_, _31536_, _06219_);
  or (_31538_, _31518_, _06220_);
  and (_31539_, _31538_, _06040_);
  and (_31540_, _31539_, _31537_);
  and (_31541_, _14681_, _07638_);
  or (_31544_, _31541_, _31527_);
  and (_31545_, _31544_, _06039_);
  or (_31546_, _31545_, _06032_);
  or (_31547_, _31546_, _31540_);
  or (_31548_, _31527_, _14708_);
  and (_31549_, _31548_, _31529_);
  or (_31550_, _31549_, _06033_);
  and (_31551_, _31550_, _06027_);
  and (_31552_, _31551_, _31547_);
  and (_31553_, _14724_, _07638_);
  or (_31554_, _31553_, _31527_);
  and (_31555_, _31554_, _06026_);
  or (_31556_, _31555_, _09818_);
  or (_31557_, _31556_, _31552_);
  and (_31558_, _09181_, _07730_);
  or (_31559_, _31510_, _07012_);
  or (_31560_, _31559_, _31558_);
  or (_31561_, _31534_, _09827_);
  and (_31562_, _31561_, _05669_);
  and (_31563_, _31562_, _31560_);
  and (_31566_, _31563_, _31557_);
  and (_31567_, _14778_, _07730_);
  or (_31568_, _31567_, _31510_);
  and (_31569_, _31568_, _09833_);
  or (_31570_, _31569_, _06019_);
  or (_31571_, _31570_, _31566_);
  and (_31572_, _31571_, _31513_);
  or (_31573_, _31572_, _06112_);
  and (_31574_, _14793_, _07730_);
  or (_31575_, _31510_, _08751_);
  or (_31576_, _31575_, _31574_);
  and (_31577_, _31576_, _08756_);
  and (_31578_, _31577_, _31573_);
  and (_31579_, _12299_, _07730_);
  or (_31580_, _31579_, _31510_);
  and (_31581_, _31580_, _06284_);
  or (_31582_, _31581_, _31578_);
  and (_31583_, _31582_, _07032_);
  or (_31584_, _31510_, _08029_);
  and (_31585_, _31512_, _06108_);
  and (_31588_, _31585_, _31584_);
  or (_31589_, _31588_, _31583_);
  and (_31590_, _31589_, _06278_);
  and (_31591_, _31518_, _06277_);
  and (_31592_, _31591_, _31584_);
  or (_31593_, _31592_, _06130_);
  or (_31594_, _31593_, _31590_);
  and (_31595_, _14792_, _07730_);
  or (_31596_, _31510_, _08777_);
  or (_31597_, _31596_, _31595_);
  and (_31598_, _31597_, _08782_);
  and (_31599_, _31598_, _31594_);
  nor (_31600_, _10988_, _13006_);
  or (_31601_, _31600_, _31510_);
  and (_31602_, _31601_, _06292_);
  or (_31603_, _31602_, _06316_);
  or (_31604_, _31603_, _31599_);
  or (_31605_, _31515_, _06718_);
  and (_31606_, _31605_, _05653_);
  and (_31607_, _31606_, _31604_);
  and (_31610_, _31544_, _05652_);
  or (_31611_, _31610_, _06047_);
  or (_31612_, _31611_, _31607_);
  and (_31613_, _14849_, _07730_);
  or (_31614_, _31510_, _06048_);
  or (_31615_, _31614_, _31613_);
  and (_31616_, _31615_, _01336_);
  and (_31617_, _31616_, _31612_);
  nor (_31618_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_31619_, _31618_, _00000_);
  or (_43454_, _31619_, _31617_);
  nor (_31620_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_31621_, _31620_, _00000_);
  and (_31622_, _13006_, \oc8051_golden_model_1.P0 [4]);
  and (_31623_, _08665_, _07730_);
  or (_31624_, _31623_, _31622_);
  or (_31625_, _31624_, _06020_);
  and (_31626_, _14887_, _07730_);
  or (_31627_, _31626_, _31622_);
  or (_31628_, _31627_, _06954_);
  and (_31631_, _07730_, \oc8051_golden_model_1.ACC [4]);
  or (_31632_, _31631_, _31622_);
  and (_31633_, _31632_, _06938_);
  and (_31634_, _06939_, \oc8051_golden_model_1.P0 [4]);
  or (_31635_, _31634_, _06102_);
  or (_31636_, _31635_, _31633_);
  and (_31637_, _31636_, _06044_);
  and (_31638_, _31637_, _31628_);
  and (_31639_, _13025_, \oc8051_golden_model_1.P0 [4]);
  and (_31640_, _14878_, _07638_);
  or (_31641_, _31640_, _31639_);
  and (_31642_, _31641_, _06043_);
  or (_31643_, _31642_, _06239_);
  or (_31644_, _31643_, _31638_);
  nor (_31645_, _08270_, _13006_);
  or (_31646_, _31645_, _31622_);
  or (_31647_, _31646_, _06848_);
  and (_31648_, _31647_, _31644_);
  or (_31649_, _31648_, _06219_);
  or (_31650_, _31632_, _06220_);
  and (_31653_, _31650_, _06040_);
  and (_31654_, _31653_, _31649_);
  and (_31655_, _14882_, _07638_);
  or (_31656_, _31655_, _31639_);
  and (_31657_, _31656_, _06039_);
  or (_31658_, _31657_, _06032_);
  or (_31659_, _31658_, _31654_);
  or (_31660_, _31639_, _14914_);
  and (_31661_, _31660_, _31641_);
  or (_31662_, _31661_, _06033_);
  and (_31663_, _31662_, _06027_);
  and (_31664_, _31663_, _31659_);
  or (_31665_, _31639_, _14879_);
  and (_31666_, _31665_, _06026_);
  and (_31667_, _31666_, _31641_);
  or (_31668_, _31667_, _09818_);
  or (_31669_, _31668_, _31664_);
  and (_31670_, _09180_, _07730_);
  or (_31671_, _31622_, _07012_);
  or (_31672_, _31671_, _31670_);
  or (_31675_, _31646_, _09827_);
  and (_31676_, _31675_, _05669_);
  and (_31677_, _31676_, _31672_);
  and (_31678_, _31677_, _31669_);
  and (_31679_, _14983_, _07730_);
  or (_31680_, _31679_, _31622_);
  and (_31681_, _31680_, _09833_);
  or (_31682_, _31681_, _06019_);
  or (_31683_, _31682_, _31678_);
  and (_31684_, _31683_, _31625_);
  or (_31685_, _31684_, _06112_);
  and (_31686_, _14876_, _07730_);
  or (_31687_, _31686_, _31622_);
  or (_31688_, _31687_, _08751_);
  and (_31689_, _31688_, _08756_);
  and (_31690_, _31689_, _31685_);
  and (_31691_, _10986_, _07730_);
  or (_31692_, _31691_, _31622_);
  and (_31693_, _31692_, _06284_);
  or (_31694_, _31693_, _31690_);
  and (_31697_, _31694_, _07032_);
  or (_31698_, _31622_, _08273_);
  and (_31699_, _31624_, _06108_);
  and (_31700_, _31699_, _31698_);
  or (_31701_, _31700_, _31697_);
  and (_31702_, _31701_, _06278_);
  and (_31703_, _31632_, _06277_);
  and (_31704_, _31703_, _31698_);
  or (_31705_, _31704_, _06130_);
  or (_31706_, _31705_, _31702_);
  and (_31707_, _14873_, _07730_);
  or (_31708_, _31622_, _08777_);
  or (_31709_, _31708_, _31707_);
  and (_31710_, _31709_, _08782_);
  and (_31711_, _31710_, _31706_);
  nor (_31712_, _10985_, _13006_);
  or (_31713_, _31712_, _31622_);
  and (_31714_, _31713_, _06292_);
  or (_31715_, _31714_, _06316_);
  or (_31716_, _31715_, _31711_);
  or (_31719_, _31627_, _06718_);
  and (_31720_, _31719_, _05653_);
  and (_31721_, _31720_, _31716_);
  and (_31722_, _31656_, _05652_);
  or (_31723_, _31722_, _06047_);
  or (_31724_, _31723_, _31721_);
  and (_31725_, _15055_, _07730_);
  or (_31726_, _31622_, _06048_);
  or (_31727_, _31726_, _31725_);
  and (_31728_, _31727_, _01336_);
  and (_31729_, _31728_, _31724_);
  or (_43455_, _31729_, _31621_);
  and (_31730_, _13006_, \oc8051_golden_model_1.P0 [5]);
  and (_31731_, _08652_, _07730_);
  or (_31732_, _31731_, _31730_);
  or (_31733_, _31732_, _06020_);
  and (_31734_, _15093_, _07730_);
  or (_31735_, _31734_, _31730_);
  or (_31736_, _31735_, _06954_);
  and (_31737_, _07730_, \oc8051_golden_model_1.ACC [5]);
  or (_31740_, _31737_, _31730_);
  and (_31741_, _31740_, _06938_);
  and (_31742_, _06939_, \oc8051_golden_model_1.P0 [5]);
  or (_31743_, _31742_, _06102_);
  or (_31744_, _31743_, _31741_);
  and (_31745_, _31744_, _06044_);
  and (_31746_, _31745_, _31736_);
  and (_31747_, _13025_, \oc8051_golden_model_1.P0 [5]);
  and (_31748_, _15073_, _07638_);
  or (_31749_, _31748_, _31747_);
  and (_31750_, _31749_, _06043_);
  or (_31751_, _31750_, _06239_);
  or (_31752_, _31751_, _31746_);
  nor (_31753_, _07977_, _13006_);
  or (_31754_, _31753_, _31730_);
  or (_31755_, _31754_, _06848_);
  and (_31756_, _31755_, _31752_);
  or (_31757_, _31756_, _06219_);
  or (_31758_, _31740_, _06220_);
  and (_31759_, _31758_, _06040_);
  and (_31762_, _31759_, _31757_);
  and (_31763_, _15077_, _07638_);
  or (_31764_, _31763_, _31747_);
  and (_31765_, _31764_, _06039_);
  or (_31766_, _31765_, _06032_);
  or (_31767_, _31766_, _31762_);
  or (_31768_, _31747_, _15110_);
  and (_31769_, _31768_, _31749_);
  or (_31770_, _31769_, _06033_);
  and (_31771_, _31770_, _06027_);
  and (_31772_, _31771_, _31767_);
  or (_31773_, _31747_, _15074_);
  and (_31774_, _31773_, _06026_);
  and (_31775_, _31774_, _31749_);
  or (_31776_, _31775_, _09818_);
  or (_31777_, _31776_, _31772_);
  and (_31778_, _09179_, _07730_);
  or (_31779_, _31730_, _07012_);
  or (_31780_, _31779_, _31778_);
  or (_31781_, _31754_, _09827_);
  and (_31784_, _31781_, _05669_);
  and (_31785_, _31784_, _31780_);
  and (_31786_, _31785_, _31777_);
  and (_31787_, _15179_, _07730_);
  or (_31788_, _31787_, _31730_);
  and (_31789_, _31788_, _09833_);
  or (_31790_, _31789_, _06019_);
  or (_31791_, _31790_, _31786_);
  and (_31792_, _31791_, _31733_);
  or (_31793_, _31792_, _06112_);
  and (_31794_, _15195_, _07730_);
  or (_31795_, _31794_, _31730_);
  or (_31796_, _31795_, _08751_);
  and (_31797_, _31796_, _08756_);
  and (_31798_, _31797_, _31793_);
  and (_31799_, _12306_, _07730_);
  or (_31800_, _31799_, _31730_);
  and (_31801_, _31800_, _06284_);
  or (_31802_, _31801_, _31798_);
  and (_31803_, _31802_, _07032_);
  or (_31806_, _31730_, _07980_);
  and (_31807_, _31732_, _06108_);
  and (_31808_, _31807_, _31806_);
  or (_31809_, _31808_, _31803_);
  and (_31810_, _31809_, _06278_);
  and (_31811_, _31740_, _06277_);
  and (_31812_, _31811_, _31806_);
  or (_31813_, _31812_, _06130_);
  or (_31814_, _31813_, _31810_);
  and (_31815_, _15194_, _07730_);
  or (_31816_, _31730_, _08777_);
  or (_31817_, _31816_, _31815_);
  and (_31818_, _31817_, _08782_);
  and (_31819_, _31818_, _31814_);
  nor (_31820_, _10982_, _13006_);
  or (_31821_, _31820_, _31730_);
  and (_31822_, _31821_, _06292_);
  or (_31823_, _31822_, _06316_);
  or (_31824_, _31823_, _31819_);
  or (_31825_, _31735_, _06718_);
  and (_31828_, _31825_, _05653_);
  and (_31829_, _31828_, _31824_);
  and (_31830_, _31764_, _05652_);
  or (_31831_, _31830_, _06047_);
  or (_31832_, _31831_, _31829_);
  and (_31833_, _15253_, _07730_);
  or (_31834_, _31730_, _06048_);
  or (_31835_, _31834_, _31833_);
  and (_31836_, _31835_, _01336_);
  and (_31837_, _31836_, _31832_);
  nor (_31838_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_31839_, _31838_, _00000_);
  or (_43456_, _31839_, _31837_);
  nor (_31840_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_31841_, _31840_, _00000_);
  and (_31842_, _13006_, \oc8051_golden_model_1.P0 [6]);
  and (_31843_, _15389_, _07730_);
  or (_31844_, _31843_, _31842_);
  or (_31845_, _31844_, _06020_);
  and (_31846_, _15293_, _07730_);
  or (_31849_, _31846_, _31842_);
  or (_31850_, _31849_, _06954_);
  and (_31851_, _07730_, \oc8051_golden_model_1.ACC [6]);
  or (_31852_, _31851_, _31842_);
  and (_31853_, _31852_, _06938_);
  and (_31854_, _06939_, \oc8051_golden_model_1.P0 [6]);
  or (_31855_, _31854_, _06102_);
  or (_31856_, _31855_, _31853_);
  and (_31857_, _31856_, _06044_);
  and (_31858_, _31857_, _31850_);
  and (_31860_, _13025_, \oc8051_golden_model_1.P0 [6]);
  and (_31861_, _15280_, _07638_);
  or (_31862_, _31861_, _31860_);
  and (_31863_, _31862_, _06043_);
  or (_31864_, _31863_, _06239_);
  or (_31865_, _31864_, _31858_);
  nor (_31866_, _07883_, _13006_);
  or (_31867_, _31866_, _31842_);
  or (_31868_, _31867_, _06848_);
  and (_31869_, _31868_, _31865_);
  or (_31871_, _31869_, _06219_);
  or (_31872_, _31852_, _06220_);
  and (_31873_, _31872_, _06040_);
  and (_31874_, _31873_, _31871_);
  and (_31875_, _15278_, _07638_);
  or (_31876_, _31875_, _31860_);
  and (_31877_, _31876_, _06039_);
  or (_31878_, _31877_, _06032_);
  or (_31879_, _31878_, _31874_);
  or (_31880_, _31860_, _15310_);
  and (_31882_, _31880_, _31862_);
  or (_31883_, _31882_, _06033_);
  and (_31884_, _31883_, _06027_);
  and (_31885_, _31884_, _31879_);
  or (_31886_, _31860_, _15326_);
  and (_31887_, _31886_, _06026_);
  and (_31888_, _31887_, _31862_);
  or (_31889_, _31888_, _09818_);
  or (_31890_, _31889_, _31885_);
  and (_31891_, _09178_, _07730_);
  or (_31893_, _31842_, _07012_);
  or (_31894_, _31893_, _31891_);
  or (_31895_, _31867_, _09827_);
  and (_31896_, _31895_, _05669_);
  and (_31897_, _31896_, _31894_);
  and (_31898_, _31897_, _31890_);
  and (_31899_, _15382_, _07730_);
  or (_31900_, _31899_, _31842_);
  and (_31901_, _31900_, _09833_);
  or (_31902_, _31901_, _06019_);
  or (_31904_, _31902_, _31898_);
  and (_31905_, _31904_, _31845_);
  or (_31906_, _31905_, _06112_);
  and (_31907_, _15399_, _07730_);
  or (_31908_, _31842_, _08751_);
  or (_31909_, _31908_, _31907_);
  and (_31910_, _31909_, _08756_);
  and (_31911_, _31910_, _31906_);
  and (_31912_, _10980_, _07730_);
  or (_31913_, _31912_, _31842_);
  and (_31915_, _31913_, _06284_);
  or (_31916_, _31915_, _31911_);
  and (_31917_, _31916_, _07032_);
  or (_31918_, _31842_, _07886_);
  and (_31919_, _31844_, _06108_);
  and (_31920_, _31919_, _31918_);
  or (_31921_, _31920_, _31917_);
  and (_31922_, _31921_, _06278_);
  and (_31923_, _31852_, _06277_);
  and (_31924_, _31923_, _31918_);
  or (_31925_, _31924_, _06130_);
  or (_31926_, _31925_, _31922_);
  and (_31927_, _15396_, _07730_);
  or (_31928_, _31842_, _08777_);
  or (_31929_, _31928_, _31927_);
  and (_31930_, _31929_, _08782_);
  and (_31931_, _31930_, _31926_);
  nor (_31932_, _10979_, _13006_);
  or (_31933_, _31932_, _31842_);
  and (_31934_, _31933_, _06292_);
  or (_31936_, _31934_, _06316_);
  or (_31937_, _31936_, _31931_);
  or (_31938_, _31849_, _06718_);
  and (_31939_, _31938_, _05653_);
  and (_31940_, _31939_, _31937_);
  and (_31941_, _31876_, _05652_);
  or (_31942_, _31941_, _06047_);
  or (_31943_, _31942_, _31940_);
  and (_31944_, _15451_, _07730_);
  or (_31945_, _31842_, _06048_);
  or (_31947_, _31945_, _31944_);
  and (_31948_, _31947_, _01336_);
  and (_31949_, _31948_, _31943_);
  or (_43457_, _31949_, _31841_);
  nor (_31950_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_31951_, _31950_, _00000_);
  and (_31952_, _07677_, \oc8051_golden_model_1.ACC [0]);
  and (_31953_, _31952_, _08127_);
  and (_31954_, _13108_, \oc8051_golden_model_1.P1 [0]);
  or (_31955_, _31954_, _06278_);
  or (_31957_, _31955_, _31953_);
  and (_31958_, _07677_, _08672_);
  or (_31959_, _31958_, _31954_);
  or (_31960_, _31959_, _06020_);
  and (_31961_, _09120_, _07677_);
  or (_31962_, _31954_, _07012_);
  or (_31963_, _31962_, _31961_);
  nor (_31964_, _08127_, _13108_);
  or (_31965_, _31964_, _31954_);
  and (_31966_, _31965_, _06102_);
  and (_31968_, _06939_, \oc8051_golden_model_1.P1 [0]);
  or (_31969_, _31952_, _31954_);
  and (_31970_, _31969_, _06938_);
  or (_31971_, _31970_, _31968_);
  and (_31972_, _31971_, _06954_);
  or (_31973_, _31972_, _06043_);
  or (_31974_, _31973_, _31966_);
  and (_31975_, _14102_, _08345_);
  and (_31976_, _13127_, \oc8051_golden_model_1.P1 [0]);
  or (_31977_, _31976_, _06044_);
  or (_31979_, _31977_, _31975_);
  and (_31980_, _31979_, _06848_);
  and (_31981_, _31980_, _31974_);
  and (_31982_, _07677_, _06931_);
  or (_31983_, _31982_, _31954_);
  and (_31984_, _31983_, _06239_);
  or (_31985_, _31984_, _06219_);
  or (_31986_, _31985_, _31981_);
  or (_31987_, _31969_, _06220_);
  and (_31988_, _31987_, _06040_);
  and (_31990_, _31988_, _31986_);
  and (_31991_, _31954_, _06039_);
  or (_31992_, _31991_, _06032_);
  or (_31993_, _31992_, _31990_);
  or (_31994_, _31965_, _06033_);
  and (_31995_, _31994_, _06027_);
  and (_31996_, _31995_, _31993_);
  and (_31997_, _14132_, _08345_);
  or (_31998_, _31997_, _31976_);
  and (_31999_, _31998_, _06026_);
  or (_32001_, _31999_, _09818_);
  or (_32002_, _32001_, _31996_);
  or (_32003_, _31983_, _09827_);
  and (_32004_, _32003_, _05669_);
  and (_32005_, _32004_, _32002_);
  and (_32006_, _32005_, _31963_);
  and (_32007_, _14186_, _07677_);
  or (_32008_, _32007_, _31954_);
  and (_32009_, _32008_, _09833_);
  or (_32010_, _32009_, _06019_);
  or (_32012_, _32010_, _32006_);
  and (_32013_, _32012_, _31960_);
  or (_32014_, _32013_, _06112_);
  and (_32015_, _14086_, _07677_);
  or (_32016_, _32015_, _31954_);
  or (_32017_, _32016_, _08751_);
  and (_32018_, _32017_, _08756_);
  and (_32019_, _32018_, _32014_);
  nor (_32020_, _12302_, _13108_);
  or (_32021_, _32020_, _31954_);
  nor (_32023_, _31953_, _08756_);
  and (_32024_, _32023_, _32021_);
  or (_32025_, _32024_, _32019_);
  and (_32026_, _32025_, _07032_);
  nand (_32027_, _31959_, _06108_);
  nor (_32028_, _32027_, _31964_);
  or (_32029_, _32028_, _06277_);
  or (_32030_, _32029_, _32026_);
  and (_32031_, _32030_, _31957_);
  or (_32032_, _32031_, _06130_);
  and (_32034_, _14083_, _07677_);
  or (_32035_, _31954_, _08777_);
  or (_32036_, _32035_, _32034_);
  and (_32037_, _32036_, _08782_);
  and (_32038_, _32037_, _32032_);
  and (_32039_, _32021_, _06292_);
  or (_32040_, _32039_, _06316_);
  or (_32041_, _32040_, _32038_);
  or (_32042_, _31965_, _06718_);
  and (_32043_, _32042_, _32041_);
  or (_32045_, _32043_, _05652_);
  or (_32046_, _31954_, _05653_);
  and (_32047_, _32046_, _32045_);
  or (_32048_, _32047_, _06047_);
  or (_32049_, _31965_, _06048_);
  and (_32050_, _32049_, _01336_);
  and (_32051_, _32050_, _32048_);
  or (_43459_, _32051_, _31951_);
  and (_32052_, _13108_, \oc8051_golden_model_1.P1 [1]);
  nor (_32053_, _10993_, _13108_);
  or (_32055_, _32053_, _32052_);
  or (_32056_, _32055_, _08782_);
  or (_32057_, _14367_, _13108_);
  or (_32058_, _07677_, \oc8051_golden_model_1.P1 [1]);
  and (_32059_, _32058_, _09833_);
  and (_32060_, _32059_, _32057_);
  nor (_32061_, _13108_, _07132_);
  or (_32062_, _32061_, _32052_);
  and (_32063_, _32062_, _06239_);
  and (_32064_, _13127_, \oc8051_golden_model_1.P1 [1]);
  and (_32066_, _14266_, _08345_);
  or (_32067_, _32066_, _32064_);
  or (_32068_, _32067_, _06044_);
  and (_32069_, _14284_, _07677_);
  not (_32070_, _32069_);
  and (_32071_, _32070_, _32058_);
  and (_32072_, _32071_, _06102_);
  and (_32073_, _06939_, \oc8051_golden_model_1.P1 [1]);
  and (_32074_, _07677_, \oc8051_golden_model_1.ACC [1]);
  or (_32075_, _32074_, _32052_);
  and (_32077_, _32075_, _06938_);
  or (_32078_, _32077_, _32073_);
  and (_32079_, _32078_, _06954_);
  or (_32080_, _32079_, _06043_);
  or (_32081_, _32080_, _32072_);
  and (_32082_, _32081_, _32068_);
  and (_32083_, _32082_, _06848_);
  or (_32084_, _32083_, _32063_);
  or (_32085_, _32084_, _06219_);
  or (_32086_, _32075_, _06220_);
  and (_32088_, _32086_, _06040_);
  and (_32089_, _32088_, _32085_);
  and (_32090_, _14273_, _08345_);
  or (_32091_, _32090_, _32064_);
  and (_32092_, _32091_, _06039_);
  or (_32093_, _32092_, _06032_);
  or (_32094_, _32093_, _32089_);
  or (_32095_, _32064_, _14302_);
  and (_32096_, _32095_, _32067_);
  or (_32097_, _32096_, _06033_);
  and (_32099_, _32097_, _06027_);
  and (_32100_, _32099_, _32094_);
  or (_32101_, _32064_, _14267_);
  and (_32102_, _32101_, _06026_);
  and (_32103_, _32102_, _32067_);
  or (_32104_, _32103_, _09815_);
  or (_32105_, _32104_, _32100_);
  or (_32106_, _32062_, _09827_);
  and (_32107_, _32106_, _32105_);
  or (_32108_, _32107_, _07011_);
  and (_32110_, _09075_, _07677_);
  or (_32111_, _32052_, _07012_);
  or (_32112_, _32111_, _32110_);
  and (_32113_, _32112_, _05669_);
  and (_32114_, _32113_, _32108_);
  or (_32115_, _32114_, _32060_);
  and (_32116_, _32115_, _06020_);
  nand (_32117_, _07677_, _06832_);
  and (_32118_, _32058_, _06019_);
  and (_32119_, _32118_, _32117_);
  or (_32121_, _32119_, _32116_);
  and (_32122_, _32121_, _08751_);
  or (_32123_, _14263_, _13108_);
  and (_32124_, _32058_, _06112_);
  and (_32125_, _32124_, _32123_);
  or (_32126_, _32125_, _06284_);
  or (_32127_, _32126_, _32122_);
  nand (_32128_, _10992_, _07677_);
  and (_32129_, _32128_, _32055_);
  or (_32130_, _32129_, _08756_);
  and (_32132_, _32130_, _07032_);
  and (_32133_, _32132_, _32127_);
  or (_32134_, _14261_, _13108_);
  and (_32135_, _32058_, _06108_);
  and (_32136_, _32135_, _32134_);
  or (_32137_, _32136_, _06277_);
  or (_32138_, _32137_, _32133_);
  nor (_32139_, _32052_, _06278_);
  nand (_32140_, _32139_, _32128_);
  and (_32141_, _32140_, _08777_);
  and (_32143_, _32141_, _32138_);
  or (_32144_, _32117_, _08078_);
  and (_32145_, _32058_, _06130_);
  and (_32146_, _32145_, _32144_);
  or (_32147_, _32146_, _06292_);
  or (_32148_, _32147_, _32143_);
  and (_32149_, _32148_, _32056_);
  or (_32150_, _32149_, _06316_);
  or (_32151_, _32071_, _06718_);
  and (_32152_, _32151_, _05653_);
  and (_32154_, _32152_, _32150_);
  and (_32155_, _32091_, _05652_);
  or (_32156_, _32155_, _06047_);
  or (_32157_, _32156_, _32154_);
  or (_32158_, _32052_, _06048_);
  or (_32159_, _32158_, _32069_);
  and (_32160_, _32159_, _01336_);
  and (_32161_, _32160_, _32157_);
  nor (_32162_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_32163_, _32162_, _00000_);
  or (_43460_, _32163_, _32161_);
  nor (_32165_, \oc8051_golden_model_1.P1 [2], rst);
  nor (_32166_, _32165_, _00000_);
  and (_32167_, _13108_, \oc8051_golden_model_1.P1 [2]);
  and (_32168_, _07677_, _08730_);
  or (_32169_, _32168_, _32167_);
  or (_32170_, _32169_, _06020_);
  nor (_32171_, _13108_, _07530_);
  or (_32172_, _32171_, _32167_);
  and (_32173_, _32172_, _06239_);
  and (_32175_, _13127_, \oc8051_golden_model_1.P1 [2]);
  and (_32176_, _14497_, _08345_);
  or (_32177_, _32176_, _32175_);
  or (_32178_, _32177_, _06044_);
  and (_32179_, _14493_, _07677_);
  or (_32180_, _32179_, _32167_);
  and (_32181_, _32180_, _06102_);
  and (_32182_, _06939_, \oc8051_golden_model_1.P1 [2]);
  and (_32183_, _07677_, \oc8051_golden_model_1.ACC [2]);
  or (_32184_, _32183_, _32167_);
  and (_32186_, _32184_, _06938_);
  or (_32187_, _32186_, _32182_);
  and (_32188_, _32187_, _06954_);
  or (_32189_, _32188_, _06043_);
  or (_32190_, _32189_, _32181_);
  and (_32191_, _32190_, _32178_);
  and (_32192_, _32191_, _06848_);
  or (_32193_, _32192_, _32173_);
  or (_32194_, _32193_, _06219_);
  or (_32195_, _32184_, _06220_);
  and (_32197_, _32195_, _06040_);
  and (_32198_, _32197_, _32194_);
  and (_32199_, _14479_, _08345_);
  or (_32200_, _32199_, _32175_);
  and (_32201_, _32200_, _06039_);
  or (_32202_, _32201_, _06032_);
  or (_32203_, _32202_, _32198_);
  or (_32204_, _32175_, _14512_);
  and (_32205_, _32204_, _32177_);
  or (_32206_, _32205_, _06033_);
  and (_32208_, _32206_, _06027_);
  and (_32209_, _32208_, _32203_);
  or (_32210_, _32175_, _14525_);
  and (_32211_, _32210_, _06026_);
  and (_32212_, _32211_, _32177_);
  or (_32213_, _32212_, _09818_);
  or (_32214_, _32213_, _32209_);
  and (_32215_, _09182_, _07677_);
  or (_32216_, _32167_, _07012_);
  or (_32217_, _32216_, _32215_);
  or (_32219_, _32172_, _09827_);
  and (_32220_, _32219_, _05669_);
  and (_32221_, _32220_, _32217_);
  and (_32222_, _32221_, _32214_);
  and (_32223_, _14580_, _07677_);
  or (_32224_, _32223_, _32167_);
  and (_32225_, _32224_, _09833_);
  or (_32226_, _32225_, _06019_);
  or (_32227_, _32226_, _32222_);
  and (_32228_, _32227_, _32170_);
  or (_32230_, _32228_, _06112_);
  and (_32231_, _14596_, _07677_);
  or (_32232_, _32167_, _08751_);
  or (_32233_, _32232_, _32231_);
  and (_32234_, _32233_, _08756_);
  and (_32235_, _32234_, _32230_);
  and (_32236_, _10991_, _07677_);
  or (_32237_, _32236_, _32167_);
  and (_32238_, _32237_, _06284_);
  or (_32239_, _32238_, _32235_);
  and (_32241_, _32239_, _07032_);
  or (_32242_, _32167_, _08177_);
  and (_32243_, _32169_, _06108_);
  and (_32244_, _32243_, _32242_);
  or (_32245_, _32244_, _32241_);
  and (_32246_, _32245_, _06278_);
  and (_32247_, _32184_, _06277_);
  and (_32248_, _32247_, _32242_);
  or (_32249_, _32248_, _06130_);
  or (_32250_, _32249_, _32246_);
  and (_32252_, _14593_, _07677_);
  or (_32253_, _32167_, _08777_);
  or (_32254_, _32253_, _32252_);
  and (_32255_, _32254_, _08782_);
  and (_32256_, _32255_, _32250_);
  nor (_32257_, _10990_, _13108_);
  or (_32258_, _32257_, _32167_);
  and (_32259_, _32258_, _06292_);
  or (_32260_, _32259_, _06316_);
  or (_32261_, _32260_, _32256_);
  or (_32263_, _32180_, _06718_);
  and (_32264_, _32263_, _05653_);
  and (_32265_, _32264_, _32261_);
  and (_32266_, _32200_, _05652_);
  or (_32267_, _32266_, _06047_);
  or (_32268_, _32267_, _32265_);
  and (_32269_, _14657_, _07677_);
  or (_32270_, _32167_, _06048_);
  or (_32271_, _32270_, _32269_);
  and (_32272_, _32271_, _01336_);
  and (_32274_, _32272_, _32268_);
  or (_43461_, _32274_, _32166_);
  and (_32275_, _13108_, \oc8051_golden_model_1.P1 [3]);
  and (_32276_, _07677_, _08662_);
  or (_32277_, _32276_, _32275_);
  or (_32278_, _32277_, _06020_);
  and (_32279_, _14672_, _07677_);
  or (_32280_, _32279_, _32275_);
  or (_32281_, _32280_, _06954_);
  and (_32282_, _07677_, \oc8051_golden_model_1.ACC [3]);
  or (_32284_, _32282_, _32275_);
  and (_32285_, _32284_, _06938_);
  and (_32286_, _06939_, \oc8051_golden_model_1.P1 [3]);
  or (_32287_, _32286_, _06102_);
  or (_32288_, _32287_, _32285_);
  and (_32289_, _32288_, _06044_);
  and (_32290_, _32289_, _32281_);
  and (_32291_, _13127_, \oc8051_golden_model_1.P1 [3]);
  and (_32292_, _14683_, _08345_);
  or (_32293_, _32292_, _32291_);
  and (_32295_, _32293_, _06043_);
  or (_32296_, _32295_, _06239_);
  or (_32297_, _32296_, _32290_);
  nor (_32298_, _13108_, _07353_);
  or (_32299_, _32298_, _32275_);
  or (_32300_, _32299_, _06848_);
  and (_32301_, _32300_, _32297_);
  or (_32302_, _32301_, _06219_);
  or (_32303_, _32284_, _06220_);
  and (_32304_, _32303_, _06040_);
  and (_32306_, _32304_, _32302_);
  and (_32307_, _14681_, _08345_);
  or (_32308_, _32307_, _32291_);
  and (_32309_, _32308_, _06039_);
  or (_32310_, _32309_, _06032_);
  or (_32311_, _32310_, _32306_);
  or (_32312_, _32291_, _14708_);
  and (_32313_, _32312_, _32293_);
  or (_32314_, _32313_, _06033_);
  and (_32315_, _32314_, _06027_);
  and (_32317_, _32315_, _32311_);
  and (_32318_, _14724_, _08345_);
  or (_32319_, _32318_, _32291_);
  and (_32320_, _32319_, _06026_);
  or (_32321_, _32320_, _09818_);
  or (_32322_, _32321_, _32317_);
  and (_32323_, _09181_, _07677_);
  or (_32324_, _32275_, _07012_);
  or (_32325_, _32324_, _32323_);
  or (_32326_, _32299_, _09827_);
  and (_32328_, _32326_, _05669_);
  and (_32329_, _32328_, _32325_);
  and (_32330_, _32329_, _32322_);
  and (_32331_, _14778_, _07677_);
  or (_32332_, _32331_, _32275_);
  and (_32333_, _32332_, _09833_);
  or (_32334_, _32333_, _06019_);
  or (_32335_, _32334_, _32330_);
  and (_32336_, _32335_, _32278_);
  or (_32337_, _32336_, _06112_);
  and (_32339_, _14793_, _07677_);
  or (_32340_, _32275_, _08751_);
  or (_32341_, _32340_, _32339_);
  and (_32342_, _32341_, _08756_);
  and (_32343_, _32342_, _32337_);
  and (_32344_, _12299_, _07677_);
  or (_32345_, _32344_, _32275_);
  and (_32346_, _32345_, _06284_);
  or (_32347_, _32346_, _32343_);
  and (_32348_, _32347_, _07032_);
  or (_32350_, _32275_, _08029_);
  and (_32351_, _32277_, _06108_);
  and (_32352_, _32351_, _32350_);
  or (_32353_, _32352_, _32348_);
  and (_32354_, _32353_, _06278_);
  and (_32355_, _32284_, _06277_);
  and (_32356_, _32355_, _32350_);
  or (_32357_, _32356_, _06130_);
  or (_32358_, _32357_, _32354_);
  and (_32359_, _14792_, _07677_);
  or (_32361_, _32275_, _08777_);
  or (_32362_, _32361_, _32359_);
  and (_32363_, _32362_, _08782_);
  and (_32364_, _32363_, _32358_);
  nor (_32365_, _10988_, _13108_);
  or (_32366_, _32365_, _32275_);
  and (_32367_, _32366_, _06292_);
  or (_32368_, _32367_, _06316_);
  or (_32369_, _32368_, _32364_);
  or (_32370_, _32280_, _06718_);
  and (_32372_, _32370_, _05653_);
  and (_32373_, _32372_, _32369_);
  and (_32374_, _32308_, _05652_);
  or (_32375_, _32374_, _06047_);
  or (_32376_, _32375_, _32373_);
  and (_32377_, _14849_, _07677_);
  or (_32378_, _32275_, _06048_);
  or (_32379_, _32378_, _32377_);
  and (_32380_, _32379_, _01336_);
  and (_32381_, _32380_, _32376_);
  nor (_32383_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_32384_, _32383_, _00000_);
  or (_43463_, _32384_, _32381_);
  and (_32385_, _13108_, \oc8051_golden_model_1.P1 [4]);
  and (_32386_, _08665_, _07677_);
  or (_32387_, _32386_, _32385_);
  or (_32388_, _32387_, _06020_);
  and (_32389_, _14887_, _07677_);
  or (_32390_, _32389_, _32385_);
  or (_32391_, _32390_, _06954_);
  and (_32393_, _07677_, \oc8051_golden_model_1.ACC [4]);
  or (_32394_, _32393_, _32385_);
  and (_32395_, _32394_, _06938_);
  and (_32396_, _06939_, \oc8051_golden_model_1.P1 [4]);
  or (_32397_, _32396_, _06102_);
  or (_32398_, _32397_, _32395_);
  and (_32399_, _32398_, _06044_);
  and (_32400_, _32399_, _32391_);
  and (_32401_, _13127_, \oc8051_golden_model_1.P1 [4]);
  and (_32402_, _14878_, _08345_);
  or (_32404_, _32402_, _32401_);
  and (_32405_, _32404_, _06043_);
  or (_32406_, _32405_, _06239_);
  or (_32407_, _32406_, _32400_);
  nor (_32408_, _08270_, _13108_);
  or (_32409_, _32408_, _32385_);
  or (_32410_, _32409_, _06848_);
  and (_32411_, _32410_, _32407_);
  or (_32412_, _32411_, _06219_);
  or (_32413_, _32394_, _06220_);
  and (_32415_, _32413_, _06040_);
  and (_32416_, _32415_, _32412_);
  and (_32417_, _14882_, _08345_);
  or (_32418_, _32417_, _32401_);
  and (_32419_, _32418_, _06039_);
  or (_32420_, _32419_, _06032_);
  or (_32421_, _32420_, _32416_);
  or (_32422_, _32401_, _14914_);
  and (_32423_, _32422_, _32404_);
  or (_32424_, _32423_, _06033_);
  and (_32426_, _32424_, _06027_);
  and (_32427_, _32426_, _32421_);
  or (_32428_, _32401_, _14879_);
  and (_32429_, _32428_, _06026_);
  and (_32430_, _32429_, _32404_);
  or (_32431_, _32430_, _09818_);
  or (_32432_, _32431_, _32427_);
  and (_32433_, _09180_, _07677_);
  or (_32434_, _32385_, _07012_);
  or (_32435_, _32434_, _32433_);
  or (_32437_, _32409_, _09827_);
  and (_32438_, _32437_, _05669_);
  and (_32439_, _32438_, _32435_);
  and (_32440_, _32439_, _32432_);
  and (_32441_, _14983_, _07677_);
  or (_32442_, _32441_, _32385_);
  and (_32443_, _32442_, _09833_);
  or (_32444_, _32443_, _06019_);
  or (_32445_, _32444_, _32440_);
  and (_32446_, _32445_, _32388_);
  or (_32448_, _32446_, _06112_);
  and (_32449_, _14876_, _07677_);
  or (_32450_, _32449_, _32385_);
  or (_32451_, _32450_, _08751_);
  and (_32452_, _32451_, _08756_);
  and (_32453_, _32452_, _32448_);
  and (_32454_, _10986_, _07677_);
  or (_32455_, _32454_, _32385_);
  and (_32456_, _32455_, _06284_);
  or (_32457_, _32456_, _32453_);
  and (_32459_, _32457_, _07032_);
  or (_32460_, _32385_, _08273_);
  and (_32461_, _32387_, _06108_);
  and (_32462_, _32461_, _32460_);
  or (_32463_, _32462_, _32459_);
  and (_32464_, _32463_, _06278_);
  and (_32465_, _32394_, _06277_);
  and (_32466_, _32465_, _32460_);
  or (_32467_, _32466_, _06130_);
  or (_32468_, _32467_, _32464_);
  and (_32470_, _14873_, _07677_);
  or (_32471_, _32385_, _08777_);
  or (_32472_, _32471_, _32470_);
  and (_32473_, _32472_, _08782_);
  and (_32474_, _32473_, _32468_);
  nor (_32475_, _10985_, _13108_);
  or (_32476_, _32475_, _32385_);
  and (_32477_, _32476_, _06292_);
  or (_32478_, _32477_, _06316_);
  or (_32479_, _32478_, _32474_);
  or (_32481_, _32390_, _06718_);
  and (_32482_, _32481_, _05653_);
  and (_32483_, _32482_, _32479_);
  and (_32484_, _32418_, _05652_);
  or (_32485_, _32484_, _06047_);
  or (_32486_, _32485_, _32483_);
  and (_32487_, _15055_, _07677_);
  or (_32488_, _32385_, _06048_);
  or (_32489_, _32488_, _32487_);
  and (_32490_, _32489_, _01336_);
  and (_32492_, _32490_, _32486_);
  nor (_32493_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_32494_, _32493_, _00000_);
  or (_43464_, _32494_, _32492_);
  and (_32495_, _13108_, \oc8051_golden_model_1.P1 [5]);
  and (_32496_, _08652_, _07677_);
  or (_32497_, _32496_, _32495_);
  or (_32498_, _32497_, _06020_);
  and (_32499_, _15093_, _07677_);
  or (_32500_, _32499_, _32495_);
  or (_32502_, _32500_, _06954_);
  and (_32503_, _07677_, \oc8051_golden_model_1.ACC [5]);
  or (_32504_, _32503_, _32495_);
  and (_32505_, _32504_, _06938_);
  and (_32506_, _06939_, \oc8051_golden_model_1.P1 [5]);
  or (_32507_, _32506_, _06102_);
  or (_32508_, _32507_, _32505_);
  and (_32509_, _32508_, _06044_);
  and (_32510_, _32509_, _32502_);
  and (_32511_, _13127_, \oc8051_golden_model_1.P1 [5]);
  and (_32513_, _15073_, _08345_);
  or (_32514_, _32513_, _32511_);
  and (_32515_, _32514_, _06043_);
  or (_32516_, _32515_, _06239_);
  or (_32517_, _32516_, _32510_);
  nor (_32518_, _07977_, _13108_);
  or (_32519_, _32518_, _32495_);
  or (_32520_, _32519_, _06848_);
  and (_32521_, _32520_, _32517_);
  or (_32522_, _32521_, _06219_);
  or (_32524_, _32504_, _06220_);
  and (_32525_, _32524_, _06040_);
  and (_32526_, _32525_, _32522_);
  and (_32527_, _15077_, _08345_);
  or (_32528_, _32527_, _32511_);
  and (_32529_, _32528_, _06039_);
  or (_32530_, _32529_, _06032_);
  or (_32531_, _32530_, _32526_);
  or (_32532_, _32511_, _15110_);
  and (_32533_, _32532_, _32514_);
  or (_32535_, _32533_, _06033_);
  and (_32536_, _32535_, _06027_);
  and (_32537_, _32536_, _32531_);
  or (_32538_, _32511_, _15074_);
  and (_32539_, _32538_, _06026_);
  and (_32540_, _32539_, _32514_);
  or (_32541_, _32540_, _09818_);
  or (_32542_, _32541_, _32537_);
  and (_32543_, _09179_, _07677_);
  or (_32544_, _32495_, _07012_);
  or (_32546_, _32544_, _32543_);
  or (_32547_, _32519_, _09827_);
  and (_32548_, _32547_, _05669_);
  and (_32549_, _32548_, _32546_);
  and (_32550_, _32549_, _32542_);
  and (_32551_, _15179_, _07677_);
  or (_32552_, _32551_, _32495_);
  and (_32553_, _32552_, _09833_);
  or (_32554_, _32553_, _06019_);
  or (_32555_, _32554_, _32550_);
  and (_32557_, _32555_, _32498_);
  or (_32558_, _32557_, _06112_);
  and (_32559_, _15195_, _07677_);
  or (_32560_, _32495_, _08751_);
  or (_32561_, _32560_, _32559_);
  and (_32562_, _32561_, _08756_);
  and (_32563_, _32562_, _32558_);
  and (_32564_, _12306_, _07677_);
  or (_32565_, _32564_, _32495_);
  and (_32566_, _32565_, _06284_);
  or (_32568_, _32566_, _32563_);
  and (_32569_, _32568_, _07032_);
  or (_32570_, _32495_, _07980_);
  and (_32571_, _32497_, _06108_);
  and (_32572_, _32571_, _32570_);
  or (_32573_, _32572_, _32569_);
  and (_32574_, _32573_, _06278_);
  and (_32575_, _32504_, _06277_);
  and (_32576_, _32575_, _32570_);
  or (_32577_, _32576_, _06130_);
  or (_32579_, _32577_, _32574_);
  and (_32580_, _15194_, _07677_);
  or (_32581_, _32495_, _08777_);
  or (_32582_, _32581_, _32580_);
  and (_32583_, _32582_, _08782_);
  and (_32584_, _32583_, _32579_);
  nor (_32585_, _10982_, _13108_);
  or (_32586_, _32585_, _32495_);
  and (_32587_, _32586_, _06292_);
  or (_32588_, _32587_, _06316_);
  or (_32590_, _32588_, _32584_);
  or (_32591_, _32500_, _06718_);
  and (_32592_, _32591_, _05653_);
  and (_32593_, _32592_, _32590_);
  and (_32594_, _32528_, _05652_);
  or (_32595_, _32594_, _06047_);
  or (_32596_, _32595_, _32593_);
  and (_32597_, _15253_, _07677_);
  or (_32598_, _32495_, _06048_);
  or (_32599_, _32598_, _32597_);
  and (_32601_, _32599_, _01336_);
  and (_32602_, _32601_, _32596_);
  nor (_32603_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_32604_, _32603_, _00000_);
  or (_43465_, _32604_, _32602_);
  and (_32605_, _13108_, \oc8051_golden_model_1.P1 [6]);
  and (_32606_, _15389_, _07677_);
  or (_32607_, _32606_, _32605_);
  or (_32608_, _32607_, _06020_);
  and (_32609_, _15293_, _07677_);
  or (_32611_, _32609_, _32605_);
  or (_32612_, _32611_, _06954_);
  and (_32613_, _07677_, \oc8051_golden_model_1.ACC [6]);
  or (_32614_, _32613_, _32605_);
  and (_32615_, _32614_, _06938_);
  and (_32616_, _06939_, \oc8051_golden_model_1.P1 [6]);
  or (_32617_, _32616_, _06102_);
  or (_32618_, _32617_, _32615_);
  and (_32619_, _32618_, _06044_);
  and (_32620_, _32619_, _32612_);
  and (_32622_, _13127_, \oc8051_golden_model_1.P1 [6]);
  and (_32623_, _15280_, _08345_);
  or (_32624_, _32623_, _32622_);
  and (_32625_, _32624_, _06043_);
  or (_32626_, _32625_, _06239_);
  or (_32627_, _32626_, _32620_);
  nor (_32628_, _07883_, _13108_);
  or (_32629_, _32628_, _32605_);
  or (_32630_, _32629_, _06848_);
  and (_32631_, _32630_, _32627_);
  or (_32633_, _32631_, _06219_);
  or (_32634_, _32614_, _06220_);
  and (_32635_, _32634_, _06040_);
  and (_32636_, _32635_, _32633_);
  and (_32637_, _15278_, _08345_);
  or (_32638_, _32637_, _32622_);
  and (_32639_, _32638_, _06039_);
  or (_32640_, _32639_, _06032_);
  or (_32641_, _32640_, _32636_);
  or (_32642_, _32622_, _15310_);
  and (_32644_, _32642_, _32624_);
  or (_32645_, _32644_, _06033_);
  and (_32646_, _32645_, _06027_);
  and (_32647_, _32646_, _32641_);
  or (_32648_, _32622_, _15326_);
  and (_32649_, _32648_, _06026_);
  and (_32650_, _32649_, _32624_);
  or (_32651_, _32650_, _09818_);
  or (_32652_, _32651_, _32647_);
  and (_32653_, _09178_, _07677_);
  or (_32654_, _32605_, _07012_);
  or (_32655_, _32654_, _32653_);
  or (_32656_, _32629_, _09827_);
  and (_32657_, _32656_, _05669_);
  and (_32658_, _32657_, _32655_);
  and (_32659_, _32658_, _32652_);
  and (_32660_, _15382_, _07677_);
  or (_32661_, _32660_, _32605_);
  and (_32662_, _32661_, _09833_);
  or (_32663_, _32662_, _06019_);
  or (_32665_, _32663_, _32659_);
  and (_32666_, _32665_, _32608_);
  or (_32667_, _32666_, _06112_);
  and (_32668_, _15399_, _07677_);
  or (_32669_, _32605_, _08751_);
  or (_32670_, _32669_, _32668_);
  and (_32671_, _32670_, _08756_);
  and (_32672_, _32671_, _32667_);
  and (_32673_, _10980_, _07677_);
  or (_32674_, _32673_, _32605_);
  and (_32676_, _32674_, _06284_);
  or (_32677_, _32676_, _32672_);
  and (_32678_, _32677_, _07032_);
  or (_32679_, _32605_, _07886_);
  and (_32680_, _32607_, _06108_);
  and (_32681_, _32680_, _32679_);
  or (_32682_, _32681_, _32678_);
  and (_32683_, _32682_, _06278_);
  and (_32684_, _32614_, _06277_);
  and (_32685_, _32684_, _32679_);
  or (_32687_, _32685_, _06130_);
  or (_32688_, _32687_, _32683_);
  and (_32689_, _15396_, _07677_);
  or (_32690_, _32605_, _08777_);
  or (_32691_, _32690_, _32689_);
  and (_32692_, _32691_, _08782_);
  and (_32693_, _32692_, _32688_);
  nor (_32694_, _10979_, _13108_);
  or (_32695_, _32694_, _32605_);
  and (_32696_, _32695_, _06292_);
  or (_32698_, _32696_, _06316_);
  or (_32699_, _32698_, _32693_);
  or (_32700_, _32611_, _06718_);
  and (_32701_, _32700_, _05653_);
  and (_32702_, _32701_, _32699_);
  and (_32703_, _32638_, _05652_);
  or (_32704_, _32703_, _06047_);
  or (_32705_, _32704_, _32702_);
  and (_32706_, _15451_, _07677_);
  or (_32707_, _32605_, _06048_);
  or (_32709_, _32707_, _32706_);
  and (_32710_, _32709_, _01336_);
  and (_32711_, _32710_, _32705_);
  nor (_32712_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_32713_, _32712_, _00000_);
  or (_43466_, _32713_, _32711_);
  not (_32714_, \oc8051_golden_model_1.IP [0]);
  nor (_32715_, _01336_, _32714_);
  nand (_32716_, _10995_, _07694_);
  nor (_32717_, _07694_, _32714_);
  nor (_32719_, _32717_, _06278_);
  nand (_32720_, _32719_, _32716_);
  and (_32721_, _07694_, _08672_);
  or (_32722_, _32721_, _32717_);
  or (_32723_, _32722_, _06020_);
  and (_32724_, _09120_, _07694_);
  or (_32725_, _32717_, _07012_);
  or (_32726_, _32725_, _32724_);
  nor (_32727_, _08127_, _13209_);
  or (_32728_, _32727_, _32717_);
  or (_32730_, _32728_, _06954_);
  and (_32731_, _07694_, \oc8051_golden_model_1.ACC [0]);
  or (_32732_, _32731_, _32717_);
  and (_32733_, _32732_, _06938_);
  nor (_32734_, _06938_, _32714_);
  or (_32735_, _32734_, _06102_);
  or (_32736_, _32735_, _32733_);
  and (_32737_, _32736_, _06044_);
  and (_32738_, _32737_, _32730_);
  nor (_32739_, _08357_, _32714_);
  and (_32741_, _14102_, _08357_);
  or (_32742_, _32741_, _32739_);
  and (_32743_, _32742_, _06043_);
  or (_32744_, _32743_, _32738_);
  and (_32745_, _32744_, _06848_);
  and (_32746_, _07694_, _06931_);
  or (_32747_, _32746_, _32717_);
  and (_32748_, _32747_, _06239_);
  or (_32749_, _32748_, _06219_);
  or (_32750_, _32749_, _32745_);
  or (_32752_, _32732_, _06220_);
  and (_32753_, _32752_, _06040_);
  and (_32754_, _32753_, _32750_);
  and (_32755_, _32717_, _06039_);
  or (_32756_, _32755_, _06032_);
  or (_32757_, _32756_, _32754_);
  or (_32758_, _32728_, _06033_);
  and (_32759_, _32758_, _06027_);
  and (_32760_, _32759_, _32757_);
  or (_32761_, _32739_, _14131_);
  and (_32763_, _32761_, _06026_);
  and (_32764_, _32763_, _32742_);
  or (_32765_, _32764_, _09818_);
  or (_32766_, _32765_, _32760_);
  or (_32767_, _32747_, _09827_);
  and (_32768_, _32767_, _05669_);
  and (_32769_, _32768_, _32766_);
  and (_32770_, _32769_, _32726_);
  and (_32771_, _14186_, _07694_);
  or (_32772_, _32771_, _32717_);
  and (_32774_, _32772_, _09833_);
  or (_32775_, _32774_, _06019_);
  or (_32776_, _32775_, _32770_);
  and (_32777_, _32776_, _32723_);
  or (_32778_, _32777_, _06112_);
  and (_32779_, _14086_, _07694_);
  or (_32780_, _32717_, _08751_);
  or (_32781_, _32780_, _32779_);
  and (_32782_, _32781_, _08756_);
  and (_32783_, _32782_, _32778_);
  nor (_32785_, _12302_, _13209_);
  or (_32786_, _32785_, _32717_);
  and (_32787_, _32716_, _06284_);
  and (_32788_, _32787_, _32786_);
  or (_32789_, _32788_, _32783_);
  and (_32790_, _32789_, _07032_);
  nand (_32791_, _32722_, _06108_);
  nor (_32792_, _32791_, _32727_);
  or (_32793_, _32792_, _06277_);
  or (_32794_, _32793_, _32790_);
  and (_32796_, _32794_, _32720_);
  or (_32797_, _32796_, _06130_);
  and (_32798_, _14083_, _07694_);
  or (_32799_, _32717_, _08777_);
  or (_32800_, _32799_, _32798_);
  and (_32801_, _32800_, _08782_);
  and (_32802_, _32801_, _32797_);
  and (_32803_, _32786_, _06292_);
  or (_32804_, _32803_, _06316_);
  or (_32805_, _32804_, _32802_);
  or (_32807_, _32728_, _06718_);
  and (_32808_, _32807_, _32805_);
  or (_32809_, _32808_, _05652_);
  or (_32810_, _32717_, _05653_);
  and (_32811_, _32810_, _32809_);
  or (_32812_, _32811_, _06047_);
  or (_32813_, _32728_, _06048_);
  and (_32814_, _32813_, _01336_);
  and (_32815_, _32814_, _32812_);
  or (_32816_, _32815_, _32715_);
  and (_43468_, _32816_, _42882_);
  not (_32818_, \oc8051_golden_model_1.IP [1]);
  nor (_32819_, _01336_, _32818_);
  nor (_32820_, _07694_, _32818_);
  nor (_32821_, _10993_, _13209_);
  or (_32822_, _32821_, _32820_);
  or (_32823_, _32822_, _08782_);
  or (_32824_, _14367_, _13209_);
  or (_32825_, _07694_, \oc8051_golden_model_1.IP [1]);
  and (_32826_, _32825_, _09833_);
  and (_32828_, _32826_, _32824_);
  nor (_32829_, _13209_, _07132_);
  or (_32830_, _32829_, _32820_);
  and (_32831_, _32830_, _06239_);
  nor (_32832_, _08357_, _32818_);
  and (_32833_, _14266_, _08357_);
  or (_32834_, _32833_, _32832_);
  or (_32835_, _32834_, _06044_);
  and (_32836_, _14284_, _07694_);
  not (_32837_, _32836_);
  and (_32839_, _32837_, _32825_);
  and (_32840_, _32839_, _06102_);
  nor (_32841_, _06938_, _32818_);
  and (_32842_, _07694_, \oc8051_golden_model_1.ACC [1]);
  or (_32843_, _32842_, _32820_);
  and (_32844_, _32843_, _06938_);
  or (_32845_, _32844_, _32841_);
  and (_32846_, _32845_, _06954_);
  or (_32847_, _32846_, _06043_);
  or (_32848_, _32847_, _32840_);
  and (_32850_, _32848_, _32835_);
  and (_32851_, _32850_, _06848_);
  or (_32852_, _32851_, _32831_);
  or (_32853_, _32852_, _06219_);
  or (_32854_, _32843_, _06220_);
  and (_32855_, _32854_, _06040_);
  and (_32856_, _32855_, _32853_);
  and (_32857_, _14273_, _08357_);
  or (_32858_, _32857_, _32832_);
  and (_32859_, _32858_, _06039_);
  or (_32861_, _32859_, _06032_);
  or (_32862_, _32861_, _32856_);
  or (_32863_, _32832_, _14302_);
  and (_32864_, _32863_, _32834_);
  or (_32865_, _32864_, _06033_);
  and (_32866_, _32865_, _06027_);
  and (_32867_, _32866_, _32862_);
  or (_32868_, _32832_, _14267_);
  and (_32869_, _32868_, _06026_);
  and (_32870_, _32869_, _32834_);
  or (_32872_, _32870_, _09815_);
  or (_32873_, _32872_, _32867_);
  or (_32874_, _32830_, _09827_);
  and (_32875_, _32874_, _32873_);
  or (_32876_, _32875_, _07011_);
  and (_32877_, _09075_, _07694_);
  or (_32878_, _32820_, _07012_);
  or (_32879_, _32878_, _32877_);
  and (_32880_, _32879_, _05669_);
  and (_32881_, _32880_, _32876_);
  or (_32883_, _32881_, _32828_);
  and (_32884_, _32883_, _06020_);
  nand (_32885_, _07694_, _06832_);
  and (_32886_, _32825_, _06019_);
  and (_32887_, _32886_, _32885_);
  or (_32888_, _32887_, _32884_);
  and (_32889_, _32888_, _08751_);
  or (_32890_, _14263_, _13209_);
  and (_32891_, _32825_, _06112_);
  and (_32892_, _32891_, _32890_);
  or (_32894_, _32892_, _06284_);
  or (_32895_, _32894_, _32889_);
  nand (_32896_, _10992_, _07694_);
  and (_32897_, _32896_, _32822_);
  or (_32898_, _32897_, _08756_);
  and (_32899_, _32898_, _07032_);
  and (_32900_, _32899_, _32895_);
  or (_32901_, _14261_, _13209_);
  and (_32902_, _32825_, _06108_);
  and (_32903_, _32902_, _32901_);
  or (_32905_, _32903_, _06277_);
  or (_32906_, _32905_, _32900_);
  nor (_32907_, _32820_, _06278_);
  nand (_32908_, _32907_, _32896_);
  and (_32909_, _32908_, _08777_);
  and (_32910_, _32909_, _32906_);
  or (_32911_, _32885_, _08078_);
  and (_32912_, _32825_, _06130_);
  and (_32913_, _32912_, _32911_);
  or (_32914_, _32913_, _06292_);
  or (_32916_, _32914_, _32910_);
  and (_32917_, _32916_, _32823_);
  or (_32918_, _32917_, _06316_);
  or (_32919_, _32839_, _06718_);
  and (_32920_, _32919_, _05653_);
  and (_32921_, _32920_, _32918_);
  and (_32922_, _32858_, _05652_);
  or (_32923_, _32922_, _06047_);
  or (_32924_, _32923_, _32921_);
  or (_32925_, _32820_, _06048_);
  or (_32927_, _32925_, _32836_);
  and (_32928_, _32927_, _01336_);
  and (_32929_, _32928_, _32924_);
  or (_32930_, _32929_, _32819_);
  and (_43469_, _32930_, _42882_);
  and (_32931_, _01340_, \oc8051_golden_model_1.IP [2]);
  and (_32932_, _13209_, \oc8051_golden_model_1.IP [2]);
  or (_32933_, _32932_, _08177_);
  and (_32934_, _07694_, _08730_);
  or (_32935_, _32934_, _32932_);
  and (_32937_, _32935_, _06108_);
  and (_32938_, _32937_, _32933_);
  or (_32939_, _32935_, _06020_);
  nor (_32940_, _13209_, _07530_);
  or (_32941_, _32940_, _32932_);
  or (_32942_, _32941_, _06848_);
  and (_32943_, _14493_, _07694_);
  or (_32944_, _32943_, _32932_);
  or (_32945_, _32944_, _06954_);
  and (_32946_, _07694_, \oc8051_golden_model_1.ACC [2]);
  or (_32948_, _32946_, _32932_);
  and (_32949_, _32948_, _06938_);
  and (_32950_, _06939_, \oc8051_golden_model_1.IP [2]);
  or (_32951_, _32950_, _06102_);
  or (_32952_, _32951_, _32949_);
  and (_32953_, _32952_, _06044_);
  and (_32954_, _32953_, _32945_);
  and (_32955_, _13228_, \oc8051_golden_model_1.IP [2]);
  and (_32956_, _14497_, _08357_);
  or (_32957_, _32956_, _32955_);
  and (_32959_, _32957_, _06043_);
  or (_32960_, _32959_, _06239_);
  or (_32961_, _32960_, _32954_);
  and (_32962_, _32961_, _32942_);
  or (_32963_, _32962_, _06219_);
  or (_32964_, _32948_, _06220_);
  and (_32965_, _32964_, _06040_);
  and (_32966_, _32965_, _32963_);
  and (_32967_, _14479_, _08357_);
  or (_32968_, _32967_, _32955_);
  and (_32970_, _32968_, _06039_);
  or (_32971_, _32970_, _06032_);
  or (_32972_, _32971_, _32966_);
  and (_32973_, _32956_, _14512_);
  or (_32974_, _32955_, _06033_);
  or (_32975_, _32974_, _32973_);
  and (_32976_, _32975_, _06027_);
  and (_32977_, _32976_, _32972_);
  or (_32978_, _32955_, _14525_);
  and (_32979_, _32978_, _06026_);
  and (_32981_, _32979_, _32957_);
  or (_32982_, _32981_, _09818_);
  or (_32983_, _32982_, _32977_);
  and (_32984_, _09182_, _07694_);
  or (_32985_, _32932_, _07012_);
  or (_32986_, _32985_, _32984_);
  or (_32987_, _32941_, _09827_);
  and (_32988_, _32987_, _05669_);
  and (_32989_, _32988_, _32986_);
  and (_32990_, _32989_, _32983_);
  and (_32992_, _14580_, _07694_);
  or (_32993_, _32992_, _32932_);
  and (_32994_, _32993_, _09833_);
  or (_32995_, _32994_, _06019_);
  or (_32996_, _32995_, _32990_);
  and (_32997_, _32996_, _32939_);
  or (_32998_, _32997_, _06112_);
  and (_32999_, _14596_, _07694_);
  or (_33000_, _32932_, _08751_);
  or (_33001_, _33000_, _32999_);
  and (_33003_, _33001_, _08756_);
  and (_33004_, _33003_, _32998_);
  and (_33005_, _10991_, _07694_);
  or (_33006_, _33005_, _32932_);
  and (_33007_, _33006_, _06284_);
  or (_33008_, _33007_, _33004_);
  and (_33009_, _33008_, _07032_);
  or (_33010_, _33009_, _32938_);
  and (_33011_, _33010_, _06278_);
  and (_33012_, _32948_, _06277_);
  and (_33014_, _33012_, _32933_);
  or (_33015_, _33014_, _06130_);
  or (_33016_, _33015_, _33011_);
  and (_33017_, _14593_, _07694_);
  or (_33018_, _32932_, _08777_);
  or (_33019_, _33018_, _33017_);
  and (_33020_, _33019_, _08782_);
  and (_33021_, _33020_, _33016_);
  nor (_33022_, _10990_, _13209_);
  or (_33023_, _33022_, _32932_);
  and (_33025_, _33023_, _06292_);
  or (_33026_, _33025_, _06316_);
  or (_33027_, _33026_, _33021_);
  or (_33028_, _32944_, _06718_);
  and (_33029_, _33028_, _05653_);
  and (_33030_, _33029_, _33027_);
  and (_33031_, _32968_, _05652_);
  or (_33032_, _33031_, _06047_);
  or (_33033_, _33032_, _33030_);
  and (_33034_, _14657_, _07694_);
  or (_33036_, _32932_, _06048_);
  or (_33037_, _33036_, _33034_);
  and (_33038_, _33037_, _01336_);
  and (_33039_, _33038_, _33033_);
  or (_33040_, _33039_, _32931_);
  and (_43470_, _33040_, _42882_);
  and (_33041_, _01340_, \oc8051_golden_model_1.IP [3]);
  and (_33042_, _13209_, \oc8051_golden_model_1.IP [3]);
  and (_33043_, _07694_, _08662_);
  or (_33044_, _33043_, _33042_);
  or (_33046_, _33044_, _06020_);
  and (_33047_, _14672_, _07694_);
  or (_33048_, _33047_, _33042_);
  or (_33049_, _33048_, _06954_);
  and (_33050_, _07694_, \oc8051_golden_model_1.ACC [3]);
  or (_33051_, _33050_, _33042_);
  and (_33052_, _33051_, _06938_);
  and (_33053_, _06939_, \oc8051_golden_model_1.IP [3]);
  or (_33054_, _33053_, _06102_);
  or (_33055_, _33054_, _33052_);
  and (_33057_, _33055_, _06044_);
  and (_33058_, _33057_, _33049_);
  and (_33059_, _13228_, \oc8051_golden_model_1.IP [3]);
  and (_33060_, _14683_, _08357_);
  or (_33061_, _33060_, _33059_);
  and (_33062_, _33061_, _06043_);
  or (_33063_, _33062_, _06239_);
  or (_33064_, _33063_, _33058_);
  nor (_33065_, _13209_, _07353_);
  or (_33066_, _33065_, _33042_);
  or (_33068_, _33066_, _06848_);
  and (_33069_, _33068_, _33064_);
  or (_33070_, _33069_, _06219_);
  or (_33071_, _33051_, _06220_);
  and (_33072_, _33071_, _06040_);
  and (_33073_, _33072_, _33070_);
  and (_33074_, _14681_, _08357_);
  or (_33075_, _33074_, _33059_);
  and (_33076_, _33075_, _06039_);
  or (_33077_, _33076_, _06032_);
  or (_33079_, _33077_, _33073_);
  or (_33080_, _33059_, _14708_);
  and (_33081_, _33080_, _33061_);
  or (_33082_, _33081_, _06033_);
  and (_33083_, _33082_, _06027_);
  and (_33084_, _33083_, _33079_);
  and (_33085_, _14724_, _08357_);
  or (_33086_, _33085_, _33059_);
  and (_33087_, _33086_, _06026_);
  or (_33088_, _33087_, _09818_);
  or (_33090_, _33088_, _33084_);
  and (_33091_, _09181_, _07694_);
  or (_33092_, _33042_, _07012_);
  or (_33093_, _33092_, _33091_);
  or (_33094_, _33066_, _09827_);
  and (_33095_, _33094_, _05669_);
  and (_33096_, _33095_, _33093_);
  and (_33097_, _33096_, _33090_);
  and (_33098_, _14778_, _07694_);
  or (_33099_, _33098_, _33042_);
  and (_33101_, _33099_, _09833_);
  or (_33102_, _33101_, _06019_);
  or (_33103_, _33102_, _33097_);
  and (_33104_, _33103_, _33046_);
  or (_33105_, _33104_, _06112_);
  and (_33106_, _14793_, _07694_);
  or (_33107_, _33042_, _08751_);
  or (_33108_, _33107_, _33106_);
  and (_33109_, _33108_, _08756_);
  and (_33110_, _33109_, _33105_);
  and (_33112_, _12299_, _07694_);
  or (_33113_, _33112_, _33042_);
  and (_33114_, _33113_, _06284_);
  or (_33115_, _33114_, _33110_);
  and (_33116_, _33115_, _07032_);
  or (_33117_, _33042_, _08029_);
  and (_33118_, _33044_, _06108_);
  and (_33119_, _33118_, _33117_);
  or (_33120_, _33119_, _33116_);
  and (_33121_, _33120_, _06278_);
  and (_33123_, _33051_, _06277_);
  and (_33124_, _33123_, _33117_);
  or (_33125_, _33124_, _06130_);
  or (_33126_, _33125_, _33121_);
  and (_33127_, _14792_, _07694_);
  or (_33128_, _33042_, _08777_);
  or (_33129_, _33128_, _33127_);
  and (_33130_, _33129_, _08782_);
  and (_33131_, _33130_, _33126_);
  nor (_33132_, _10988_, _13209_);
  or (_33134_, _33132_, _33042_);
  and (_33135_, _33134_, _06292_);
  or (_33136_, _33135_, _06316_);
  or (_33137_, _33136_, _33131_);
  or (_33138_, _33048_, _06718_);
  and (_33139_, _33138_, _05653_);
  and (_33140_, _33139_, _33137_);
  and (_33141_, _33075_, _05652_);
  or (_33142_, _33141_, _06047_);
  or (_33143_, _33142_, _33140_);
  and (_33145_, _14849_, _07694_);
  or (_33146_, _33042_, _06048_);
  or (_33147_, _33146_, _33145_);
  and (_33148_, _33147_, _01336_);
  and (_33149_, _33148_, _33143_);
  or (_33150_, _33149_, _33041_);
  and (_43471_, _33150_, _42882_);
  and (_33151_, _01340_, \oc8051_golden_model_1.IP [4]);
  and (_33152_, _13209_, \oc8051_golden_model_1.IP [4]);
  and (_33153_, _08665_, _07694_);
  or (_33155_, _33153_, _33152_);
  or (_33156_, _33155_, _06020_);
  and (_33157_, _14887_, _07694_);
  or (_33158_, _33157_, _33152_);
  or (_33159_, _33158_, _06954_);
  and (_33160_, _07694_, \oc8051_golden_model_1.ACC [4]);
  or (_33161_, _33160_, _33152_);
  and (_33162_, _33161_, _06938_);
  and (_33163_, _06939_, \oc8051_golden_model_1.IP [4]);
  or (_33164_, _33163_, _06102_);
  or (_33166_, _33164_, _33162_);
  and (_33167_, _33166_, _06044_);
  and (_33168_, _33167_, _33159_);
  and (_33169_, _13228_, \oc8051_golden_model_1.IP [4]);
  and (_33170_, _14878_, _08357_);
  or (_33171_, _33170_, _33169_);
  and (_33172_, _33171_, _06043_);
  or (_33173_, _33172_, _06239_);
  or (_33174_, _33173_, _33168_);
  nor (_33175_, _08270_, _13209_);
  or (_33177_, _33175_, _33152_);
  or (_33178_, _33177_, _06848_);
  and (_33179_, _33178_, _33174_);
  or (_33180_, _33179_, _06219_);
  or (_33181_, _33161_, _06220_);
  and (_33182_, _33181_, _06040_);
  and (_33183_, _33182_, _33180_);
  and (_33184_, _14882_, _08357_);
  or (_33185_, _33184_, _33169_);
  and (_33186_, _33185_, _06039_);
  or (_33188_, _33186_, _06032_);
  or (_33189_, _33188_, _33183_);
  or (_33190_, _33169_, _14914_);
  and (_33191_, _33190_, _33171_);
  or (_33192_, _33191_, _06033_);
  and (_33193_, _33192_, _06027_);
  and (_33194_, _33193_, _33189_);
  or (_33195_, _33169_, _14879_);
  and (_33196_, _33195_, _06026_);
  and (_33197_, _33196_, _33171_);
  or (_33199_, _33197_, _09818_);
  or (_33200_, _33199_, _33194_);
  and (_33201_, _09180_, _07694_);
  or (_33202_, _33152_, _07012_);
  or (_33203_, _33202_, _33201_);
  or (_33204_, _33177_, _09827_);
  and (_33205_, _33204_, _05669_);
  and (_33206_, _33205_, _33203_);
  and (_33207_, _33206_, _33200_);
  and (_33208_, _14983_, _07694_);
  or (_33210_, _33208_, _33152_);
  and (_33211_, _33210_, _09833_);
  or (_33212_, _33211_, _06019_);
  or (_33213_, _33212_, _33207_);
  and (_33214_, _33213_, _33156_);
  or (_33215_, _33214_, _06112_);
  and (_33216_, _14876_, _07694_);
  or (_33217_, _33216_, _33152_);
  or (_33218_, _33217_, _08751_);
  and (_33219_, _33218_, _08756_);
  and (_33221_, _33219_, _33215_);
  and (_33222_, _10986_, _07694_);
  or (_33223_, _33222_, _33152_);
  and (_33224_, _33223_, _06284_);
  or (_33225_, _33224_, _33221_);
  and (_33226_, _33225_, _07032_);
  or (_33227_, _33152_, _08273_);
  and (_33228_, _33155_, _06108_);
  and (_33229_, _33228_, _33227_);
  or (_33230_, _33229_, _33226_);
  and (_33232_, _33230_, _06278_);
  and (_33233_, _33161_, _06277_);
  and (_33234_, _33233_, _33227_);
  or (_33235_, _33234_, _06130_);
  or (_33236_, _33235_, _33232_);
  and (_33237_, _14873_, _07694_);
  or (_33238_, _33152_, _08777_);
  or (_33239_, _33238_, _33237_);
  and (_33240_, _33239_, _08782_);
  and (_33241_, _33240_, _33236_);
  nor (_33243_, _10985_, _13209_);
  or (_33244_, _33243_, _33152_);
  and (_33245_, _33244_, _06292_);
  or (_33246_, _33245_, _06316_);
  or (_33247_, _33246_, _33241_);
  or (_33248_, _33158_, _06718_);
  and (_33249_, _33248_, _05653_);
  and (_33250_, _33249_, _33247_);
  and (_33251_, _33185_, _05652_);
  or (_33252_, _33251_, _06047_);
  or (_33254_, _33252_, _33250_);
  and (_33255_, _15055_, _07694_);
  or (_33256_, _33152_, _06048_);
  or (_33257_, _33256_, _33255_);
  and (_33258_, _33257_, _01336_);
  and (_33259_, _33258_, _33254_);
  or (_33260_, _33259_, _33151_);
  and (_43472_, _33260_, _42882_);
  and (_33261_, _01340_, \oc8051_golden_model_1.IP [5]);
  and (_33262_, _13209_, \oc8051_golden_model_1.IP [5]);
  and (_33264_, _08652_, _07694_);
  or (_33265_, _33264_, _33262_);
  or (_33266_, _33265_, _06020_);
  and (_33267_, _15093_, _07694_);
  or (_33268_, _33267_, _33262_);
  or (_33269_, _33268_, _06954_);
  and (_33270_, _07694_, \oc8051_golden_model_1.ACC [5]);
  or (_33271_, _33270_, _33262_);
  and (_33272_, _33271_, _06938_);
  and (_33273_, _06939_, \oc8051_golden_model_1.IP [5]);
  or (_33275_, _33273_, _06102_);
  or (_33276_, _33275_, _33272_);
  and (_33277_, _33276_, _06044_);
  and (_33278_, _33277_, _33269_);
  and (_33279_, _13228_, \oc8051_golden_model_1.IP [5]);
  and (_33280_, _15073_, _08357_);
  or (_33281_, _33280_, _33279_);
  and (_33282_, _33281_, _06043_);
  or (_33283_, _33282_, _06239_);
  or (_33284_, _33283_, _33278_);
  nor (_33286_, _07977_, _13209_);
  or (_33287_, _33286_, _33262_);
  or (_33288_, _33287_, _06848_);
  and (_33289_, _33288_, _33284_);
  or (_33290_, _33289_, _06219_);
  or (_33291_, _33271_, _06220_);
  and (_33292_, _33291_, _06040_);
  and (_33293_, _33292_, _33290_);
  and (_33294_, _15077_, _08357_);
  or (_33295_, _33294_, _33279_);
  and (_33297_, _33295_, _06039_);
  or (_33298_, _33297_, _06032_);
  or (_33299_, _33298_, _33293_);
  or (_33300_, _33279_, _15110_);
  and (_33301_, _33300_, _33281_);
  or (_33302_, _33301_, _06033_);
  and (_33303_, _33302_, _06027_);
  and (_33304_, _33303_, _33299_);
  or (_33305_, _33279_, _15074_);
  and (_33306_, _33305_, _06026_);
  and (_33308_, _33306_, _33281_);
  or (_33309_, _33308_, _09818_);
  or (_33310_, _33309_, _33304_);
  and (_33311_, _09179_, _07694_);
  or (_33312_, _33262_, _07012_);
  or (_33313_, _33312_, _33311_);
  or (_33314_, _33287_, _09827_);
  and (_33315_, _33314_, _05669_);
  and (_33316_, _33315_, _33313_);
  and (_33317_, _33316_, _33310_);
  and (_33319_, _15179_, _07694_);
  or (_33320_, _33319_, _33262_);
  and (_33321_, _33320_, _09833_);
  or (_33322_, _33321_, _06019_);
  or (_33323_, _33322_, _33317_);
  and (_33324_, _33323_, _33266_);
  or (_33325_, _33324_, _06112_);
  and (_33326_, _15195_, _07694_);
  or (_33327_, _33262_, _08751_);
  or (_33328_, _33327_, _33326_);
  and (_33330_, _33328_, _08756_);
  and (_33331_, _33330_, _33325_);
  and (_33332_, _12306_, _07694_);
  or (_33333_, _33332_, _33262_);
  and (_33334_, _33333_, _06284_);
  or (_33335_, _33334_, _33331_);
  and (_33336_, _33335_, _07032_);
  or (_33337_, _33262_, _07980_);
  and (_33338_, _33265_, _06108_);
  and (_33339_, _33338_, _33337_);
  or (_33341_, _33339_, _33336_);
  and (_33342_, _33341_, _06278_);
  and (_33343_, _33271_, _06277_);
  and (_33344_, _33343_, _33337_);
  or (_33345_, _33344_, _06130_);
  or (_33346_, _33345_, _33342_);
  and (_33347_, _15194_, _07694_);
  or (_33348_, _33262_, _08777_);
  or (_33349_, _33348_, _33347_);
  and (_33350_, _33349_, _08782_);
  and (_33352_, _33350_, _33346_);
  nor (_33353_, _10982_, _13209_);
  or (_33354_, _33353_, _33262_);
  and (_33355_, _33354_, _06292_);
  or (_33356_, _33355_, _06316_);
  or (_33357_, _33356_, _33352_);
  or (_33358_, _33268_, _06718_);
  and (_33359_, _33358_, _05653_);
  and (_33360_, _33359_, _33357_);
  and (_33361_, _33295_, _05652_);
  or (_33363_, _33361_, _06047_);
  or (_33364_, _33363_, _33360_);
  and (_33365_, _15253_, _07694_);
  or (_33366_, _33262_, _06048_);
  or (_33367_, _33366_, _33365_);
  and (_33368_, _33367_, _01336_);
  and (_33369_, _33368_, _33364_);
  or (_33370_, _33369_, _33261_);
  and (_43473_, _33370_, _42882_);
  and (_33371_, _01340_, \oc8051_golden_model_1.IP [6]);
  and (_33373_, _13209_, \oc8051_golden_model_1.IP [6]);
  and (_33374_, _15389_, _07694_);
  or (_33375_, _33374_, _33373_);
  or (_33376_, _33375_, _06020_);
  and (_33377_, _15293_, _07694_);
  or (_33378_, _33377_, _33373_);
  or (_33379_, _33378_, _06954_);
  and (_33380_, _07694_, \oc8051_golden_model_1.ACC [6]);
  or (_33381_, _33380_, _33373_);
  and (_33382_, _33381_, _06938_);
  and (_33384_, _06939_, \oc8051_golden_model_1.IP [6]);
  or (_33385_, _33384_, _06102_);
  or (_33386_, _33385_, _33382_);
  and (_33387_, _33386_, _06044_);
  and (_33388_, _33387_, _33379_);
  and (_33389_, _13228_, \oc8051_golden_model_1.IP [6]);
  and (_33390_, _15280_, _08357_);
  or (_33391_, _33390_, _33389_);
  and (_33392_, _33391_, _06043_);
  or (_33393_, _33392_, _06239_);
  or (_33395_, _33393_, _33388_);
  nor (_33396_, _07883_, _13209_);
  or (_33397_, _33396_, _33373_);
  or (_33398_, _33397_, _06848_);
  and (_33399_, _33398_, _33395_);
  or (_33400_, _33399_, _06219_);
  or (_33401_, _33381_, _06220_);
  and (_33402_, _33401_, _06040_);
  and (_33403_, _33402_, _33400_);
  and (_33404_, _15278_, _08357_);
  or (_33406_, _33404_, _33389_);
  and (_33407_, _33406_, _06039_);
  or (_33408_, _33407_, _06032_);
  or (_33409_, _33408_, _33403_);
  or (_33410_, _33389_, _15310_);
  and (_33411_, _33410_, _33391_);
  or (_33412_, _33411_, _06033_);
  and (_33413_, _33412_, _06027_);
  and (_33414_, _33413_, _33409_);
  or (_33415_, _33389_, _15326_);
  and (_33416_, _33415_, _06026_);
  and (_33417_, _33416_, _33391_);
  or (_33418_, _33417_, _09818_);
  or (_33419_, _33418_, _33414_);
  and (_33420_, _09178_, _07694_);
  or (_33421_, _33373_, _07012_);
  or (_33422_, _33421_, _33420_);
  or (_33423_, _33397_, _09827_);
  and (_33424_, _33423_, _05669_);
  and (_33425_, _33424_, _33422_);
  and (_33427_, _33425_, _33419_);
  and (_33428_, _15382_, _07694_);
  or (_33429_, _33428_, _33373_);
  and (_33430_, _33429_, _09833_);
  or (_33431_, _33430_, _06019_);
  or (_33432_, _33431_, _33427_);
  and (_33433_, _33432_, _33376_);
  or (_33434_, _33433_, _06112_);
  and (_33435_, _15399_, _07694_);
  or (_33436_, _33435_, _33373_);
  or (_33438_, _33436_, _08751_);
  and (_33439_, _33438_, _08756_);
  and (_33440_, _33439_, _33434_);
  and (_33441_, _10980_, _07694_);
  or (_33442_, _33441_, _33373_);
  and (_33443_, _33442_, _06284_);
  or (_33444_, _33443_, _33440_);
  and (_33445_, _33444_, _07032_);
  or (_33446_, _33373_, _07886_);
  and (_33447_, _33375_, _06108_);
  and (_33449_, _33447_, _33446_);
  or (_33450_, _33449_, _33445_);
  and (_33451_, _33450_, _06278_);
  and (_33452_, _33381_, _06277_);
  and (_33453_, _33452_, _33446_);
  or (_33454_, _33453_, _06130_);
  or (_33455_, _33454_, _33451_);
  and (_33456_, _15396_, _07694_);
  or (_33457_, _33373_, _08777_);
  or (_33458_, _33457_, _33456_);
  and (_33460_, _33458_, _08782_);
  and (_33461_, _33460_, _33455_);
  nor (_33462_, _10979_, _13209_);
  or (_33463_, _33462_, _33373_);
  and (_33464_, _33463_, _06292_);
  or (_33465_, _33464_, _06316_);
  or (_33466_, _33465_, _33461_);
  or (_33467_, _33378_, _06718_);
  and (_33468_, _33467_, _05653_);
  and (_33469_, _33468_, _33466_);
  and (_33471_, _33406_, _05652_);
  or (_33472_, _33471_, _06047_);
  or (_33473_, _33472_, _33469_);
  and (_33474_, _15451_, _07694_);
  or (_33475_, _33373_, _06048_);
  or (_33476_, _33475_, _33474_);
  and (_33477_, _33476_, _01336_);
  and (_33478_, _33477_, _33473_);
  or (_33479_, _33478_, _33371_);
  and (_43474_, _33479_, _42882_);
  not (_33481_, \oc8051_golden_model_1.IE [0]);
  nor (_33482_, _01336_, _33481_);
  nor (_33483_, _07688_, _33481_);
  and (_33484_, _07688_, _08672_);
  or (_33485_, _33484_, _33483_);
  or (_33486_, _33485_, _06020_);
  and (_33487_, _09120_, _07688_);
  or (_33488_, _33483_, _07012_);
  or (_33489_, _33488_, _33487_);
  nor (_33490_, _08127_, _13311_);
  or (_33492_, _33490_, _33483_);
  or (_33493_, _33492_, _06954_);
  and (_33494_, _07688_, \oc8051_golden_model_1.ACC [0]);
  or (_33495_, _33494_, _33483_);
  and (_33496_, _33495_, _06938_);
  nor (_33497_, _06938_, _33481_);
  or (_33498_, _33497_, _06102_);
  or (_33499_, _33498_, _33496_);
  and (_33500_, _33499_, _06044_);
  and (_33501_, _33500_, _33493_);
  nor (_33503_, _08351_, _33481_);
  and (_33504_, _14102_, _08351_);
  or (_33505_, _33504_, _33503_);
  and (_33506_, _33505_, _06043_);
  or (_33507_, _33506_, _33501_);
  and (_33508_, _33507_, _06848_);
  and (_33509_, _07688_, _06931_);
  or (_33510_, _33509_, _33483_);
  and (_33511_, _33510_, _06239_);
  or (_33512_, _33511_, _06219_);
  or (_33514_, _33512_, _33508_);
  or (_33515_, _33495_, _06220_);
  and (_33516_, _33515_, _06040_);
  and (_33517_, _33516_, _33514_);
  and (_33518_, _33483_, _06039_);
  or (_33519_, _33518_, _06032_);
  or (_33520_, _33519_, _33517_);
  or (_33521_, _33492_, _06033_);
  and (_33522_, _33521_, _06027_);
  and (_33523_, _33522_, _33520_);
  or (_33525_, _33503_, _14131_);
  and (_33526_, _33525_, _06026_);
  and (_33527_, _33526_, _33505_);
  or (_33528_, _33527_, _09818_);
  or (_33529_, _33528_, _33523_);
  or (_33530_, _33510_, _09827_);
  and (_33531_, _33530_, _05669_);
  and (_33532_, _33531_, _33529_);
  and (_33533_, _33532_, _33489_);
  and (_33534_, _14186_, _07688_);
  or (_33536_, _33534_, _33483_);
  and (_33537_, _33536_, _09833_);
  or (_33538_, _33537_, _06019_);
  or (_33539_, _33538_, _33533_);
  and (_33540_, _33539_, _33486_);
  or (_33541_, _33540_, _06112_);
  and (_33542_, _14086_, _07688_);
  or (_33543_, _33483_, _08751_);
  or (_33544_, _33543_, _33542_);
  and (_33545_, _33544_, _08756_);
  and (_33547_, _33545_, _33541_);
  nor (_33548_, _12302_, _13311_);
  or (_33549_, _33548_, _33483_);
  nand (_33550_, _10995_, _07688_);
  and (_33551_, _33550_, _06284_);
  and (_33552_, _33551_, _33549_);
  or (_33553_, _33552_, _33547_);
  and (_33554_, _33553_, _07032_);
  nand (_33555_, _33485_, _06108_);
  nor (_33556_, _33555_, _33490_);
  or (_33558_, _33556_, _06277_);
  or (_33559_, _33558_, _33554_);
  nor (_33560_, _33483_, _06278_);
  nand (_33561_, _33560_, _33550_);
  and (_33562_, _33561_, _33559_);
  or (_33563_, _33562_, _06130_);
  and (_33564_, _14083_, _07688_);
  or (_33565_, _33483_, _08777_);
  or (_33566_, _33565_, _33564_);
  and (_33567_, _33566_, _08782_);
  and (_33569_, _33567_, _33563_);
  and (_33570_, _33549_, _06292_);
  or (_33571_, _33570_, _06316_);
  or (_33572_, _33571_, _33569_);
  or (_33573_, _33492_, _06718_);
  and (_33574_, _33573_, _33572_);
  or (_33575_, _33574_, _05652_);
  or (_33576_, _33483_, _05653_);
  and (_33577_, _33576_, _33575_);
  or (_33578_, _33577_, _06047_);
  or (_33580_, _33492_, _06048_);
  and (_33581_, _33580_, _01336_);
  and (_33582_, _33581_, _33578_);
  or (_33583_, _33582_, _33482_);
  and (_43476_, _33583_, _42882_);
  not (_33584_, \oc8051_golden_model_1.IE [1]);
  nor (_33585_, _01336_, _33584_);
  nor (_33586_, _07688_, _33584_);
  nor (_33587_, _10993_, _13311_);
  or (_33588_, _33587_, _33586_);
  or (_33590_, _33588_, _08782_);
  or (_33591_, _14367_, _13311_);
  or (_33592_, _07688_, \oc8051_golden_model_1.IE [1]);
  and (_33593_, _33592_, _09833_);
  and (_33594_, _33593_, _33591_);
  nor (_33595_, _13311_, _07132_);
  or (_33596_, _33595_, _33586_);
  or (_33597_, _33596_, _06848_);
  and (_33598_, _14284_, _07688_);
  not (_33599_, _33598_);
  and (_33601_, _33599_, _33592_);
  or (_33602_, _33601_, _06954_);
  and (_33603_, _07688_, \oc8051_golden_model_1.ACC [1]);
  or (_33604_, _33603_, _33586_);
  and (_33605_, _33604_, _06938_);
  nor (_33606_, _06938_, _33584_);
  or (_33607_, _33606_, _06102_);
  or (_33608_, _33607_, _33605_);
  and (_33609_, _33608_, _06044_);
  and (_33610_, _33609_, _33602_);
  nor (_33612_, _08351_, _33584_);
  and (_33613_, _14266_, _08351_);
  or (_33614_, _33613_, _33612_);
  and (_33615_, _33614_, _06043_);
  or (_33616_, _33615_, _06239_);
  or (_33617_, _33616_, _33610_);
  and (_33618_, _33617_, _33597_);
  or (_33619_, _33618_, _06219_);
  or (_33620_, _33604_, _06220_);
  and (_33621_, _33620_, _06040_);
  and (_33623_, _33621_, _33619_);
  and (_33624_, _14273_, _08351_);
  or (_33625_, _33624_, _33612_);
  and (_33626_, _33625_, _06039_);
  or (_33627_, _33626_, _06032_);
  or (_33628_, _33627_, _33623_);
  and (_33629_, _33613_, _14302_);
  or (_33630_, _33612_, _06033_);
  or (_33631_, _33630_, _33629_);
  and (_33632_, _33631_, _06027_);
  and (_33634_, _33632_, _33628_);
  or (_33635_, _33612_, _14267_);
  and (_33636_, _33635_, _06026_);
  and (_33637_, _33636_, _33614_);
  or (_33638_, _33637_, _09818_);
  or (_33639_, _33638_, _33634_);
  and (_33640_, _09075_, _07688_);
  or (_33641_, _33586_, _07012_);
  or (_33642_, _33641_, _33640_);
  or (_33643_, _33596_, _09827_);
  and (_33645_, _33643_, _05669_);
  and (_33646_, _33645_, _33642_);
  and (_33647_, _33646_, _33639_);
  or (_33648_, _33647_, _33594_);
  and (_33649_, _33648_, _06020_);
  nand (_33650_, _07688_, _06832_);
  and (_33651_, _33592_, _06019_);
  and (_33652_, _33651_, _33650_);
  or (_33653_, _33652_, _33649_);
  and (_33654_, _33653_, _08751_);
  or (_33656_, _14263_, _13311_);
  and (_33657_, _33592_, _06112_);
  and (_33658_, _33657_, _33656_);
  or (_33659_, _33658_, _06284_);
  or (_33660_, _33659_, _33654_);
  nand (_33661_, _10992_, _07688_);
  and (_33662_, _33661_, _33588_);
  or (_33663_, _33662_, _08756_);
  and (_33664_, _33663_, _07032_);
  and (_33665_, _33664_, _33660_);
  or (_33667_, _14261_, _13311_);
  and (_33668_, _33592_, _06108_);
  and (_33669_, _33668_, _33667_);
  or (_33670_, _33669_, _06277_);
  or (_33671_, _33670_, _33665_);
  nor (_33672_, _33586_, _06278_);
  nand (_33673_, _33672_, _33661_);
  and (_33674_, _33673_, _08777_);
  and (_33675_, _33674_, _33671_);
  or (_33676_, _33650_, _08078_);
  and (_33678_, _33592_, _06130_);
  and (_33679_, _33678_, _33676_);
  or (_33680_, _33679_, _06292_);
  or (_33681_, _33680_, _33675_);
  and (_33682_, _33681_, _33590_);
  or (_33683_, _33682_, _06316_);
  or (_33684_, _33601_, _06718_);
  and (_33685_, _33684_, _05653_);
  and (_33686_, _33685_, _33683_);
  and (_33687_, _33625_, _05652_);
  or (_33689_, _33687_, _06047_);
  or (_33690_, _33689_, _33686_);
  or (_33691_, _33586_, _06048_);
  or (_33692_, _33691_, _33598_);
  and (_33693_, _33692_, _01336_);
  and (_33694_, _33693_, _33690_);
  or (_33695_, _33694_, _33585_);
  and (_43477_, _33695_, _42882_);
  and (_33696_, _01340_, \oc8051_golden_model_1.IE [2]);
  and (_33697_, _13311_, \oc8051_golden_model_1.IE [2]);
  and (_33699_, _07688_, _08730_);
  or (_33700_, _33699_, _33697_);
  or (_33701_, _33700_, _06020_);
  nor (_33702_, _13311_, _07530_);
  or (_33703_, _33702_, _33697_);
  and (_33704_, _33703_, _06239_);
  and (_33705_, _13330_, \oc8051_golden_model_1.IE [2]);
  and (_33706_, _14497_, _08351_);
  or (_33707_, _33706_, _33705_);
  or (_33708_, _33707_, _06044_);
  and (_33710_, _14493_, _07688_);
  or (_33711_, _33710_, _33697_);
  and (_33712_, _33711_, _06102_);
  and (_33713_, _06939_, \oc8051_golden_model_1.IE [2]);
  and (_33714_, _07688_, \oc8051_golden_model_1.ACC [2]);
  or (_33715_, _33714_, _33697_);
  and (_33716_, _33715_, _06938_);
  or (_33717_, _33716_, _33713_);
  and (_33718_, _33717_, _06954_);
  or (_33719_, _33718_, _06043_);
  or (_33721_, _33719_, _33712_);
  and (_33722_, _33721_, _33708_);
  and (_33723_, _33722_, _06848_);
  or (_33724_, _33723_, _33704_);
  or (_33725_, _33724_, _06219_);
  or (_33726_, _33715_, _06220_);
  and (_33727_, _33726_, _06040_);
  and (_33728_, _33727_, _33725_);
  and (_33729_, _14479_, _08351_);
  or (_33730_, _33729_, _33705_);
  and (_33732_, _33730_, _06039_);
  or (_33733_, _33732_, _06032_);
  or (_33734_, _33733_, _33728_);
  or (_33735_, _33705_, _14512_);
  and (_33736_, _33735_, _33707_);
  or (_33737_, _33736_, _06033_);
  and (_33738_, _33737_, _06027_);
  and (_33739_, _33738_, _33734_);
  or (_33740_, _33705_, _14525_);
  and (_33741_, _33740_, _06026_);
  and (_33743_, _33741_, _33707_);
  or (_33744_, _33743_, _09818_);
  or (_33745_, _33744_, _33739_);
  and (_33746_, _09182_, _07688_);
  or (_33747_, _33697_, _07012_);
  or (_33748_, _33747_, _33746_);
  or (_33749_, _33703_, _09827_);
  and (_33750_, _33749_, _05669_);
  and (_33751_, _33750_, _33748_);
  and (_33752_, _33751_, _33745_);
  and (_33754_, _14580_, _07688_);
  or (_33755_, _33754_, _33697_);
  and (_33756_, _33755_, _09833_);
  or (_33757_, _33756_, _06019_);
  or (_33758_, _33757_, _33752_);
  and (_33759_, _33758_, _33701_);
  or (_33760_, _33759_, _06112_);
  and (_33761_, _14596_, _07688_);
  or (_33762_, _33697_, _08751_);
  or (_33763_, _33762_, _33761_);
  and (_33765_, _33763_, _08756_);
  and (_33766_, _33765_, _33760_);
  and (_33767_, _10991_, _07688_);
  or (_33768_, _33767_, _33697_);
  and (_33769_, _33768_, _06284_);
  or (_33770_, _33769_, _33766_);
  and (_33771_, _33770_, _07032_);
  or (_33772_, _33697_, _08177_);
  and (_33773_, _33700_, _06108_);
  and (_33774_, _33773_, _33772_);
  or (_33776_, _33774_, _33771_);
  and (_33777_, _33776_, _06278_);
  and (_33778_, _33715_, _06277_);
  and (_33779_, _33778_, _33772_);
  or (_33780_, _33779_, _06130_);
  or (_33781_, _33780_, _33777_);
  and (_33782_, _14593_, _07688_);
  or (_33783_, _33697_, _08777_);
  or (_33784_, _33783_, _33782_);
  and (_33785_, _33784_, _08782_);
  and (_33787_, _33785_, _33781_);
  nor (_33788_, _10990_, _13311_);
  or (_33789_, _33788_, _33697_);
  and (_33790_, _33789_, _06292_);
  or (_33791_, _33790_, _06316_);
  or (_33792_, _33791_, _33787_);
  or (_33793_, _33711_, _06718_);
  and (_33794_, _33793_, _05653_);
  and (_33795_, _33794_, _33792_);
  and (_33796_, _33730_, _05652_);
  or (_33798_, _33796_, _06047_);
  or (_33799_, _33798_, _33795_);
  and (_33800_, _14657_, _07688_);
  or (_33801_, _33697_, _06048_);
  or (_33802_, _33801_, _33800_);
  and (_33803_, _33802_, _01336_);
  and (_33804_, _33803_, _33799_);
  or (_33805_, _33804_, _33696_);
  and (_43478_, _33805_, _42882_);
  and (_33806_, _01340_, \oc8051_golden_model_1.IE [3]);
  and (_33808_, _13311_, \oc8051_golden_model_1.IE [3]);
  and (_33809_, _07688_, _08662_);
  or (_33810_, _33809_, _33808_);
  or (_33811_, _33810_, _06020_);
  and (_33812_, _14672_, _07688_);
  or (_33813_, _33812_, _33808_);
  or (_33814_, _33813_, _06954_);
  and (_33815_, _07688_, \oc8051_golden_model_1.ACC [3]);
  or (_33816_, _33815_, _33808_);
  and (_33817_, _33816_, _06938_);
  and (_33819_, _06939_, \oc8051_golden_model_1.IE [3]);
  or (_33820_, _33819_, _06102_);
  or (_33821_, _33820_, _33817_);
  and (_33822_, _33821_, _06044_);
  and (_33823_, _33822_, _33814_);
  and (_33824_, _13330_, \oc8051_golden_model_1.IE [3]);
  and (_33825_, _14683_, _08351_);
  or (_33826_, _33825_, _33824_);
  and (_33827_, _33826_, _06043_);
  or (_33828_, _33827_, _06239_);
  or (_33830_, _33828_, _33823_);
  nor (_33831_, _13311_, _07353_);
  or (_33832_, _33831_, _33808_);
  or (_33833_, _33832_, _06848_);
  and (_33834_, _33833_, _33830_);
  or (_33835_, _33834_, _06219_);
  or (_33836_, _33816_, _06220_);
  and (_33837_, _33836_, _06040_);
  and (_33838_, _33837_, _33835_);
  and (_33839_, _14681_, _08351_);
  or (_33841_, _33839_, _33824_);
  and (_33842_, _33841_, _06039_);
  or (_33843_, _33842_, _06032_);
  or (_33844_, _33843_, _33838_);
  or (_33845_, _33824_, _14708_);
  and (_33846_, _33845_, _33826_);
  or (_33847_, _33846_, _06033_);
  and (_33848_, _33847_, _06027_);
  and (_33849_, _33848_, _33844_);
  and (_33850_, _14724_, _08351_);
  or (_33852_, _33850_, _33824_);
  and (_33853_, _33852_, _06026_);
  or (_33854_, _33853_, _09818_);
  or (_33855_, _33854_, _33849_);
  and (_33856_, _09181_, _07688_);
  or (_33857_, _33808_, _07012_);
  or (_33858_, _33857_, _33856_);
  or (_33859_, _33832_, _09827_);
  and (_33860_, _33859_, _05669_);
  and (_33861_, _33860_, _33858_);
  and (_33863_, _33861_, _33855_);
  and (_33864_, _14778_, _07688_);
  or (_33865_, _33864_, _33808_);
  and (_33866_, _33865_, _09833_);
  or (_33867_, _33866_, _06019_);
  or (_33868_, _33867_, _33863_);
  and (_33869_, _33868_, _33811_);
  or (_33870_, _33869_, _06112_);
  and (_33871_, _14793_, _07688_);
  or (_33872_, _33808_, _08751_);
  or (_33874_, _33872_, _33871_);
  and (_33875_, _33874_, _08756_);
  and (_33876_, _33875_, _33870_);
  and (_33877_, _12299_, _07688_);
  or (_33878_, _33877_, _33808_);
  and (_33879_, _33878_, _06284_);
  or (_33880_, _33879_, _33876_);
  and (_33881_, _33880_, _07032_);
  or (_33882_, _33808_, _08029_);
  and (_33883_, _33810_, _06108_);
  and (_33885_, _33883_, _33882_);
  or (_33886_, _33885_, _33881_);
  and (_33887_, _33886_, _06278_);
  and (_33888_, _33816_, _06277_);
  and (_33889_, _33888_, _33882_);
  or (_33890_, _33889_, _06130_);
  or (_33891_, _33890_, _33887_);
  and (_33892_, _14792_, _07688_);
  or (_33893_, _33808_, _08777_);
  or (_33894_, _33893_, _33892_);
  and (_33896_, _33894_, _08782_);
  and (_33897_, _33896_, _33891_);
  nor (_33898_, _10988_, _13311_);
  or (_33899_, _33898_, _33808_);
  and (_33900_, _33899_, _06292_);
  or (_33901_, _33900_, _06316_);
  or (_33902_, _33901_, _33897_);
  or (_33903_, _33813_, _06718_);
  and (_33904_, _33903_, _05653_);
  and (_33905_, _33904_, _33902_);
  and (_33907_, _33841_, _05652_);
  or (_33908_, _33907_, _06047_);
  or (_33909_, _33908_, _33905_);
  and (_33910_, _14849_, _07688_);
  or (_33911_, _33808_, _06048_);
  or (_33912_, _33911_, _33910_);
  and (_33913_, _33912_, _01336_);
  and (_33914_, _33913_, _33909_);
  or (_33915_, _33914_, _33806_);
  and (_43479_, _33915_, _42882_);
  and (_33917_, _01340_, \oc8051_golden_model_1.IE [4]);
  and (_33918_, _13311_, \oc8051_golden_model_1.IE [4]);
  and (_33919_, _08665_, _07688_);
  or (_33920_, _33919_, _33918_);
  or (_33921_, _33920_, _06020_);
  and (_33922_, _14887_, _07688_);
  or (_33923_, _33922_, _33918_);
  or (_33924_, _33923_, _06954_);
  and (_33925_, _07688_, \oc8051_golden_model_1.ACC [4]);
  or (_33926_, _33925_, _33918_);
  and (_33928_, _33926_, _06938_);
  and (_33929_, _06939_, \oc8051_golden_model_1.IE [4]);
  or (_33930_, _33929_, _06102_);
  or (_33931_, _33930_, _33928_);
  and (_33932_, _33931_, _06044_);
  and (_33933_, _33932_, _33924_);
  and (_33934_, _13330_, \oc8051_golden_model_1.IE [4]);
  and (_33935_, _14878_, _08351_);
  or (_33936_, _33935_, _33934_);
  and (_33937_, _33936_, _06043_);
  or (_33939_, _33937_, _06239_);
  or (_33940_, _33939_, _33933_);
  nor (_33941_, _08270_, _13311_);
  or (_33942_, _33941_, _33918_);
  or (_33943_, _33942_, _06848_);
  and (_33944_, _33943_, _33940_);
  or (_33945_, _33944_, _06219_);
  or (_33946_, _33926_, _06220_);
  and (_33947_, _33946_, _06040_);
  and (_33948_, _33947_, _33945_);
  and (_33950_, _14882_, _08351_);
  or (_33951_, _33950_, _33934_);
  and (_33952_, _33951_, _06039_);
  or (_33953_, _33952_, _06032_);
  or (_33954_, _33953_, _33948_);
  or (_33955_, _33934_, _14914_);
  and (_33956_, _33955_, _33936_);
  or (_33957_, _33956_, _06033_);
  and (_33958_, _33957_, _06027_);
  and (_33959_, _33958_, _33954_);
  or (_33961_, _33934_, _14879_);
  and (_33962_, _33961_, _06026_);
  and (_33963_, _33962_, _33936_);
  or (_33964_, _33963_, _09818_);
  or (_33965_, _33964_, _33959_);
  and (_33966_, _09180_, _07688_);
  or (_33967_, _33918_, _07012_);
  or (_33968_, _33967_, _33966_);
  or (_33969_, _33942_, _09827_);
  and (_33970_, _33969_, _05669_);
  and (_33972_, _33970_, _33968_);
  and (_33973_, _33972_, _33965_);
  and (_33974_, _14983_, _07688_);
  or (_33975_, _33974_, _33918_);
  and (_33976_, _33975_, _09833_);
  or (_33977_, _33976_, _06019_);
  or (_33978_, _33977_, _33973_);
  and (_33979_, _33978_, _33921_);
  or (_33980_, _33979_, _06112_);
  and (_33981_, _14876_, _07688_);
  or (_33983_, _33918_, _08751_);
  or (_33984_, _33983_, _33981_);
  and (_33985_, _33984_, _08756_);
  and (_33986_, _33985_, _33980_);
  and (_33987_, _10986_, _07688_);
  or (_33988_, _33987_, _33918_);
  and (_33989_, _33988_, _06284_);
  or (_33990_, _33989_, _33986_);
  and (_33991_, _33990_, _07032_);
  or (_33992_, _33918_, _08273_);
  and (_33994_, _33920_, _06108_);
  and (_33995_, _33994_, _33992_);
  or (_33996_, _33995_, _33991_);
  and (_33997_, _33996_, _06278_);
  and (_33998_, _33926_, _06277_);
  and (_33999_, _33998_, _33992_);
  or (_34000_, _33999_, _06130_);
  or (_34001_, _34000_, _33997_);
  and (_34002_, _14873_, _07688_);
  or (_34003_, _33918_, _08777_);
  or (_34005_, _34003_, _34002_);
  and (_34006_, _34005_, _08782_);
  and (_34007_, _34006_, _34001_);
  nor (_34008_, _10985_, _13311_);
  or (_34009_, _34008_, _33918_);
  and (_34010_, _34009_, _06292_);
  or (_34011_, _34010_, _06316_);
  or (_34012_, _34011_, _34007_);
  or (_34013_, _33923_, _06718_);
  and (_34014_, _34013_, _05653_);
  and (_34016_, _34014_, _34012_);
  and (_34017_, _33951_, _05652_);
  or (_34018_, _34017_, _06047_);
  or (_34019_, _34018_, _34016_);
  and (_34020_, _15055_, _07688_);
  or (_34021_, _33918_, _06048_);
  or (_34022_, _34021_, _34020_);
  and (_34023_, _34022_, _01336_);
  and (_34024_, _34023_, _34019_);
  or (_34025_, _34024_, _33917_);
  and (_43480_, _34025_, _42882_);
  and (_34027_, _01340_, \oc8051_golden_model_1.IE [5]);
  and (_34028_, _13311_, \oc8051_golden_model_1.IE [5]);
  and (_34029_, _08652_, _07688_);
  or (_34030_, _34029_, _34028_);
  or (_34031_, _34030_, _06020_);
  and (_34032_, _15093_, _07688_);
  or (_34033_, _34032_, _34028_);
  or (_34034_, _34033_, _06954_);
  and (_34035_, _07688_, \oc8051_golden_model_1.ACC [5]);
  or (_34037_, _34035_, _34028_);
  and (_34038_, _34037_, _06938_);
  and (_34039_, _06939_, \oc8051_golden_model_1.IE [5]);
  or (_34040_, _34039_, _06102_);
  or (_34041_, _34040_, _34038_);
  and (_34042_, _34041_, _06044_);
  and (_34043_, _34042_, _34034_);
  and (_34044_, _13330_, \oc8051_golden_model_1.IE [5]);
  and (_34045_, _15073_, _08351_);
  or (_34046_, _34045_, _34044_);
  and (_34048_, _34046_, _06043_);
  or (_34049_, _34048_, _06239_);
  or (_34050_, _34049_, _34043_);
  nor (_34051_, _07977_, _13311_);
  or (_34052_, _34051_, _34028_);
  or (_34053_, _34052_, _06848_);
  and (_34054_, _34053_, _34050_);
  or (_34055_, _34054_, _06219_);
  or (_34056_, _34037_, _06220_);
  and (_34057_, _34056_, _06040_);
  and (_34059_, _34057_, _34055_);
  and (_34060_, _15077_, _08351_);
  or (_34061_, _34060_, _34044_);
  and (_34062_, _34061_, _06039_);
  or (_34063_, _34062_, _06032_);
  or (_34064_, _34063_, _34059_);
  or (_34065_, _34044_, _15110_);
  and (_34066_, _34065_, _34046_);
  or (_34067_, _34066_, _06033_);
  and (_34068_, _34067_, _06027_);
  and (_34070_, _34068_, _34064_);
  or (_34071_, _34044_, _15074_);
  and (_34072_, _34071_, _06026_);
  and (_34073_, _34072_, _34046_);
  or (_34074_, _34073_, _09818_);
  or (_34075_, _34074_, _34070_);
  and (_34076_, _09179_, _07688_);
  or (_34077_, _34028_, _07012_);
  or (_34078_, _34077_, _34076_);
  or (_34079_, _34052_, _09827_);
  and (_34081_, _34079_, _05669_);
  and (_34082_, _34081_, _34078_);
  and (_34083_, _34082_, _34075_);
  and (_34084_, _15179_, _07688_);
  or (_34085_, _34084_, _34028_);
  and (_34086_, _34085_, _09833_);
  or (_34087_, _34086_, _06019_);
  or (_34088_, _34087_, _34083_);
  and (_34089_, _34088_, _34031_);
  or (_34090_, _34089_, _06112_);
  and (_34092_, _15195_, _07688_);
  or (_34093_, _34092_, _34028_);
  or (_34094_, _34093_, _08751_);
  and (_34095_, _34094_, _08756_);
  and (_34096_, _34095_, _34090_);
  and (_34097_, _12306_, _07688_);
  or (_34098_, _34097_, _34028_);
  and (_34099_, _34098_, _06284_);
  or (_34100_, _34099_, _34096_);
  and (_34101_, _34100_, _07032_);
  or (_34103_, _34028_, _07980_);
  and (_34104_, _34030_, _06108_);
  and (_34105_, _34104_, _34103_);
  or (_34106_, _34105_, _34101_);
  and (_34107_, _34106_, _06278_);
  and (_34108_, _34037_, _06277_);
  and (_34109_, _34108_, _34103_);
  or (_34110_, _34109_, _06130_);
  or (_34111_, _34110_, _34107_);
  and (_34112_, _15194_, _07688_);
  or (_34113_, _34028_, _08777_);
  or (_34114_, _34113_, _34112_);
  and (_34115_, _34114_, _08782_);
  and (_34116_, _34115_, _34111_);
  nor (_34117_, _10982_, _13311_);
  or (_34118_, _34117_, _34028_);
  and (_34119_, _34118_, _06292_);
  or (_34120_, _34119_, _06316_);
  or (_34121_, _34120_, _34116_);
  or (_34122_, _34033_, _06718_);
  and (_34124_, _34122_, _05653_);
  and (_34125_, _34124_, _34121_);
  and (_34126_, _34061_, _05652_);
  or (_34127_, _34126_, _06047_);
  or (_34128_, _34127_, _34125_);
  and (_34129_, _15253_, _07688_);
  or (_34130_, _34028_, _06048_);
  or (_34131_, _34130_, _34129_);
  and (_34132_, _34131_, _01336_);
  and (_34133_, _34132_, _34128_);
  or (_34135_, _34133_, _34027_);
  and (_43482_, _34135_, _42882_);
  and (_34136_, _01340_, \oc8051_golden_model_1.IE [6]);
  and (_34137_, _13311_, \oc8051_golden_model_1.IE [6]);
  and (_34138_, _15389_, _07688_);
  or (_34139_, _34138_, _34137_);
  or (_34140_, _34139_, _06020_);
  and (_34141_, _15293_, _07688_);
  or (_34142_, _34141_, _34137_);
  or (_34143_, _34142_, _06954_);
  and (_34145_, _07688_, \oc8051_golden_model_1.ACC [6]);
  or (_34146_, _34145_, _34137_);
  and (_34147_, _34146_, _06938_);
  and (_34148_, _06939_, \oc8051_golden_model_1.IE [6]);
  or (_34149_, _34148_, _06102_);
  or (_34150_, _34149_, _34147_);
  and (_34151_, _34150_, _06044_);
  and (_34152_, _34151_, _34143_);
  and (_34153_, _13330_, \oc8051_golden_model_1.IE [6]);
  and (_34154_, _15280_, _08351_);
  or (_34156_, _34154_, _34153_);
  and (_34157_, _34156_, _06043_);
  or (_34158_, _34157_, _06239_);
  or (_34159_, _34158_, _34152_);
  nor (_34160_, _07883_, _13311_);
  or (_34161_, _34160_, _34137_);
  or (_34162_, _34161_, _06848_);
  and (_34163_, _34162_, _34159_);
  or (_34164_, _34163_, _06219_);
  or (_34165_, _34146_, _06220_);
  and (_34167_, _34165_, _06040_);
  and (_34168_, _34167_, _34164_);
  and (_34169_, _15278_, _08351_);
  or (_34170_, _34169_, _34153_);
  and (_34171_, _34170_, _06039_);
  or (_34172_, _34171_, _06032_);
  or (_34173_, _34172_, _34168_);
  or (_34174_, _34153_, _15310_);
  and (_34175_, _34174_, _34156_);
  or (_34176_, _34175_, _06033_);
  and (_34178_, _34176_, _06027_);
  and (_34179_, _34178_, _34173_);
  or (_34180_, _34153_, _15326_);
  and (_34181_, _34180_, _06026_);
  and (_34182_, _34181_, _34156_);
  or (_34183_, _34182_, _09818_);
  or (_34184_, _34183_, _34179_);
  and (_34185_, _09178_, _07688_);
  or (_34186_, _34137_, _07012_);
  or (_34187_, _34186_, _34185_);
  or (_34189_, _34161_, _09827_);
  and (_34190_, _34189_, _05669_);
  and (_34191_, _34190_, _34187_);
  and (_34192_, _34191_, _34184_);
  and (_34193_, _15382_, _07688_);
  or (_34194_, _34193_, _34137_);
  and (_34195_, _34194_, _09833_);
  or (_34196_, _34195_, _06019_);
  or (_34197_, _34196_, _34192_);
  and (_34198_, _34197_, _34140_);
  or (_34200_, _34198_, _06112_);
  and (_34201_, _15399_, _07688_);
  or (_34202_, _34201_, _34137_);
  or (_34203_, _34202_, _08751_);
  and (_34204_, _34203_, _08756_);
  and (_34205_, _34204_, _34200_);
  and (_34206_, _10980_, _07688_);
  or (_34207_, _34206_, _34137_);
  and (_34208_, _34207_, _06284_);
  or (_34209_, _34208_, _34205_);
  and (_34211_, _34209_, _07032_);
  or (_34212_, _34137_, _07886_);
  and (_34213_, _34139_, _06108_);
  and (_34214_, _34213_, _34212_);
  or (_34215_, _34214_, _34211_);
  and (_34216_, _34215_, _06278_);
  and (_34217_, _34146_, _06277_);
  and (_34218_, _34217_, _34212_);
  or (_34219_, _34218_, _06130_);
  or (_34220_, _34219_, _34216_);
  and (_34222_, _15396_, _07688_);
  or (_34223_, _34137_, _08777_);
  or (_34224_, _34223_, _34222_);
  and (_34225_, _34224_, _08782_);
  and (_34226_, _34225_, _34220_);
  nor (_34227_, _10979_, _13311_);
  or (_34228_, _34227_, _34137_);
  and (_34229_, _34228_, _06292_);
  or (_34230_, _34229_, _06316_);
  or (_34231_, _34230_, _34226_);
  or (_34233_, _34142_, _06718_);
  and (_34234_, _34233_, _05653_);
  and (_34235_, _34234_, _34231_);
  and (_34236_, _34170_, _05652_);
  or (_34237_, _34236_, _06047_);
  or (_34238_, _34237_, _34235_);
  and (_34239_, _15451_, _07688_);
  or (_34240_, _34137_, _06048_);
  or (_34241_, _34240_, _34239_);
  and (_34242_, _34241_, _01336_);
  and (_34244_, _34242_, _34238_);
  or (_34245_, _34244_, _34136_);
  and (_43483_, _34245_, _42882_);
  and (_34246_, _01340_, \oc8051_golden_model_1.SCON [0]);
  and (_34247_, _07679_, \oc8051_golden_model_1.ACC [0]);
  and (_34248_, _34247_, _08127_);
  and (_34249_, _13413_, \oc8051_golden_model_1.SCON [0]);
  or (_34250_, _34249_, _06278_);
  or (_34251_, _34250_, _34248_);
  and (_34252_, _07679_, _08672_);
  or (_34254_, _34252_, _34249_);
  or (_34255_, _34254_, _06020_);
  and (_34256_, _09120_, _07679_);
  or (_34257_, _34249_, _07012_);
  or (_34258_, _34257_, _34256_);
  nor (_34259_, _08127_, _13413_);
  or (_34260_, _34259_, _34249_);
  or (_34261_, _34260_, _06954_);
  or (_34262_, _34247_, _34249_);
  and (_34263_, _34262_, _06938_);
  and (_34265_, _06939_, \oc8051_golden_model_1.SCON [0]);
  or (_34266_, _34265_, _06102_);
  or (_34267_, _34266_, _34263_);
  and (_34268_, _34267_, _06044_);
  and (_34269_, _34268_, _34261_);
  and (_34270_, _13432_, \oc8051_golden_model_1.SCON [0]);
  and (_34271_, _14102_, _08347_);
  or (_34272_, _34271_, _34270_);
  and (_34274_, _34272_, _06043_);
  or (_34276_, _34274_, _34269_);
  and (_34279_, _34276_, _06848_);
  and (_34281_, _07679_, _06931_);
  or (_34283_, _34281_, _34249_);
  and (_34285_, _34283_, _06239_);
  or (_34287_, _34285_, _06219_);
  or (_34289_, _34287_, _34279_);
  or (_34291_, _34262_, _06220_);
  and (_34293_, _34291_, _06040_);
  and (_34294_, _34293_, _34289_);
  and (_34295_, _34249_, _06039_);
  or (_34297_, _34295_, _06032_);
  or (_34298_, _34297_, _34294_);
  or (_34299_, _34260_, _06033_);
  and (_34300_, _34299_, _06027_);
  and (_34301_, _34300_, _34298_);
  or (_34302_, _34270_, _14131_);
  and (_34303_, _34302_, _06026_);
  and (_34304_, _34303_, _34272_);
  or (_34305_, _34304_, _09818_);
  or (_34306_, _34305_, _34301_);
  or (_34308_, _34283_, _09827_);
  and (_34309_, _34308_, _05669_);
  and (_34310_, _34309_, _34306_);
  and (_34311_, _34310_, _34258_);
  and (_34312_, _14186_, _07679_);
  or (_34313_, _34312_, _34249_);
  and (_34314_, _34313_, _09833_);
  or (_34315_, _34314_, _06019_);
  or (_34316_, _34315_, _34311_);
  and (_34317_, _34316_, _34255_);
  or (_34319_, _34317_, _06112_);
  and (_34320_, _14086_, _07679_);
  or (_34321_, _34249_, _08751_);
  or (_34322_, _34321_, _34320_);
  and (_34323_, _34322_, _08756_);
  and (_34324_, _34323_, _34319_);
  nor (_34325_, _12302_, _13413_);
  or (_34326_, _34325_, _34249_);
  nor (_34327_, _34248_, _08756_);
  and (_34328_, _34327_, _34326_);
  or (_34330_, _34328_, _34324_);
  and (_34331_, _34330_, _07032_);
  nand (_34332_, _34254_, _06108_);
  nor (_34333_, _34332_, _34259_);
  or (_34334_, _34333_, _06277_);
  or (_34335_, _34334_, _34331_);
  and (_34336_, _34335_, _34251_);
  or (_34337_, _34336_, _06130_);
  and (_34338_, _14083_, _07679_);
  or (_34339_, _34249_, _08777_);
  or (_34341_, _34339_, _34338_);
  and (_34342_, _34341_, _08782_);
  and (_34343_, _34342_, _34337_);
  and (_34344_, _34326_, _06292_);
  or (_34345_, _34344_, _06316_);
  or (_34346_, _34345_, _34343_);
  or (_34347_, _34260_, _06718_);
  and (_34348_, _34347_, _34346_);
  or (_34349_, _34348_, _05652_);
  or (_34350_, _34249_, _05653_);
  and (_34352_, _34350_, _34349_);
  or (_34353_, _34352_, _06047_);
  or (_34354_, _34260_, _06048_);
  and (_34355_, _34354_, _01336_);
  and (_34356_, _34355_, _34353_);
  or (_34357_, _34356_, _34246_);
  and (_43484_, _34357_, _42882_);
  not (_34358_, \oc8051_golden_model_1.SCON [1]);
  nor (_34359_, _01336_, _34358_);
  nor (_34360_, _07679_, _34358_);
  nor (_34362_, _10993_, _13413_);
  or (_34363_, _34362_, _34360_);
  or (_34364_, _34363_, _08782_);
  nor (_34365_, _13413_, _07132_);
  or (_34366_, _34365_, _34360_);
  or (_34367_, _34366_, _06848_);
  or (_34368_, _07679_, \oc8051_golden_model_1.SCON [1]);
  and (_34369_, _14284_, _07679_);
  not (_34370_, _34369_);
  and (_34371_, _34370_, _34368_);
  or (_34373_, _34371_, _06954_);
  and (_34374_, _07679_, \oc8051_golden_model_1.ACC [1]);
  or (_34375_, _34374_, _34360_);
  and (_34376_, _34375_, _06938_);
  nor (_34377_, _06938_, _34358_);
  or (_34378_, _34377_, _06102_);
  or (_34379_, _34378_, _34376_);
  and (_34380_, _34379_, _06044_);
  and (_34381_, _34380_, _34373_);
  nor (_34382_, _08347_, _34358_);
  and (_34384_, _14266_, _08347_);
  or (_34385_, _34384_, _34382_);
  and (_34386_, _34385_, _06043_);
  or (_34387_, _34386_, _06239_);
  or (_34388_, _34387_, _34381_);
  and (_34389_, _34388_, _34367_);
  or (_34390_, _34389_, _06219_);
  or (_34391_, _34375_, _06220_);
  and (_34392_, _34391_, _06040_);
  and (_34393_, _34392_, _34390_);
  and (_34395_, _14273_, _08347_);
  or (_34396_, _34395_, _34382_);
  and (_34397_, _34396_, _06039_);
  or (_34398_, _34397_, _06032_);
  or (_34399_, _34398_, _34393_);
  and (_34400_, _34384_, _14302_);
  or (_34401_, _34382_, _06033_);
  or (_34402_, _34401_, _34400_);
  and (_34403_, _34402_, _06027_);
  and (_34404_, _34403_, _34399_);
  or (_34406_, _34382_, _14267_);
  and (_34407_, _34406_, _06026_);
  and (_34408_, _34407_, _34385_);
  or (_34409_, _34408_, _09818_);
  or (_34410_, _34409_, _34404_);
  and (_34411_, _09075_, _07679_);
  or (_34412_, _34360_, _07012_);
  or (_34413_, _34412_, _34411_);
  or (_34414_, _34366_, _09827_);
  and (_34415_, _34414_, _05669_);
  and (_34417_, _34415_, _34413_);
  and (_34418_, _34417_, _34410_);
  and (_34419_, _14367_, _07679_);
  or (_34420_, _34419_, _34360_);
  and (_34421_, _34420_, _09833_);
  or (_34422_, _34421_, _34418_);
  and (_34423_, _34422_, _06020_);
  nand (_34424_, _07679_, _06832_);
  and (_34425_, _34368_, _06019_);
  and (_34426_, _34425_, _34424_);
  or (_34428_, _34426_, _34423_);
  and (_34429_, _34428_, _08751_);
  or (_34430_, _14263_, _13413_);
  and (_34431_, _34368_, _06112_);
  and (_34432_, _34431_, _34430_);
  or (_34433_, _34432_, _06284_);
  or (_34434_, _34433_, _34429_);
  nand (_34435_, _10992_, _07679_);
  and (_34436_, _34435_, _34363_);
  or (_34437_, _34436_, _08756_);
  and (_34439_, _34437_, _07032_);
  and (_34440_, _34439_, _34434_);
  or (_34441_, _14261_, _13413_);
  and (_34442_, _34368_, _06108_);
  and (_34443_, _34442_, _34441_);
  or (_34444_, _34443_, _06277_);
  or (_34445_, _34444_, _34440_);
  nor (_34446_, _34360_, _06278_);
  nand (_34447_, _34446_, _34435_);
  and (_34448_, _34447_, _08777_);
  and (_34450_, _34448_, _34445_);
  or (_34451_, _34424_, _08078_);
  and (_34452_, _34368_, _06130_);
  and (_34453_, _34452_, _34451_);
  or (_34454_, _34453_, _06292_);
  or (_34455_, _34454_, _34450_);
  and (_34456_, _34455_, _34364_);
  or (_34457_, _34456_, _06316_);
  or (_34458_, _34371_, _06718_);
  and (_34459_, _34458_, _05653_);
  and (_34461_, _34459_, _34457_);
  and (_34462_, _34396_, _05652_);
  or (_34463_, _34462_, _06047_);
  or (_34464_, _34463_, _34461_);
  or (_34465_, _34360_, _06048_);
  or (_34466_, _34465_, _34369_);
  and (_34467_, _34466_, _01336_);
  and (_34468_, _34467_, _34464_);
  or (_34469_, _34468_, _34359_);
  and (_43486_, _34469_, _42882_);
  and (_34471_, _01340_, \oc8051_golden_model_1.SCON [2]);
  and (_34472_, _13413_, \oc8051_golden_model_1.SCON [2]);
  and (_34473_, _07679_, _08730_);
  or (_34474_, _34473_, _34472_);
  or (_34475_, _34474_, _06020_);
  nor (_34476_, _13413_, _07530_);
  or (_34477_, _34476_, _34472_);
  and (_34478_, _34477_, _06239_);
  and (_34479_, _13432_, \oc8051_golden_model_1.SCON [2]);
  and (_34480_, _14497_, _08347_);
  or (_34482_, _34480_, _34479_);
  or (_34483_, _34482_, _06044_);
  and (_34484_, _14493_, _07679_);
  or (_34485_, _34484_, _34472_);
  and (_34486_, _34485_, _06102_);
  and (_34487_, _06939_, \oc8051_golden_model_1.SCON [2]);
  and (_34488_, _07679_, \oc8051_golden_model_1.ACC [2]);
  or (_34489_, _34488_, _34472_);
  and (_34490_, _34489_, _06938_);
  or (_34491_, _34490_, _34487_);
  and (_34493_, _34491_, _06954_);
  or (_34494_, _34493_, _06043_);
  or (_34495_, _34494_, _34486_);
  and (_34496_, _34495_, _34483_);
  and (_34497_, _34496_, _06848_);
  or (_34498_, _34497_, _34478_);
  or (_34499_, _34498_, _06219_);
  or (_34500_, _34489_, _06220_);
  and (_34501_, _34500_, _06040_);
  and (_34502_, _34501_, _34499_);
  and (_34504_, _14479_, _08347_);
  or (_34505_, _34504_, _34479_);
  and (_34506_, _34505_, _06039_);
  or (_34507_, _34506_, _06032_);
  or (_34508_, _34507_, _34502_);
  or (_34509_, _34479_, _14512_);
  and (_34510_, _34509_, _34482_);
  or (_34511_, _34510_, _06033_);
  and (_34512_, _34511_, _06027_);
  and (_34513_, _34512_, _34508_);
  or (_34515_, _34479_, _14525_);
  and (_34516_, _34515_, _06026_);
  and (_34517_, _34516_, _34482_);
  or (_34518_, _34517_, _09818_);
  or (_34519_, _34518_, _34513_);
  and (_34520_, _09182_, _07679_);
  or (_34521_, _34472_, _07012_);
  or (_34522_, _34521_, _34520_);
  or (_34523_, _34477_, _09827_);
  and (_34524_, _34523_, _05669_);
  and (_34526_, _34524_, _34522_);
  and (_34527_, _34526_, _34519_);
  and (_34528_, _14580_, _07679_);
  or (_34529_, _34528_, _34472_);
  and (_34530_, _34529_, _09833_);
  or (_34531_, _34530_, _06019_);
  or (_34532_, _34531_, _34527_);
  and (_34533_, _34532_, _34475_);
  or (_34534_, _34533_, _06112_);
  and (_34535_, _14596_, _07679_);
  or (_34537_, _34535_, _34472_);
  or (_34538_, _34537_, _08751_);
  and (_34539_, _34538_, _08756_);
  and (_34540_, _34539_, _34534_);
  and (_34541_, _10991_, _07679_);
  or (_34542_, _34541_, _34472_);
  and (_34543_, _34542_, _06284_);
  or (_34544_, _34543_, _34540_);
  and (_34545_, _34544_, _07032_);
  or (_34546_, _34472_, _08177_);
  and (_34548_, _34474_, _06108_);
  and (_34549_, _34548_, _34546_);
  or (_34550_, _34549_, _34545_);
  and (_34551_, _34550_, _06278_);
  and (_34552_, _34489_, _06277_);
  and (_34553_, _34552_, _34546_);
  or (_34554_, _34553_, _06130_);
  or (_34555_, _34554_, _34551_);
  and (_34556_, _14593_, _07679_);
  or (_34557_, _34472_, _08777_);
  or (_34559_, _34557_, _34556_);
  and (_34560_, _34559_, _08782_);
  and (_34561_, _34560_, _34555_);
  nor (_34562_, _10990_, _13413_);
  or (_34563_, _34562_, _34472_);
  and (_34564_, _34563_, _06292_);
  or (_34565_, _34564_, _06316_);
  or (_34566_, _34565_, _34561_);
  or (_34567_, _34485_, _06718_);
  and (_34568_, _34567_, _05653_);
  and (_34570_, _34568_, _34566_);
  and (_34571_, _34505_, _05652_);
  or (_34572_, _34571_, _06047_);
  or (_34573_, _34572_, _34570_);
  and (_34574_, _14657_, _07679_);
  or (_34575_, _34472_, _06048_);
  or (_34576_, _34575_, _34574_);
  and (_34577_, _34576_, _01336_);
  and (_34578_, _34577_, _34573_);
  or (_34579_, _34578_, _34471_);
  and (_43487_, _34579_, _42882_);
  and (_34581_, _01340_, \oc8051_golden_model_1.SCON [3]);
  and (_34582_, _13413_, \oc8051_golden_model_1.SCON [3]);
  and (_34583_, _07679_, _08662_);
  or (_34584_, _34583_, _34582_);
  or (_34585_, _34584_, _06020_);
  and (_34586_, _14672_, _07679_);
  or (_34587_, _34586_, _34582_);
  or (_34588_, _34587_, _06954_);
  and (_34589_, _07679_, \oc8051_golden_model_1.ACC [3]);
  or (_34591_, _34589_, _34582_);
  and (_34592_, _34591_, _06938_);
  and (_34593_, _06939_, \oc8051_golden_model_1.SCON [3]);
  or (_34594_, _34593_, _06102_);
  or (_34595_, _34594_, _34592_);
  and (_34596_, _34595_, _06044_);
  and (_34597_, _34596_, _34588_);
  and (_34598_, _13432_, \oc8051_golden_model_1.SCON [3]);
  and (_34599_, _14683_, _08347_);
  or (_34600_, _34599_, _34598_);
  and (_34602_, _34600_, _06043_);
  or (_34603_, _34602_, _06239_);
  or (_34604_, _34603_, _34597_);
  nor (_34605_, _13413_, _07353_);
  or (_34606_, _34605_, _34582_);
  or (_34607_, _34606_, _06848_);
  and (_34608_, _34607_, _34604_);
  or (_34609_, _34608_, _06219_);
  or (_34610_, _34591_, _06220_);
  and (_34611_, _34610_, _06040_);
  and (_34613_, _34611_, _34609_);
  and (_34614_, _14681_, _08347_);
  or (_34615_, _34614_, _34598_);
  and (_34616_, _34615_, _06039_);
  or (_34617_, _34616_, _06032_);
  or (_34618_, _34617_, _34613_);
  or (_34619_, _34598_, _14708_);
  and (_34620_, _34619_, _34600_);
  or (_34621_, _34620_, _06033_);
  and (_34622_, _34621_, _06027_);
  and (_34624_, _34622_, _34618_);
  and (_34625_, _14724_, _08347_);
  or (_34626_, _34625_, _34598_);
  and (_34627_, _34626_, _06026_);
  or (_34628_, _34627_, _09818_);
  or (_34629_, _34628_, _34624_);
  and (_34630_, _09181_, _07679_);
  or (_34631_, _34582_, _07012_);
  or (_34632_, _34631_, _34630_);
  or (_34633_, _34606_, _09827_);
  and (_34635_, _34633_, _05669_);
  and (_34636_, _34635_, _34632_);
  and (_34637_, _34636_, _34629_);
  and (_34638_, _14778_, _07679_);
  or (_34639_, _34638_, _34582_);
  and (_34640_, _34639_, _09833_);
  or (_34641_, _34640_, _06019_);
  or (_34642_, _34641_, _34637_);
  and (_34643_, _34642_, _34585_);
  or (_34644_, _34643_, _06112_);
  and (_34646_, _14793_, _07679_);
  or (_34647_, _34582_, _08751_);
  or (_34648_, _34647_, _34646_);
  and (_34649_, _34648_, _08756_);
  and (_34650_, _34649_, _34644_);
  and (_34651_, _12299_, _07679_);
  or (_34652_, _34651_, _34582_);
  and (_34653_, _34652_, _06284_);
  or (_34654_, _34653_, _34650_);
  and (_34655_, _34654_, _07032_);
  or (_34657_, _34582_, _08029_);
  and (_34658_, _34584_, _06108_);
  and (_34659_, _34658_, _34657_);
  or (_34660_, _34659_, _34655_);
  and (_34661_, _34660_, _06278_);
  and (_34662_, _34591_, _06277_);
  and (_34663_, _34662_, _34657_);
  or (_34664_, _34663_, _06130_);
  or (_34665_, _34664_, _34661_);
  and (_34666_, _14792_, _07679_);
  or (_34668_, _34582_, _08777_);
  or (_34669_, _34668_, _34666_);
  and (_34670_, _34669_, _08782_);
  and (_34671_, _34670_, _34665_);
  nor (_34672_, _10988_, _13413_);
  or (_34673_, _34672_, _34582_);
  and (_34674_, _34673_, _06292_);
  or (_34675_, _34674_, _06316_);
  or (_34676_, _34675_, _34671_);
  or (_34677_, _34587_, _06718_);
  and (_34679_, _34677_, _05653_);
  and (_34680_, _34679_, _34676_);
  and (_34681_, _34615_, _05652_);
  or (_34682_, _34681_, _06047_);
  or (_34683_, _34682_, _34680_);
  and (_34684_, _14849_, _07679_);
  or (_34685_, _34582_, _06048_);
  or (_34686_, _34685_, _34684_);
  and (_34687_, _34686_, _01336_);
  and (_34688_, _34687_, _34683_);
  or (_34690_, _34688_, _34581_);
  and (_43488_, _34690_, _42882_);
  and (_34691_, _01340_, \oc8051_golden_model_1.SCON [4]);
  and (_34692_, _13413_, \oc8051_golden_model_1.SCON [4]);
  and (_34693_, _08665_, _07679_);
  or (_34694_, _34693_, _34692_);
  or (_34695_, _34694_, _06020_);
  and (_34696_, _14887_, _07679_);
  or (_34697_, _34696_, _34692_);
  or (_34698_, _34697_, _06954_);
  and (_34700_, _07679_, \oc8051_golden_model_1.ACC [4]);
  or (_34701_, _34700_, _34692_);
  and (_34702_, _34701_, _06938_);
  and (_34703_, _06939_, \oc8051_golden_model_1.SCON [4]);
  or (_34704_, _34703_, _06102_);
  or (_34705_, _34704_, _34702_);
  and (_34706_, _34705_, _06044_);
  and (_34707_, _34706_, _34698_);
  and (_34708_, _13432_, \oc8051_golden_model_1.SCON [4]);
  and (_34709_, _14878_, _08347_);
  or (_34711_, _34709_, _34708_);
  and (_34712_, _34711_, _06043_);
  or (_34713_, _34712_, _06239_);
  or (_34714_, _34713_, _34707_);
  nor (_34715_, _08270_, _13413_);
  or (_34716_, _34715_, _34692_);
  or (_34717_, _34716_, _06848_);
  and (_34718_, _34717_, _34714_);
  or (_34719_, _34718_, _06219_);
  or (_34720_, _34701_, _06220_);
  and (_34722_, _34720_, _06040_);
  and (_34723_, _34722_, _34719_);
  and (_34724_, _14882_, _08347_);
  or (_34725_, _34724_, _34708_);
  and (_34726_, _34725_, _06039_);
  or (_34727_, _34726_, _06032_);
  or (_34728_, _34727_, _34723_);
  or (_34729_, _34708_, _14914_);
  and (_34730_, _34729_, _34711_);
  or (_34731_, _34730_, _06033_);
  and (_34733_, _34731_, _06027_);
  and (_34734_, _34733_, _34728_);
  or (_34735_, _34708_, _14879_);
  and (_34736_, _34735_, _06026_);
  and (_34737_, _34736_, _34711_);
  or (_34738_, _34737_, _09818_);
  or (_34739_, _34738_, _34734_);
  and (_34740_, _09180_, _07679_);
  or (_34741_, _34692_, _07012_);
  or (_34742_, _34741_, _34740_);
  or (_34744_, _34716_, _09827_);
  and (_34745_, _34744_, _05669_);
  and (_34746_, _34745_, _34742_);
  and (_34747_, _34746_, _34739_);
  and (_34748_, _14983_, _07679_);
  or (_34749_, _34748_, _34692_);
  and (_34750_, _34749_, _09833_);
  or (_34751_, _34750_, _06019_);
  or (_34752_, _34751_, _34747_);
  and (_34753_, _34752_, _34695_);
  or (_34755_, _34753_, _06112_);
  and (_34756_, _14876_, _07679_);
  or (_34757_, _34756_, _34692_);
  or (_34758_, _34757_, _08751_);
  and (_34759_, _34758_, _08756_);
  and (_34760_, _34759_, _34755_);
  and (_34761_, _10986_, _07679_);
  or (_34762_, _34761_, _34692_);
  and (_34763_, _34762_, _06284_);
  or (_34764_, _34763_, _34760_);
  and (_34766_, _34764_, _07032_);
  or (_34767_, _34692_, _08273_);
  and (_34768_, _34694_, _06108_);
  and (_34769_, _34768_, _34767_);
  or (_34770_, _34769_, _34766_);
  and (_34771_, _34770_, _06278_);
  and (_34772_, _34701_, _06277_);
  and (_34773_, _34772_, _34767_);
  or (_34774_, _34773_, _06130_);
  or (_34775_, _34774_, _34771_);
  and (_34777_, _14873_, _07679_);
  or (_34778_, _34692_, _08777_);
  or (_34779_, _34778_, _34777_);
  and (_34780_, _34779_, _08782_);
  and (_34781_, _34780_, _34775_);
  nor (_34782_, _10985_, _13413_);
  or (_34783_, _34782_, _34692_);
  and (_34784_, _34783_, _06292_);
  or (_34785_, _34784_, _06316_);
  or (_34786_, _34785_, _34781_);
  or (_34788_, _34697_, _06718_);
  and (_34789_, _34788_, _05653_);
  and (_34790_, _34789_, _34786_);
  and (_34791_, _34725_, _05652_);
  or (_34792_, _34791_, _06047_);
  or (_34793_, _34792_, _34790_);
  and (_34794_, _15055_, _07679_);
  or (_34795_, _34692_, _06048_);
  or (_34796_, _34795_, _34794_);
  and (_34797_, _34796_, _01336_);
  and (_34799_, _34797_, _34793_);
  or (_34800_, _34799_, _34691_);
  and (_43489_, _34800_, _42882_);
  and (_34801_, _01340_, \oc8051_golden_model_1.SCON [5]);
  and (_34802_, _13413_, \oc8051_golden_model_1.SCON [5]);
  and (_34803_, _08652_, _07679_);
  or (_34804_, _34803_, _34802_);
  or (_34805_, _34804_, _06020_);
  and (_34806_, _15093_, _07679_);
  or (_34807_, _34806_, _34802_);
  or (_34809_, _34807_, _06954_);
  and (_34810_, _07679_, \oc8051_golden_model_1.ACC [5]);
  or (_34811_, _34810_, _34802_);
  and (_34812_, _34811_, _06938_);
  and (_34813_, _06939_, \oc8051_golden_model_1.SCON [5]);
  or (_34814_, _34813_, _06102_);
  or (_34815_, _34814_, _34812_);
  and (_34816_, _34815_, _06044_);
  and (_34817_, _34816_, _34809_);
  and (_34818_, _13432_, \oc8051_golden_model_1.SCON [5]);
  and (_34820_, _15073_, _08347_);
  or (_34821_, _34820_, _34818_);
  and (_34822_, _34821_, _06043_);
  or (_34823_, _34822_, _06239_);
  or (_34824_, _34823_, _34817_);
  nor (_34825_, _07977_, _13413_);
  or (_34826_, _34825_, _34802_);
  or (_34827_, _34826_, _06848_);
  and (_34828_, _34827_, _34824_);
  or (_34829_, _34828_, _06219_);
  or (_34831_, _34811_, _06220_);
  and (_34832_, _34831_, _06040_);
  and (_34833_, _34832_, _34829_);
  and (_34834_, _15077_, _08347_);
  or (_34835_, _34834_, _34818_);
  and (_34836_, _34835_, _06039_);
  or (_34837_, _34836_, _06032_);
  or (_34838_, _34837_, _34833_);
  or (_34839_, _34818_, _15110_);
  and (_34840_, _34839_, _34821_);
  or (_34842_, _34840_, _06033_);
  and (_34843_, _34842_, _06027_);
  and (_34844_, _34843_, _34838_);
  or (_34845_, _34818_, _15074_);
  and (_34846_, _34845_, _06026_);
  and (_34847_, _34846_, _34821_);
  or (_34848_, _34847_, _09818_);
  or (_34849_, _34848_, _34844_);
  and (_34850_, _09179_, _07679_);
  or (_34851_, _34802_, _07012_);
  or (_34853_, _34851_, _34850_);
  or (_34854_, _34826_, _09827_);
  and (_34855_, _34854_, _05669_);
  and (_34856_, _34855_, _34853_);
  and (_34857_, _34856_, _34849_);
  and (_34858_, _15179_, _07679_);
  or (_34859_, _34858_, _34802_);
  and (_34860_, _34859_, _09833_);
  or (_34861_, _34860_, _06019_);
  or (_34862_, _34861_, _34857_);
  and (_34864_, _34862_, _34805_);
  or (_34865_, _34864_, _06112_);
  and (_34866_, _15195_, _07679_);
  or (_34867_, _34802_, _08751_);
  or (_34868_, _34867_, _34866_);
  and (_34869_, _34868_, _08756_);
  and (_34870_, _34869_, _34865_);
  and (_34871_, _12306_, _07679_);
  or (_34872_, _34871_, _34802_);
  and (_34873_, _34872_, _06284_);
  or (_34875_, _34873_, _34870_);
  and (_34876_, _34875_, _07032_);
  or (_34877_, _34802_, _07980_);
  and (_34878_, _34804_, _06108_);
  and (_34879_, _34878_, _34877_);
  or (_34880_, _34879_, _34876_);
  and (_34881_, _34880_, _06278_);
  and (_34882_, _34811_, _06277_);
  and (_34883_, _34882_, _34877_);
  or (_34884_, _34883_, _06130_);
  or (_34886_, _34884_, _34881_);
  and (_34887_, _15194_, _07679_);
  or (_34888_, _34802_, _08777_);
  or (_34889_, _34888_, _34887_);
  and (_34890_, _34889_, _08782_);
  and (_34891_, _34890_, _34886_);
  nor (_34892_, _10982_, _13413_);
  or (_34893_, _34892_, _34802_);
  and (_34894_, _34893_, _06292_);
  or (_34895_, _34894_, _06316_);
  or (_34897_, _34895_, _34891_);
  or (_34898_, _34807_, _06718_);
  and (_34899_, _34898_, _05653_);
  and (_34900_, _34899_, _34897_);
  and (_34901_, _34835_, _05652_);
  or (_34902_, _34901_, _06047_);
  or (_34903_, _34902_, _34900_);
  and (_34904_, _15253_, _07679_);
  or (_34905_, _34802_, _06048_);
  or (_34906_, _34905_, _34904_);
  and (_34907_, _34906_, _01336_);
  and (_34908_, _34907_, _34903_);
  or (_34909_, _34908_, _34801_);
  and (_43490_, _34909_, _42882_);
  and (_34910_, _01340_, \oc8051_golden_model_1.SCON [6]);
  and (_34911_, _13413_, \oc8051_golden_model_1.SCON [6]);
  and (_34912_, _15389_, _07679_);
  or (_34913_, _34912_, _34911_);
  or (_34914_, _34913_, _06020_);
  and (_34915_, _15293_, _07679_);
  or (_34917_, _34915_, _34911_);
  or (_34918_, _34917_, _06954_);
  and (_34919_, _07679_, \oc8051_golden_model_1.ACC [6]);
  or (_34920_, _34919_, _34911_);
  and (_34921_, _34920_, _06938_);
  and (_34922_, _06939_, \oc8051_golden_model_1.SCON [6]);
  or (_34923_, _34922_, _06102_);
  or (_34924_, _34923_, _34921_);
  and (_34925_, _34924_, _06044_);
  and (_34926_, _34925_, _34918_);
  and (_34928_, _13432_, \oc8051_golden_model_1.SCON [6]);
  and (_34929_, _15280_, _08347_);
  or (_34930_, _34929_, _34928_);
  and (_34931_, _34930_, _06043_);
  or (_34932_, _34931_, _06239_);
  or (_34933_, _34932_, _34926_);
  nor (_34934_, _07883_, _13413_);
  or (_34935_, _34934_, _34911_);
  or (_34936_, _34935_, _06848_);
  and (_34937_, _34936_, _34933_);
  or (_34939_, _34937_, _06219_);
  or (_34940_, _34920_, _06220_);
  and (_34941_, _34940_, _06040_);
  and (_34942_, _34941_, _34939_);
  and (_34943_, _15278_, _08347_);
  or (_34944_, _34943_, _34928_);
  and (_34945_, _34944_, _06039_);
  or (_34946_, _34945_, _06032_);
  or (_34947_, _34946_, _34942_);
  or (_34948_, _34928_, _15310_);
  and (_34950_, _34948_, _34930_);
  or (_34951_, _34950_, _06033_);
  and (_34952_, _34951_, _06027_);
  and (_34953_, _34952_, _34947_);
  or (_34954_, _34928_, _15326_);
  and (_34955_, _34954_, _06026_);
  and (_34956_, _34955_, _34930_);
  or (_34957_, _34956_, _09818_);
  or (_34958_, _34957_, _34953_);
  and (_34959_, _09178_, _07679_);
  or (_34961_, _34911_, _07012_);
  or (_34962_, _34961_, _34959_);
  or (_34963_, _34935_, _09827_);
  and (_34964_, _34963_, _05669_);
  and (_34965_, _34964_, _34962_);
  and (_34966_, _34965_, _34958_);
  and (_34967_, _15382_, _07679_);
  or (_34968_, _34967_, _34911_);
  and (_34969_, _34968_, _09833_);
  or (_34970_, _34969_, _06019_);
  or (_34972_, _34970_, _34966_);
  and (_34973_, _34972_, _34914_);
  or (_34974_, _34973_, _06112_);
  and (_34975_, _15399_, _07679_);
  or (_34976_, _34975_, _34911_);
  or (_34977_, _34976_, _08751_);
  and (_34978_, _34977_, _08756_);
  and (_34979_, _34978_, _34974_);
  and (_34980_, _10980_, _07679_);
  or (_34981_, _34980_, _34911_);
  and (_34983_, _34981_, _06284_);
  or (_34984_, _34983_, _34979_);
  and (_34985_, _34984_, _07032_);
  or (_34986_, _34911_, _07886_);
  and (_34987_, _34913_, _06108_);
  and (_34988_, _34987_, _34986_);
  or (_34989_, _34988_, _34985_);
  and (_34990_, _34989_, _06278_);
  and (_34991_, _34920_, _06277_);
  and (_34992_, _34991_, _34986_);
  or (_34994_, _34992_, _06130_);
  or (_34995_, _34994_, _34990_);
  and (_34996_, _15396_, _07679_);
  or (_34997_, _34911_, _08777_);
  or (_34998_, _34997_, _34996_);
  and (_34999_, _34998_, _08782_);
  and (_35000_, _34999_, _34995_);
  nor (_35001_, _10979_, _13413_);
  or (_35002_, _35001_, _34911_);
  and (_35003_, _35002_, _06292_);
  or (_35005_, _35003_, _06316_);
  or (_35006_, _35005_, _35000_);
  or (_35007_, _34917_, _06718_);
  and (_35008_, _35007_, _05653_);
  and (_35009_, _35008_, _35006_);
  and (_35010_, _34944_, _05652_);
  or (_35011_, _35010_, _06047_);
  or (_35012_, _35011_, _35009_);
  and (_35013_, _15451_, _07679_);
  or (_35014_, _34911_, _06048_);
  or (_35016_, _35014_, _35013_);
  and (_35017_, _35016_, _01336_);
  and (_35018_, _35017_, _35012_);
  or (_35019_, _35018_, _34910_);
  and (_43491_, _35019_, _42882_);
  nor (_35020_, _01336_, _06029_);
  nor (_35021_, _07727_, _06029_);
  and (_35022_, _07833_, \oc8051_golden_model_1.ACC [0]);
  and (_35023_, _35022_, _08127_);
  or (_35024_, _35023_, _35021_);
  or (_35026_, _35024_, _06278_);
  or (_35027_, _35021_, _07012_);
  and (_35028_, _09120_, _07833_);
  or (_35029_, _35028_, _35027_);
  and (_35030_, _07727_, _06931_);
  or (_35031_, _35021_, _09827_);
  or (_35032_, _35031_, _35030_);
  nor (_35033_, _08127_, _13575_);
  or (_35034_, _35033_, _35021_);
  or (_35035_, _35034_, _06954_);
  nor (_35037_, _35022_, _35021_);
  nor (_35038_, _35037_, _06939_);
  nor (_35039_, _06938_, _06029_);
  or (_35040_, _35039_, _06102_);
  or (_35041_, _35040_, _35038_);
  and (_35042_, _35041_, _06848_);
  nand (_35043_, _35042_, _35035_);
  and (_35044_, _35043_, _06544_);
  and (_35045_, _35037_, _06219_);
  or (_35046_, _35045_, _06038_);
  or (_35048_, _35046_, _35044_);
  and (_35049_, _07012_, _06982_);
  and (_35050_, _35049_, _09827_);
  nand (_35051_, _35050_, _35048_);
  and (_35052_, _35051_, _35032_);
  and (_35053_, _35052_, _35029_);
  or (_35054_, _35053_, _09833_);
  and (_35055_, _14186_, _07727_);
  or (_35056_, _35021_, _05669_);
  or (_35057_, _35056_, _35055_);
  and (_35059_, _35057_, _06020_);
  and (_35060_, _35059_, _35054_);
  and (_35061_, _07833_, _08672_);
  or (_35062_, _35061_, _35021_);
  and (_35063_, _35062_, _06019_);
  or (_35064_, _35063_, _06112_);
  or (_35065_, _35064_, _35060_);
  and (_35066_, _14086_, _07833_);
  or (_35067_, _35066_, _35021_);
  or (_35068_, _35067_, _08751_);
  and (_35070_, _35068_, _08756_);
  and (_35071_, _35070_, _35065_);
  nor (_35072_, _12302_, _13575_);
  or (_35073_, _35072_, _35021_);
  nor (_35074_, _35023_, _08756_);
  and (_35075_, _35074_, _35073_);
  or (_35076_, _35075_, _35071_);
  and (_35077_, _35076_, _07032_);
  nand (_35078_, _35062_, _06108_);
  nor (_35079_, _35078_, _35033_);
  or (_35081_, _35079_, _06277_);
  or (_35082_, _35081_, _35077_);
  and (_35083_, _35082_, _35026_);
  or (_35084_, _35083_, _06130_);
  and (_35085_, _14083_, _07727_);
  or (_35086_, _35021_, _08777_);
  or (_35087_, _35086_, _35085_);
  and (_35088_, _35087_, _08782_);
  and (_35089_, _35088_, _35084_);
  and (_35090_, _35073_, _06292_);
  or (_35092_, _35090_, _19256_);
  or (_35093_, _35092_, _35089_);
  or (_35094_, _35034_, _06408_);
  and (_35095_, _35094_, _01336_);
  and (_35096_, _35095_, _35093_);
  or (_35097_, _35096_, _35020_);
  and (_43493_, _35097_, _42882_);
  nand (_35098_, _06298_, \oc8051_golden_model_1.SP [1]);
  nand (_35099_, _07727_, _06832_);
  or (_35100_, _35099_, _08078_);
  or (_35102_, _07727_, \oc8051_golden_model_1.SP [1]);
  and (_35103_, _35102_, _06130_);
  and (_35104_, _35103_, _35100_);
  and (_35105_, _35102_, _09833_);
  or (_35106_, _14367_, _13575_);
  and (_35107_, _35106_, _35105_);
  and (_35108_, _14284_, _07727_);
  not (_35109_, _35108_);
  and (_35110_, _35109_, _35102_);
  or (_35111_, _35110_, _06954_);
  nand (_35113_, _06943_, \oc8051_golden_model_1.SP [1]);
  nor (_35114_, _07727_, _06847_);
  and (_35115_, _07833_, \oc8051_golden_model_1.ACC [1]);
  or (_35116_, _35115_, _35114_);
  and (_35117_, _35116_, _06938_);
  nor (_35118_, _06938_, _06847_);
  or (_35119_, _35118_, _06943_);
  or (_35120_, _35119_, _35117_);
  and (_35121_, _35120_, _35113_);
  or (_35122_, _35121_, _06102_);
  and (_35124_, _35122_, _05690_);
  and (_35125_, _35124_, _35111_);
  nor (_35126_, _05690_, \oc8051_golden_model_1.SP [1]);
  or (_35127_, _35126_, _06239_);
  or (_35128_, _35127_, _35125_);
  nand (_35129_, _07083_, _06239_);
  and (_35130_, _35129_, _35128_);
  or (_35131_, _35130_, _06219_);
  or (_35132_, _35116_, _06220_);
  and (_35133_, _35132_, _07364_);
  and (_35135_, _35133_, _35131_);
  or (_35136_, _13568_, _07169_);
  or (_35137_, _35136_, _35135_);
  or (_35138_, _07271_, _06847_);
  and (_35139_, _35138_, _09827_);
  and (_35140_, _35139_, _35137_);
  nand (_35141_, _07727_, _07132_);
  and (_35142_, _35102_, _09815_);
  and (_35143_, _35142_, _35141_);
  or (_35144_, _35143_, _07011_);
  or (_35146_, _35144_, _35140_);
  or (_35147_, _35114_, _07012_);
  and (_35148_, _09075_, _07833_);
  or (_35149_, _35148_, _35147_);
  and (_35150_, _35149_, _05669_);
  and (_35151_, _35150_, _35146_);
  or (_35152_, _35151_, _35107_);
  and (_35153_, _35152_, _06020_);
  and (_35154_, _35102_, _06019_);
  and (_35155_, _35154_, _35099_);
  or (_35157_, _35155_, _05724_);
  or (_35158_, _35157_, _35153_);
  and (_35159_, _05724_, \oc8051_golden_model_1.SP [1]);
  nor (_35160_, _35159_, _06112_);
  and (_35161_, _35160_, _35158_);
  or (_35162_, _14263_, _13575_);
  and (_35163_, _35102_, _06112_);
  and (_35164_, _35163_, _35162_);
  or (_35165_, _35164_, _06284_);
  or (_35166_, _35165_, _35161_);
  and (_35168_, _10994_, _07833_);
  or (_35169_, _35168_, _35114_);
  or (_35170_, _35169_, _08756_);
  and (_35171_, _35170_, _07032_);
  and (_35172_, _35171_, _35166_);
  or (_35173_, _14261_, _13575_);
  and (_35174_, _35102_, _06108_);
  and (_35175_, _35174_, _35173_);
  or (_35176_, _35175_, _06277_);
  or (_35177_, _35176_, _35172_);
  and (_35179_, _35115_, _08078_);
  or (_35180_, _35179_, _35114_);
  or (_35181_, _35180_, _06278_);
  and (_35182_, _35181_, _35177_);
  or (_35183_, _35182_, _05736_);
  and (_35184_, _05736_, \oc8051_golden_model_1.SP [1]);
  nor (_35185_, _35184_, _06130_);
  and (_35186_, _35185_, _35183_);
  or (_35187_, _35186_, _35104_);
  and (_35188_, _35187_, _08782_);
  nor (_35190_, _10993_, _13575_);
  or (_35191_, _35190_, _35114_);
  and (_35192_, _35191_, _06292_);
  or (_35193_, _35192_, _06298_);
  or (_35194_, _35193_, _35188_);
  nand (_35195_, _35194_, _35098_);
  nor (_35196_, _06049_, _05732_);
  nand (_35197_, _35196_, _35195_);
  or (_35198_, _35196_, _06847_);
  and (_35199_, _35198_, _06718_);
  and (_35201_, _35199_, _35197_);
  and (_35202_, _35110_, _06316_);
  or (_35203_, _35202_, _07458_);
  or (_35204_, _35203_, _35201_);
  or (_35205_, _07059_, _06847_);
  and (_35206_, _35205_, _06048_);
  and (_35207_, _35206_, _35204_);
  or (_35208_, _35108_, _35114_);
  and (_35209_, _35208_, _06047_);
  or (_35210_, _35209_, _01340_);
  or (_35212_, _35210_, _35207_);
  or (_35213_, _01336_, \oc8051_golden_model_1.SP [1]);
  and (_35214_, _35213_, _42882_);
  and (_43494_, _35214_, _35212_);
  nor (_35215_, _01336_, _06447_);
  nand (_35216_, _14449_, _05724_);
  nor (_35217_, _13575_, _07530_);
  nor (_35218_, _07727_, _06447_);
  or (_35219_, _35218_, _09827_);
  or (_35220_, _35219_, _35217_);
  and (_35222_, _14493_, _07727_);
  or (_35223_, _35222_, _35218_);
  or (_35224_, _35223_, _06954_);
  and (_35225_, _07833_, \oc8051_golden_model_1.ACC [2]);
  or (_35226_, _35225_, _35218_);
  or (_35227_, _35226_, _06939_);
  or (_35228_, _06938_, \oc8051_golden_model_1.SP [2]);
  and (_35229_, _35228_, _07233_);
  and (_35230_, _35229_, _35227_);
  and (_35231_, _07622_, _06943_);
  or (_35233_, _35231_, _06102_);
  or (_35234_, _35233_, _35230_);
  and (_35235_, _35234_, _05690_);
  and (_35236_, _35235_, _35224_);
  nor (_35237_, _14449_, _05690_);
  or (_35238_, _35237_, _06239_);
  or (_35239_, _35238_, _35236_);
  nand (_35240_, _08415_, _06239_);
  and (_35241_, _35240_, _35239_);
  or (_35242_, _35241_, _06219_);
  or (_35244_, _35226_, _06220_);
  and (_35245_, _35244_, _07364_);
  and (_35246_, _35245_, _35242_);
  or (_35247_, _07561_, _07355_);
  or (_35248_, _35247_, _35246_);
  or (_35249_, _07622_, _05686_);
  and (_35250_, _35249_, _05673_);
  and (_35251_, _35250_, _35248_);
  nor (_35252_, _14449_, _05673_);
  or (_35253_, _35252_, _09815_);
  or (_35255_, _35253_, _35251_);
  and (_35256_, _35255_, _35220_);
  or (_35257_, _35256_, _07011_);
  or (_35258_, _35218_, _07012_);
  and (_35259_, _09182_, _07833_);
  or (_35260_, _35259_, _35258_);
  and (_35261_, _35260_, _05669_);
  and (_35262_, _35261_, _35257_);
  and (_35263_, _14580_, _07833_);
  or (_35264_, _35263_, _35218_);
  and (_35266_, _35264_, _09833_);
  or (_35267_, _35266_, _06019_);
  or (_35268_, _35267_, _35262_);
  and (_35269_, _07833_, _08730_);
  or (_35270_, _35269_, _35218_);
  or (_35271_, _35270_, _06020_);
  and (_35272_, _35271_, _35268_);
  or (_35273_, _35272_, _05724_);
  and (_35274_, _35273_, _35216_);
  or (_35275_, _35274_, _06112_);
  and (_35277_, _14596_, _07833_);
  or (_35278_, _35277_, _35218_);
  or (_35279_, _35278_, _08751_);
  and (_35280_, _35279_, _08756_);
  and (_35281_, _35280_, _35275_);
  and (_35282_, _10991_, _07833_);
  or (_35283_, _35282_, _35218_);
  and (_35284_, _35283_, _06284_);
  or (_35285_, _35284_, _35281_);
  and (_35286_, _35285_, _07032_);
  or (_35288_, _35218_, _08177_);
  and (_35289_, _35270_, _06108_);
  and (_35290_, _35289_, _35288_);
  or (_35291_, _35290_, _35286_);
  and (_35292_, _35291_, _12494_);
  and (_35293_, _35226_, _06277_);
  and (_35294_, _35293_, _35288_);
  and (_35295_, _07622_, _05736_);
  or (_35296_, _35295_, _06130_);
  or (_35297_, _35296_, _35294_);
  or (_35299_, _35297_, _35292_);
  and (_35300_, _14593_, _07727_);
  or (_35301_, _35218_, _08777_);
  or (_35302_, _35301_, _35300_);
  and (_35303_, _35302_, _35299_);
  or (_35304_, _35303_, _06292_);
  nor (_35305_, _10990_, _13575_);
  or (_35306_, _35305_, _35218_);
  or (_35307_, _35306_, _08782_);
  and (_35308_, _35307_, _13619_);
  and (_35310_, _35308_, _35304_);
  and (_35311_, _14449_, _06298_);
  or (_35312_, _35311_, _05732_);
  or (_35313_, _35312_, _35310_);
  nand (_35314_, _14449_, _05732_);
  and (_35315_, _35314_, _06050_);
  and (_35316_, _35315_, _35313_);
  and (_35317_, _14449_, _06049_);
  or (_35318_, _35317_, _06316_);
  or (_35319_, _35318_, _35316_);
  or (_35321_, _35223_, _06718_);
  and (_35322_, _35321_, _07059_);
  and (_35323_, _35322_, _35319_);
  nor (_35324_, _14449_, _07059_);
  or (_35325_, _35324_, _06047_);
  or (_35326_, _35325_, _35323_);
  and (_35327_, _14657_, _07727_);
  or (_35328_, _35218_, _06048_);
  or (_35329_, _35328_, _35327_);
  and (_35330_, _35329_, _01336_);
  and (_35332_, _35330_, _35326_);
  or (_35333_, _35332_, _35215_);
  and (_43495_, _35333_, _42882_);
  nor (_35334_, _01336_, _06238_);
  or (_35335_, _07625_, _07059_);
  nand (_35336_, _14453_, _05724_);
  nor (_35337_, _13575_, _07353_);
  nor (_35338_, _07727_, _06238_);
  or (_35339_, _35338_, _07011_);
  or (_35340_, _35339_, _35337_);
  and (_35342_, _35340_, _09818_);
  and (_35343_, _14672_, _07727_);
  or (_35344_, _35343_, _35338_);
  or (_35345_, _35344_, _06954_);
  and (_35346_, _07833_, \oc8051_golden_model_1.ACC [3]);
  or (_35347_, _35346_, _35338_);
  or (_35348_, _35347_, _06939_);
  or (_35349_, _06938_, \oc8051_golden_model_1.SP [3]);
  and (_35350_, _35349_, _07233_);
  and (_35351_, _35350_, _35348_);
  and (_35353_, _07625_, _06943_);
  or (_35354_, _35353_, _06102_);
  or (_35355_, _35354_, _35351_);
  and (_35356_, _35355_, _05690_);
  and (_35357_, _35356_, _35345_);
  nor (_35358_, _14453_, _05690_);
  or (_35359_, _35358_, _06239_);
  or (_35360_, _35359_, _35357_);
  nand (_35361_, _08405_, _06239_);
  and (_35362_, _35361_, _35360_);
  or (_35364_, _35362_, _06219_);
  or (_35365_, _35347_, _06220_);
  and (_35366_, _35365_, _07364_);
  and (_35367_, _35366_, _35364_);
  or (_35368_, _07404_, _13568_);
  or (_35369_, _35368_, _35367_);
  or (_35370_, _07625_, _07271_);
  and (_35371_, _35370_, _09827_);
  and (_35372_, _35371_, _35369_);
  or (_35373_, _35372_, _35342_);
  or (_35375_, _35338_, _07012_);
  and (_35376_, _09181_, _07833_);
  or (_35377_, _35376_, _35375_);
  and (_35378_, _35377_, _05669_);
  and (_35379_, _35378_, _35373_);
  and (_35380_, _14778_, _07833_);
  or (_35381_, _35380_, _35338_);
  and (_35382_, _35381_, _09833_);
  or (_35383_, _35382_, _06019_);
  or (_35384_, _35383_, _35379_);
  and (_35386_, _07833_, _08662_);
  or (_35387_, _35386_, _35338_);
  or (_35388_, _35387_, _06020_);
  and (_35389_, _35388_, _35384_);
  or (_35390_, _35389_, _05724_);
  and (_35391_, _35390_, _35336_);
  or (_35392_, _35391_, _06112_);
  and (_35393_, _14793_, _07833_);
  or (_35394_, _35393_, _35338_);
  or (_35395_, _35394_, _08751_);
  and (_35397_, _35395_, _08756_);
  and (_35398_, _35397_, _35392_);
  and (_35399_, _12299_, _07833_);
  or (_35400_, _35399_, _35338_);
  and (_35401_, _35400_, _06284_);
  or (_35402_, _35401_, _35398_);
  and (_35403_, _35402_, _07032_);
  or (_35404_, _35338_, _08029_);
  and (_35405_, _35387_, _06108_);
  and (_35406_, _35405_, _35404_);
  or (_35408_, _35406_, _35403_);
  and (_35409_, _35408_, _12494_);
  and (_35410_, _35347_, _06277_);
  and (_35411_, _35410_, _35404_);
  and (_35412_, _07625_, _05736_);
  or (_35413_, _35412_, _06130_);
  or (_35414_, _35413_, _35411_);
  or (_35415_, _35414_, _35409_);
  and (_35416_, _14792_, _07727_);
  or (_35417_, _35338_, _08777_);
  or (_35419_, _35417_, _35416_);
  and (_35420_, _35419_, _35415_);
  or (_35421_, _35420_, _06292_);
  nor (_35422_, _10988_, _13575_);
  or (_35423_, _35422_, _35338_);
  or (_35424_, _35423_, _08782_);
  and (_35425_, _35424_, _13619_);
  and (_35426_, _35425_, _35421_);
  nor (_35427_, _08402_, _06238_);
  or (_35428_, _35427_, _08403_);
  and (_35430_, _35428_, _06298_);
  or (_35431_, _35430_, _05732_);
  or (_35432_, _35431_, _35426_);
  nand (_35433_, _14453_, _05732_);
  and (_35434_, _35433_, _35432_);
  or (_35435_, _35434_, _06049_);
  or (_35436_, _35428_, _06050_);
  and (_35437_, _35436_, _06718_);
  and (_35438_, _35437_, _35435_);
  and (_35439_, _35344_, _06316_);
  or (_35441_, _35439_, _07458_);
  or (_35442_, _35441_, _35438_);
  and (_35443_, _35442_, _35335_);
  or (_35444_, _35443_, _06047_);
  and (_35445_, _14849_, _07727_);
  or (_35446_, _35338_, _06048_);
  or (_35447_, _35446_, _35445_);
  and (_35448_, _35447_, _01336_);
  and (_35449_, _35448_, _35444_);
  or (_35450_, _35449_, _35334_);
  and (_43496_, _35450_, _42882_);
  nor (_35452_, _01336_, _13552_);
  nor (_35453_, _07360_, \oc8051_golden_model_1.SP [4]);
  nor (_35454_, _35453_, _13516_);
  or (_35455_, _35454_, _07059_);
  or (_35456_, _35454_, _05734_);
  or (_35457_, _35454_, _07271_);
  nor (_35458_, _07727_, _13552_);
  and (_35459_, _14887_, _07727_);
  or (_35460_, _35459_, _35458_);
  or (_35462_, _35460_, _06954_);
  and (_35463_, _07833_, \oc8051_golden_model_1.ACC [4]);
  or (_35464_, _35463_, _35458_);
  or (_35465_, _35464_, _06939_);
  or (_35466_, _06938_, \oc8051_golden_model_1.SP [4]);
  and (_35467_, _35466_, _07233_);
  and (_35468_, _35467_, _35465_);
  and (_35469_, _35454_, _06943_);
  or (_35470_, _35469_, _06102_);
  or (_35471_, _35470_, _35468_);
  and (_35473_, _35471_, _05690_);
  and (_35474_, _35473_, _35462_);
  and (_35475_, _35454_, _07272_);
  or (_35476_, _35475_, _06239_);
  or (_35477_, _35476_, _35474_);
  and (_35478_, _13553_, _06029_);
  nor (_35479_, _08404_, _13552_);
  nor (_35480_, _35479_, _35478_);
  nand (_35481_, _35480_, _06239_);
  and (_35482_, _35481_, _35477_);
  or (_35484_, _35482_, _06219_);
  or (_35485_, _35464_, _06220_);
  and (_35486_, _35485_, _07364_);
  and (_35487_, _35486_, _35484_);
  and (_35488_, _07361_, \oc8051_golden_model_1.SP [4]);
  nor (_35489_, _07361_, \oc8051_golden_model_1.SP [4]);
  nor (_35490_, _35489_, _35488_);
  nand (_35491_, _35490_, _06038_);
  nand (_35492_, _35491_, _07271_);
  or (_35493_, _35492_, _35487_);
  and (_35495_, _35493_, _35457_);
  nor (_35496_, _11995_, _05660_);
  and (_35497_, _06227_, _05659_);
  and (_35498_, _06133_, _05659_);
  nor (_35499_, _35498_, _35497_);
  not (_35500_, _35499_);
  or (_35501_, _35500_, _35496_);
  or (_35502_, _35501_, _35495_);
  and (_35503_, _06096_, _05659_);
  not (_35504_, _35501_);
  nor (_35506_, _08270_, _13575_);
  or (_35507_, _35506_, _35458_);
  nor (_35508_, _35507_, _35504_);
  nor (_35509_, _35508_, _35503_);
  and (_35510_, _35509_, _35502_);
  and (_35511_, _35507_, _35503_);
  or (_35512_, _35511_, _07011_);
  or (_35513_, _35512_, _35510_);
  or (_35514_, _35458_, _07012_);
  and (_35515_, _09180_, _07833_);
  or (_35517_, _35515_, _35514_);
  and (_35518_, _35517_, _35513_);
  or (_35519_, _35518_, _09833_);
  and (_35520_, _14983_, _07833_);
  or (_35521_, _35520_, _35458_);
  or (_35522_, _35521_, _05669_);
  and (_35523_, _35522_, _06020_);
  and (_35524_, _35523_, _35519_);
  and (_35525_, _08665_, _07833_);
  or (_35526_, _35525_, _35458_);
  and (_35528_, _35526_, _06019_);
  or (_35529_, _35528_, _05724_);
  or (_35530_, _35529_, _35524_);
  or (_35531_, _35454_, _13587_);
  and (_35532_, _35531_, _35530_);
  or (_35533_, _35532_, _06112_);
  and (_35534_, _14876_, _07727_);
  or (_35535_, _35458_, _08751_);
  or (_35536_, _35535_, _35534_);
  and (_35537_, _35536_, _08756_);
  and (_35539_, _35537_, _35533_);
  and (_35540_, _10986_, _07833_);
  or (_35541_, _35540_, _35458_);
  and (_35542_, _35541_, _06284_);
  or (_35543_, _35542_, _35539_);
  and (_35544_, _35543_, _07032_);
  or (_35545_, _35458_, _08273_);
  and (_35546_, _35526_, _06108_);
  and (_35547_, _35546_, _35545_);
  or (_35548_, _35547_, _35544_);
  and (_35550_, _35548_, _12494_);
  and (_35551_, _35464_, _06277_);
  and (_35552_, _35551_, _35545_);
  and (_35553_, _35454_, _05736_);
  or (_35554_, _35553_, _06130_);
  or (_35555_, _35554_, _35552_);
  or (_35556_, _35555_, _35550_);
  and (_35557_, _14873_, _07727_);
  or (_35558_, _35458_, _08777_);
  or (_35559_, _35558_, _35557_);
  and (_35561_, _35559_, _35556_);
  or (_35562_, _35561_, _06292_);
  nor (_35563_, _10985_, _13575_);
  or (_35564_, _35563_, _35458_);
  or (_35565_, _35564_, _08782_);
  and (_35566_, _35565_, _13619_);
  and (_35567_, _35566_, _35562_);
  nor (_35568_, _08403_, _13552_);
  or (_35569_, _35568_, _13553_);
  and (_35570_, _35569_, _06298_);
  or (_35572_, _35570_, _05732_);
  or (_35573_, _35572_, _35567_);
  and (_35574_, _35573_, _35456_);
  or (_35575_, _35574_, _06049_);
  or (_35576_, _35569_, _06050_);
  and (_35577_, _35576_, _06718_);
  and (_35578_, _35577_, _35575_);
  and (_35579_, _35460_, _06316_);
  or (_35580_, _35579_, _07458_);
  or (_35581_, _35580_, _35578_);
  and (_35583_, _35581_, _35455_);
  or (_35584_, _35583_, _06047_);
  and (_35585_, _15055_, _07727_);
  or (_35586_, _35458_, _06048_);
  or (_35587_, _35586_, _35585_);
  and (_35588_, _35587_, _01336_);
  and (_35589_, _35588_, _35584_);
  or (_35590_, _35589_, _35452_);
  and (_43497_, _35590_, _42882_);
  nor (_35591_, _01336_, _13551_);
  nor (_35593_, _13516_, \oc8051_golden_model_1.SP [5]);
  nor (_35594_, _35593_, _13517_);
  or (_35595_, _35594_, _07059_);
  or (_35596_, _35594_, _05734_);
  nor (_35597_, _07977_, _13575_);
  nor (_35598_, _07727_, _13551_);
  or (_35599_, _35598_, _07011_);
  or (_35600_, _35599_, _35597_);
  and (_35601_, _35600_, _09818_);
  and (_35602_, _15093_, _07727_);
  or (_35604_, _35602_, _35598_);
  or (_35605_, _35604_, _06954_);
  and (_35606_, _07833_, \oc8051_golden_model_1.ACC [5]);
  or (_35607_, _35606_, _35598_);
  or (_35608_, _35607_, _06939_);
  or (_35609_, _06938_, \oc8051_golden_model_1.SP [5]);
  and (_35610_, _35609_, _07233_);
  and (_35611_, _35610_, _35608_);
  and (_35612_, _35594_, _06943_);
  or (_35613_, _35612_, _06102_);
  or (_35615_, _35613_, _35611_);
  and (_35616_, _35615_, _05690_);
  and (_35617_, _35616_, _35605_);
  and (_35618_, _35594_, _07272_);
  or (_35619_, _35618_, _06239_);
  or (_35620_, _35619_, _35617_);
  and (_35621_, _13554_, _06029_);
  nor (_35622_, _35478_, _13551_);
  nor (_35623_, _35622_, _35621_);
  nand (_35624_, _35623_, _06239_);
  and (_35626_, _35624_, _35620_);
  or (_35627_, _35626_, _06219_);
  or (_35628_, _35607_, _06220_);
  and (_35629_, _35628_, _07364_);
  and (_35630_, _35629_, _35627_);
  nor (_35631_, _35488_, \oc8051_golden_model_1.SP [5]);
  nor (_35632_, _35631_, _13527_);
  nand (_35633_, _35632_, _06038_);
  nand (_35634_, _35633_, _07271_);
  or (_35635_, _35634_, _35630_);
  or (_35636_, _35594_, _07271_);
  and (_35637_, _35636_, _09827_);
  and (_35638_, _35637_, _35635_);
  or (_35639_, _35638_, _35601_);
  or (_35640_, _35598_, _07012_);
  and (_35641_, _09179_, _07833_);
  or (_35642_, _35641_, _35640_);
  and (_35643_, _35642_, _05669_);
  and (_35644_, _35643_, _35639_);
  and (_35645_, _15179_, _07833_);
  or (_35647_, _35645_, _35598_);
  and (_35648_, _35647_, _09833_);
  or (_35649_, _35648_, _06019_);
  or (_35650_, _35649_, _35644_);
  and (_35651_, _08652_, _07833_);
  or (_35652_, _35651_, _35598_);
  or (_35653_, _35652_, _06020_);
  and (_35654_, _35653_, _35650_);
  or (_35655_, _35654_, _05724_);
  or (_35656_, _35594_, _13587_);
  and (_35658_, _35656_, _35655_);
  or (_35659_, _35658_, _06112_);
  and (_35660_, _15195_, _07727_);
  or (_35661_, _35598_, _08751_);
  or (_35662_, _35661_, _35660_);
  and (_35663_, _35662_, _08756_);
  and (_35664_, _35663_, _35659_);
  and (_35665_, _12306_, _07833_);
  or (_35666_, _35665_, _35598_);
  and (_35667_, _35666_, _06284_);
  or (_35669_, _35667_, _35664_);
  and (_35670_, _35669_, _07032_);
  or (_35671_, _35598_, _07980_);
  and (_35672_, _35652_, _06108_);
  and (_35673_, _35672_, _35671_);
  or (_35674_, _35673_, _35670_);
  and (_35675_, _35674_, _12494_);
  and (_35676_, _35607_, _06277_);
  and (_35677_, _35676_, _35671_);
  and (_35678_, _35594_, _05736_);
  or (_35680_, _35678_, _06130_);
  or (_35681_, _35680_, _35677_);
  or (_35682_, _35681_, _35675_);
  and (_35683_, _15194_, _07727_);
  or (_35684_, _35598_, _08777_);
  or (_35685_, _35684_, _35683_);
  and (_35686_, _35685_, _35682_);
  or (_35687_, _35686_, _06292_);
  nor (_35688_, _10982_, _13575_);
  or (_35689_, _35688_, _35598_);
  or (_35691_, _35689_, _08782_);
  and (_35692_, _35691_, _13619_);
  and (_35693_, _35692_, _35687_);
  nor (_35694_, _13553_, _13551_);
  or (_35695_, _35694_, _13554_);
  and (_35696_, _35695_, _06298_);
  or (_35697_, _35696_, _05732_);
  or (_35698_, _35697_, _35693_);
  and (_35699_, _35698_, _35596_);
  or (_35700_, _35699_, _06049_);
  or (_35702_, _35695_, _06050_);
  and (_35703_, _35702_, _06718_);
  and (_35704_, _35703_, _35700_);
  and (_35705_, _35604_, _06316_);
  or (_35706_, _35705_, _07458_);
  or (_35707_, _35706_, _35704_);
  and (_35708_, _35707_, _35595_);
  or (_35709_, _35708_, _06047_);
  and (_35710_, _15253_, _07727_);
  or (_35711_, _35598_, _06048_);
  or (_35713_, _35711_, _35710_);
  and (_35714_, _35713_, _01336_);
  and (_35715_, _35714_, _35709_);
  or (_35716_, _35715_, _35591_);
  and (_43498_, _35716_, _42882_);
  nor (_35717_, _01336_, _13550_);
  nor (_35718_, _07883_, _13575_);
  nor (_35719_, _07727_, _13550_);
  or (_35720_, _35719_, _09827_);
  or (_35721_, _35720_, _35718_);
  and (_35723_, _15293_, _07727_);
  or (_35724_, _35723_, _35719_);
  or (_35725_, _35724_, _06954_);
  and (_35726_, _07833_, \oc8051_golden_model_1.ACC [6]);
  or (_35727_, _35726_, _35719_);
  or (_35728_, _35727_, _06939_);
  or (_35729_, _06938_, \oc8051_golden_model_1.SP [6]);
  and (_35730_, _35729_, _07233_);
  and (_35731_, _35730_, _35728_);
  nor (_35732_, _13517_, \oc8051_golden_model_1.SP [6]);
  nor (_35734_, _35732_, _13518_);
  and (_35735_, _35734_, _06943_);
  or (_35736_, _35735_, _06102_);
  or (_35737_, _35736_, _35731_);
  and (_35738_, _35737_, _05690_);
  and (_35739_, _35738_, _35725_);
  and (_35740_, _35734_, _07272_);
  or (_35741_, _35740_, _06239_);
  or (_35742_, _35741_, _35739_);
  nor (_35743_, _35621_, _13550_);
  nor (_35745_, _35743_, _13556_);
  nand (_35746_, _35745_, _06239_);
  and (_35747_, _35746_, _35742_);
  or (_35748_, _35747_, _06219_);
  or (_35749_, _35727_, _06220_);
  and (_35750_, _35749_, _07364_);
  and (_35751_, _35750_, _35748_);
  nor (_35752_, _13527_, \oc8051_golden_model_1.SP [6]);
  nor (_35753_, _35752_, _13528_);
  and (_35754_, _35753_, _06038_);
  or (_35756_, _35754_, _35751_);
  and (_35757_, _35756_, _07271_);
  and (_35758_, _35734_, _13568_);
  or (_35759_, _35758_, _09815_);
  or (_35760_, _35759_, _35757_);
  and (_35761_, _35760_, _35721_);
  or (_35762_, _35761_, _07011_);
  or (_35763_, _35719_, _07012_);
  and (_35764_, _09178_, _07833_);
  or (_35765_, _35764_, _35763_);
  and (_35767_, _35765_, _05669_);
  and (_35768_, _35767_, _35762_);
  and (_35769_, _15382_, _07833_);
  or (_35770_, _35769_, _35719_);
  and (_35771_, _35770_, _09833_);
  or (_35772_, _35771_, _06019_);
  or (_35773_, _35772_, _35768_);
  and (_35774_, _15389_, _07833_);
  or (_35775_, _35774_, _35719_);
  or (_35776_, _35775_, _06020_);
  and (_35778_, _35776_, _35773_);
  or (_35779_, _35778_, _05724_);
  or (_35780_, _35734_, _13587_);
  and (_35781_, _35780_, _35779_);
  or (_35782_, _35781_, _06112_);
  and (_35783_, _15399_, _07727_);
  or (_35784_, _35719_, _08751_);
  or (_35785_, _35784_, _35783_);
  and (_35786_, _35785_, _08756_);
  and (_35787_, _35786_, _35782_);
  and (_35789_, _10980_, _07833_);
  or (_35790_, _35789_, _35719_);
  and (_35791_, _35790_, _06284_);
  or (_35792_, _35791_, _35787_);
  and (_35793_, _35792_, _07032_);
  or (_35794_, _35719_, _07886_);
  and (_35795_, _35775_, _06108_);
  and (_35796_, _35795_, _35794_);
  or (_35797_, _35796_, _35793_);
  and (_35798_, _35797_, _12494_);
  and (_35800_, _35727_, _06277_);
  and (_35801_, _35800_, _35794_);
  and (_35802_, _35734_, _05736_);
  or (_35803_, _35802_, _06130_);
  or (_35804_, _35803_, _35801_);
  or (_35805_, _35804_, _35798_);
  and (_35806_, _15396_, _07727_);
  or (_35807_, _35719_, _08777_);
  or (_35808_, _35807_, _35806_);
  and (_35809_, _35808_, _35805_);
  or (_35811_, _35809_, _06292_);
  nor (_35812_, _10979_, _13575_);
  or (_35813_, _35812_, _35719_);
  or (_35814_, _35813_, _08782_);
  and (_35815_, _35814_, _13619_);
  and (_35816_, _35815_, _35811_);
  nor (_35817_, _13554_, _13550_);
  or (_35818_, _35817_, _13555_);
  and (_35819_, _35818_, _06298_);
  or (_35820_, _35819_, _05732_);
  or (_35822_, _35820_, _35816_);
  or (_35823_, _35734_, _05734_);
  and (_35824_, _35823_, _35822_);
  or (_35825_, _35824_, _06049_);
  or (_35826_, _35818_, _06050_);
  and (_35827_, _35826_, _35825_);
  or (_35828_, _35827_, _06316_);
  or (_35829_, _35724_, _06718_);
  and (_35830_, _35829_, _07059_);
  and (_35831_, _35830_, _35828_);
  and (_35833_, _35734_, _07458_);
  or (_35834_, _35833_, _06047_);
  or (_35835_, _35834_, _35831_);
  and (_35836_, _15451_, _07727_);
  or (_35837_, _35719_, _06048_);
  or (_35838_, _35837_, _35836_);
  and (_35839_, _35838_, _01336_);
  and (_35840_, _35839_, _35835_);
  or (_35841_, _35840_, _35717_);
  and (_43499_, _35841_, _42882_);
  not (_35843_, \oc8051_golden_model_1.SBUF [0]);
  nor (_35844_, _01336_, _35843_);
  nand (_35845_, _10995_, _07681_);
  nor (_35846_, _07681_, _35843_);
  nor (_35847_, _35846_, _06278_);
  nand (_35848_, _35847_, _35845_);
  and (_35849_, _09120_, _07681_);
  or (_35850_, _35846_, _07012_);
  or (_35851_, _35850_, _35849_);
  and (_35852_, _07681_, _06931_);
  nor (_35854_, _35852_, _35846_);
  nand (_35855_, _35854_, _09815_);
  nor (_35856_, _08127_, _13650_);
  or (_35857_, _35856_, _35846_);
  or (_35858_, _35857_, _06954_);
  and (_35859_, _07681_, \oc8051_golden_model_1.ACC [0]);
  nor (_35860_, _35859_, _35846_);
  nor (_35861_, _35860_, _06939_);
  nor (_35862_, _06938_, _35843_);
  or (_35863_, _35862_, _06102_);
  or (_35865_, _35863_, _35861_);
  and (_35866_, _35865_, _06848_);
  and (_35867_, _35866_, _35858_);
  nor (_35868_, _35854_, _06848_);
  or (_35869_, _35868_, _35867_);
  nand (_35870_, _35869_, _06220_);
  or (_35871_, _35860_, _06220_);
  and (_35872_, _35871_, _09817_);
  nand (_35873_, _35872_, _35870_);
  and (_35874_, _35873_, _35855_);
  and (_35876_, _35874_, _35851_);
  or (_35877_, _35876_, _09833_);
  and (_35878_, _14186_, _07681_);
  or (_35879_, _35878_, _35846_);
  or (_35880_, _35879_, _05669_);
  and (_35881_, _35880_, _06020_);
  and (_35882_, _35881_, _35877_);
  and (_35883_, _07681_, _08672_);
  or (_35884_, _35883_, _35846_);
  and (_35885_, _35884_, _06019_);
  or (_35887_, _35885_, _06112_);
  or (_35888_, _35887_, _35882_);
  and (_35889_, _14086_, _07681_);
  or (_35890_, _35846_, _08751_);
  or (_35891_, _35890_, _35889_);
  and (_35892_, _35891_, _08756_);
  and (_35893_, _35892_, _35888_);
  nor (_35894_, _12302_, _13650_);
  or (_35895_, _35894_, _35846_);
  and (_35896_, _35845_, _06284_);
  and (_35898_, _35896_, _35895_);
  or (_35899_, _35898_, _35893_);
  and (_35900_, _35899_, _07032_);
  nand (_35901_, _35884_, _06108_);
  nor (_35902_, _35901_, _35856_);
  or (_35903_, _35902_, _06277_);
  or (_35904_, _35903_, _35900_);
  and (_35905_, _35904_, _35848_);
  or (_35906_, _35905_, _06130_);
  and (_35907_, _14083_, _07681_);
  or (_35909_, _35846_, _08777_);
  or (_35910_, _35909_, _35907_);
  and (_35911_, _35910_, _08782_);
  and (_35912_, _35911_, _35906_);
  and (_35913_, _35895_, _06292_);
  or (_35914_, _35913_, _19256_);
  or (_35915_, _35914_, _35912_);
  or (_35916_, _35857_, _06408_);
  and (_35917_, _35916_, _01336_);
  and (_35918_, _35917_, _35915_);
  or (_35920_, _35918_, _35844_);
  and (_43501_, _35920_, _42882_);
  not (_35921_, \oc8051_golden_model_1.SBUF [1]);
  nor (_35922_, _01336_, _35921_);
  or (_35923_, _14367_, _13650_);
  or (_35924_, _07681_, \oc8051_golden_model_1.SBUF [1]);
  and (_35925_, _35924_, _09833_);
  and (_35926_, _35925_, _35923_);
  and (_35927_, _09075_, _07681_);
  nor (_35928_, _07681_, _35921_);
  or (_35930_, _35928_, _07012_);
  or (_35931_, _35930_, _35927_);
  and (_35932_, _14284_, _07681_);
  not (_35933_, _35932_);
  and (_35934_, _35933_, _35924_);
  or (_35935_, _35934_, _06954_);
  and (_35936_, _07681_, \oc8051_golden_model_1.ACC [1]);
  or (_35937_, _35936_, _35928_);
  and (_35938_, _35937_, _06938_);
  nor (_35939_, _06938_, _35921_);
  or (_35941_, _35939_, _06102_);
  or (_35942_, _35941_, _35938_);
  and (_35943_, _35942_, _06848_);
  and (_35944_, _35943_, _35935_);
  nor (_35945_, _13650_, _07132_);
  or (_35946_, _35945_, _35928_);
  and (_35947_, _35946_, _06239_);
  or (_35948_, _35947_, _35944_);
  and (_35949_, _35948_, _06220_);
  and (_35950_, _35937_, _06219_);
  or (_35952_, _35950_, _09818_);
  or (_35953_, _35952_, _35949_);
  or (_35954_, _35946_, _09827_);
  and (_35955_, _35954_, _05669_);
  and (_35956_, _35955_, _35953_);
  and (_35957_, _35956_, _35931_);
  or (_35958_, _35957_, _35926_);
  and (_35959_, _35958_, _06020_);
  nand (_35960_, _07681_, _06832_);
  and (_35961_, _35924_, _06019_);
  and (_35963_, _35961_, _35960_);
  or (_35964_, _35963_, _35959_);
  and (_35965_, _35964_, _08751_);
  or (_35966_, _14263_, _13650_);
  and (_35967_, _35924_, _06112_);
  and (_35968_, _35967_, _35966_);
  or (_35969_, _35968_, _06284_);
  or (_35970_, _35969_, _35965_);
  nor (_35971_, _10993_, _13650_);
  or (_35972_, _35971_, _35928_);
  nand (_35974_, _10992_, _07681_);
  and (_35975_, _35974_, _35972_);
  or (_35976_, _35975_, _08756_);
  and (_35977_, _35976_, _07032_);
  and (_35978_, _35977_, _35970_);
  or (_35979_, _14261_, _13650_);
  and (_35980_, _35924_, _06108_);
  and (_35981_, _35980_, _35979_);
  or (_35982_, _35981_, _06277_);
  or (_35983_, _35982_, _35978_);
  nor (_35985_, _35928_, _06278_);
  nand (_35986_, _35985_, _35974_);
  and (_35987_, _35986_, _08777_);
  and (_35988_, _35987_, _35983_);
  or (_35989_, _35960_, _08078_);
  and (_35990_, _35924_, _06130_);
  and (_35991_, _35990_, _35989_);
  or (_35992_, _35991_, _06292_);
  or (_35993_, _35992_, _35988_);
  or (_35994_, _35972_, _08782_);
  and (_35996_, _35994_, _06718_);
  and (_35997_, _35996_, _35993_);
  and (_35998_, _35934_, _06316_);
  or (_35999_, _35998_, _06047_);
  or (_36000_, _35999_, _35997_);
  or (_36001_, _35928_, _06048_);
  or (_36002_, _36001_, _35932_);
  and (_36003_, _36002_, _01336_);
  and (_36004_, _36003_, _36000_);
  or (_36005_, _36004_, _35922_);
  and (_43502_, _36005_, _42882_);
  not (_36007_, \oc8051_golden_model_1.SBUF [2]);
  nor (_36008_, _01336_, _36007_);
  nor (_36009_, _07681_, _36007_);
  or (_36010_, _36009_, _08177_);
  and (_36011_, _07681_, _08730_);
  or (_36012_, _36011_, _36009_);
  and (_36013_, _36012_, _06108_);
  and (_36014_, _36013_, _36010_);
  and (_36015_, _09182_, _07681_);
  or (_36017_, _36009_, _07012_);
  or (_36018_, _36017_, _36015_);
  nor (_36019_, _13650_, _07530_);
  nor (_36020_, _36019_, _36009_);
  nand (_36021_, _36020_, _09815_);
  and (_36022_, _14493_, _07681_);
  or (_36023_, _36022_, _36009_);
  or (_36024_, _36023_, _06954_);
  and (_36025_, _07681_, \oc8051_golden_model_1.ACC [2]);
  nor (_36026_, _36025_, _36009_);
  nor (_36028_, _36026_, _06939_);
  nor (_36029_, _06938_, _36007_);
  or (_36030_, _36029_, _06102_);
  or (_36031_, _36030_, _36028_);
  and (_36032_, _36031_, _06848_);
  and (_36033_, _36032_, _36024_);
  nor (_36034_, _36020_, _06848_);
  or (_36035_, _36034_, _36033_);
  nand (_36036_, _36035_, _06220_);
  or (_36037_, _36026_, _06220_);
  and (_36039_, _36037_, _09817_);
  nand (_36040_, _36039_, _36036_);
  and (_36041_, _36040_, _36021_);
  and (_36042_, _36041_, _36018_);
  or (_36043_, _36042_, _09833_);
  and (_36044_, _14580_, _07681_);
  or (_36045_, _36044_, _36009_);
  or (_36046_, _36045_, _05669_);
  and (_36047_, _36046_, _06020_);
  and (_36048_, _36047_, _36043_);
  and (_36050_, _36012_, _06019_);
  or (_36051_, _36050_, _06112_);
  or (_36052_, _36051_, _36048_);
  and (_36053_, _14596_, _07681_);
  or (_36054_, _36009_, _08751_);
  or (_36055_, _36054_, _36053_);
  and (_36056_, _36055_, _08756_);
  and (_36057_, _36056_, _36052_);
  and (_36058_, _10991_, _07681_);
  or (_36059_, _36058_, _36009_);
  and (_36061_, _36059_, _06284_);
  or (_36062_, _36061_, _36057_);
  and (_36063_, _36062_, _07032_);
  or (_36064_, _36063_, _36014_);
  and (_36065_, _36064_, _06278_);
  nor (_36066_, _36026_, _06278_);
  and (_36067_, _36066_, _36010_);
  or (_36068_, _36067_, _06130_);
  or (_36069_, _36068_, _36065_);
  and (_36070_, _14593_, _07681_);
  or (_36072_, _36009_, _08777_);
  or (_36073_, _36072_, _36070_);
  and (_36074_, _36073_, _08782_);
  and (_36075_, _36074_, _36069_);
  nor (_36076_, _10990_, _13650_);
  or (_36077_, _36076_, _36009_);
  and (_36078_, _36077_, _06292_);
  or (_36079_, _36078_, _36075_);
  and (_36080_, _36079_, _06718_);
  and (_36081_, _36023_, _06316_);
  or (_36083_, _36081_, _06047_);
  or (_36084_, _36083_, _36080_);
  and (_36085_, _14657_, _07681_);
  or (_36086_, _36009_, _06048_);
  or (_36087_, _36086_, _36085_);
  and (_36088_, _36087_, _01336_);
  and (_36089_, _36088_, _36084_);
  or (_36090_, _36089_, _36008_);
  and (_43503_, _36090_, _42882_);
  and (_36091_, _01340_, \oc8051_golden_model_1.SBUF [3]);
  and (_36093_, _13650_, \oc8051_golden_model_1.SBUF [3]);
  and (_36094_, _07681_, _08662_);
  or (_36095_, _36094_, _36093_);
  or (_36096_, _36095_, _06020_);
  and (_36097_, _09181_, _07681_);
  or (_36098_, _36093_, _07012_);
  or (_36099_, _36098_, _36097_);
  and (_36100_, _14672_, _07681_);
  or (_36101_, _36100_, _36093_);
  or (_36102_, _36101_, _06954_);
  and (_36104_, _07681_, \oc8051_golden_model_1.ACC [3]);
  or (_36105_, _36104_, _36093_);
  and (_36106_, _36105_, _06938_);
  and (_36107_, _06939_, \oc8051_golden_model_1.SBUF [3]);
  or (_36108_, _36107_, _06102_);
  or (_36109_, _36108_, _36106_);
  and (_36110_, _36109_, _06848_);
  and (_36111_, _36110_, _36102_);
  nor (_36112_, _13650_, _07353_);
  or (_36113_, _36112_, _36093_);
  and (_36115_, _36113_, _06239_);
  or (_36116_, _36115_, _36111_);
  and (_36117_, _36116_, _06220_);
  and (_36118_, _36105_, _06219_);
  or (_36119_, _36118_, _09818_);
  or (_36120_, _36119_, _36117_);
  or (_36121_, _36113_, _09827_);
  and (_36122_, _36121_, _05669_);
  and (_36123_, _36122_, _36120_);
  and (_36124_, _36123_, _36099_);
  and (_36126_, _14778_, _07681_);
  or (_36127_, _36126_, _36093_);
  and (_36128_, _36127_, _09833_);
  or (_36129_, _36128_, _06019_);
  or (_36130_, _36129_, _36124_);
  and (_36131_, _36130_, _36096_);
  or (_36132_, _36131_, _06112_);
  and (_36133_, _14793_, _07681_);
  or (_36134_, _36133_, _36093_);
  or (_36135_, _36134_, _08751_);
  and (_36137_, _36135_, _08756_);
  and (_36138_, _36137_, _36132_);
  and (_36139_, _12299_, _07681_);
  or (_36140_, _36139_, _36093_);
  and (_36141_, _36140_, _06284_);
  or (_36142_, _36141_, _36138_);
  and (_36143_, _36142_, _07032_);
  or (_36144_, _36093_, _08029_);
  and (_36145_, _36095_, _06108_);
  and (_36146_, _36145_, _36144_);
  or (_36148_, _36146_, _36143_);
  and (_36149_, _36148_, _06278_);
  and (_36150_, _36105_, _06277_);
  and (_36151_, _36150_, _36144_);
  or (_36152_, _36151_, _06130_);
  or (_36153_, _36152_, _36149_);
  and (_36154_, _14792_, _07681_);
  or (_36155_, _36093_, _08777_);
  or (_36156_, _36155_, _36154_);
  and (_36157_, _36156_, _08782_);
  and (_36159_, _36157_, _36153_);
  nor (_36160_, _10988_, _13650_);
  or (_36161_, _36160_, _36093_);
  and (_36162_, _36161_, _06292_);
  or (_36163_, _36162_, _36159_);
  and (_36164_, _36163_, _06718_);
  and (_36165_, _36101_, _06316_);
  or (_36166_, _36165_, _06047_);
  or (_36167_, _36166_, _36164_);
  and (_36168_, _14849_, _07681_);
  or (_36170_, _36093_, _06048_);
  or (_36171_, _36170_, _36168_);
  and (_36172_, _36171_, _01336_);
  and (_36173_, _36172_, _36167_);
  or (_36174_, _36173_, _36091_);
  and (_43505_, _36174_, _42882_);
  and (_36175_, _01340_, \oc8051_golden_model_1.SBUF [4]);
  and (_36176_, _13650_, \oc8051_golden_model_1.SBUF [4]);
  or (_36177_, _36176_, _08273_);
  and (_36178_, _08665_, _07681_);
  or (_36180_, _36178_, _36176_);
  and (_36181_, _36180_, _06108_);
  and (_36182_, _36181_, _36177_);
  and (_36183_, _14887_, _07681_);
  or (_36184_, _36183_, _36176_);
  or (_36185_, _36184_, _06954_);
  and (_36186_, _07681_, \oc8051_golden_model_1.ACC [4]);
  or (_36187_, _36186_, _36176_);
  and (_36188_, _36187_, _06938_);
  and (_36189_, _06939_, \oc8051_golden_model_1.SBUF [4]);
  or (_36191_, _36189_, _06102_);
  or (_36192_, _36191_, _36188_);
  and (_36193_, _36192_, _06848_);
  and (_36194_, _36193_, _36185_);
  nor (_36195_, _08270_, _13650_);
  or (_36196_, _36195_, _36176_);
  and (_36197_, _36196_, _06239_);
  or (_36198_, _36197_, _36194_);
  and (_36199_, _36198_, _06220_);
  and (_36200_, _36187_, _06219_);
  or (_36202_, _36200_, _09815_);
  or (_36203_, _36202_, _36199_);
  or (_36204_, _36196_, _09827_);
  and (_36205_, _36204_, _07012_);
  and (_36206_, _36205_, _36203_);
  and (_36207_, _09180_, _07681_);
  or (_36208_, _36207_, _36176_);
  and (_36209_, _36208_, _07011_);
  or (_36210_, _36209_, _09833_);
  or (_36211_, _36210_, _36206_);
  and (_36213_, _14983_, _07681_);
  or (_36214_, _36176_, _05669_);
  or (_36215_, _36214_, _36213_);
  and (_36216_, _36215_, _06020_);
  and (_36217_, _36216_, _36211_);
  and (_36218_, _36180_, _06019_);
  or (_36219_, _36218_, _06112_);
  or (_36220_, _36219_, _36217_);
  and (_36221_, _14876_, _07681_);
  or (_36222_, _36176_, _08751_);
  or (_36224_, _36222_, _36221_);
  and (_36225_, _36224_, _08756_);
  and (_36226_, _36225_, _36220_);
  and (_36227_, _10986_, _07681_);
  or (_36228_, _36227_, _36176_);
  and (_36229_, _36228_, _06284_);
  or (_36230_, _36229_, _36226_);
  and (_36231_, _36230_, _07032_);
  or (_36232_, _36231_, _36182_);
  and (_36233_, _36232_, _06278_);
  and (_36235_, _36187_, _06277_);
  and (_36236_, _36235_, _36177_);
  or (_36237_, _36236_, _06130_);
  or (_36238_, _36237_, _36233_);
  and (_36239_, _14873_, _07681_);
  or (_36240_, _36176_, _08777_);
  or (_36241_, _36240_, _36239_);
  and (_36242_, _36241_, _08782_);
  and (_36243_, _36242_, _36238_);
  nor (_36244_, _10985_, _13650_);
  or (_36246_, _36244_, _36176_);
  and (_36247_, _36246_, _06292_);
  or (_36248_, _36247_, _36243_);
  and (_36249_, _36248_, _06718_);
  and (_36250_, _36184_, _06316_);
  or (_36251_, _36250_, _06047_);
  or (_36252_, _36251_, _36249_);
  and (_36253_, _15055_, _07681_);
  or (_36254_, _36176_, _06048_);
  or (_36255_, _36254_, _36253_);
  and (_36257_, _36255_, _01336_);
  and (_36258_, _36257_, _36252_);
  or (_36259_, _36258_, _36175_);
  and (_43506_, _36259_, _42882_);
  and (_36260_, _01340_, \oc8051_golden_model_1.SBUF [5]);
  and (_36261_, _13650_, \oc8051_golden_model_1.SBUF [5]);
  or (_36262_, _36261_, _07980_);
  and (_36263_, _08652_, _07681_);
  or (_36264_, _36263_, _36261_);
  and (_36265_, _36264_, _06108_);
  and (_36267_, _36265_, _36262_);
  or (_36268_, _36264_, _06020_);
  and (_36269_, _15093_, _07681_);
  or (_36270_, _36269_, _36261_);
  or (_36271_, _36270_, _06954_);
  and (_36272_, _07681_, \oc8051_golden_model_1.ACC [5]);
  or (_36273_, _36272_, _36261_);
  and (_36274_, _36273_, _06938_);
  and (_36275_, _06939_, \oc8051_golden_model_1.SBUF [5]);
  or (_36276_, _36275_, _06102_);
  or (_36278_, _36276_, _36274_);
  and (_36279_, _36278_, _06848_);
  and (_36280_, _36279_, _36271_);
  nor (_36281_, _07977_, _13650_);
  or (_36282_, _36281_, _36261_);
  and (_36283_, _36282_, _06239_);
  or (_36284_, _36283_, _36280_);
  and (_36285_, _36284_, _06220_);
  and (_36286_, _36273_, _06219_);
  or (_36287_, _36286_, _09818_);
  or (_36289_, _36287_, _36285_);
  and (_36290_, _09179_, _07681_);
  or (_36291_, _36261_, _07012_);
  or (_36292_, _36291_, _36290_);
  or (_36293_, _36282_, _09827_);
  and (_36294_, _36293_, _05669_);
  and (_36295_, _36294_, _36292_);
  and (_36296_, _36295_, _36289_);
  and (_36297_, _15179_, _07681_);
  or (_36298_, _36297_, _36261_);
  and (_36300_, _36298_, _09833_);
  or (_36301_, _36300_, _06019_);
  or (_36302_, _36301_, _36296_);
  and (_36303_, _36302_, _36268_);
  or (_36304_, _36303_, _06112_);
  and (_36305_, _15195_, _07681_);
  or (_36306_, _36305_, _36261_);
  or (_36307_, _36306_, _08751_);
  and (_36308_, _36307_, _08756_);
  and (_36309_, _36308_, _36304_);
  and (_36311_, _12306_, _07681_);
  or (_36312_, _36311_, _36261_);
  and (_36313_, _36312_, _06284_);
  or (_36314_, _36313_, _36309_);
  and (_36315_, _36314_, _07032_);
  or (_36316_, _36315_, _36267_);
  and (_36317_, _36316_, _06278_);
  and (_36318_, _36273_, _06277_);
  and (_36319_, _36318_, _36262_);
  or (_36320_, _36319_, _06130_);
  or (_36322_, _36320_, _36317_);
  and (_36323_, _15194_, _07681_);
  or (_36324_, _36261_, _08777_);
  or (_36325_, _36324_, _36323_);
  and (_36326_, _36325_, _08782_);
  and (_36327_, _36326_, _36322_);
  nor (_36328_, _10982_, _13650_);
  or (_36329_, _36328_, _36261_);
  and (_36330_, _36329_, _06292_);
  or (_36331_, _36330_, _36327_);
  and (_36333_, _36331_, _06718_);
  and (_36334_, _36270_, _06316_);
  or (_36335_, _36334_, _06047_);
  or (_36336_, _36335_, _36333_);
  and (_36337_, _15253_, _07681_);
  or (_36338_, _36261_, _06048_);
  or (_36339_, _36338_, _36337_);
  and (_36340_, _36339_, _01336_);
  and (_36341_, _36340_, _36336_);
  or (_36342_, _36341_, _36260_);
  and (_43507_, _36342_, _42882_);
  and (_36344_, _01340_, \oc8051_golden_model_1.SBUF [6]);
  and (_36345_, _13650_, \oc8051_golden_model_1.SBUF [6]);
  and (_36346_, _15389_, _07681_);
  or (_36347_, _36346_, _36345_);
  or (_36348_, _36347_, _06020_);
  and (_36349_, _15293_, _07681_);
  or (_36350_, _36349_, _36345_);
  or (_36351_, _36350_, _06954_);
  and (_36352_, _07681_, \oc8051_golden_model_1.ACC [6]);
  or (_36354_, _36352_, _36345_);
  and (_36355_, _36354_, _06938_);
  and (_36356_, _06939_, \oc8051_golden_model_1.SBUF [6]);
  or (_36357_, _36356_, _06102_);
  or (_36358_, _36357_, _36355_);
  and (_36359_, _36358_, _06848_);
  and (_36360_, _36359_, _36351_);
  nor (_36361_, _07883_, _13650_);
  or (_36362_, _36361_, _36345_);
  and (_36363_, _36362_, _06239_);
  or (_36364_, _36363_, _36360_);
  and (_36365_, _36364_, _06220_);
  and (_36366_, _36354_, _06219_);
  or (_36367_, _36366_, _09818_);
  or (_36368_, _36367_, _36365_);
  and (_36369_, _09178_, _07681_);
  or (_36370_, _36345_, _07012_);
  or (_36371_, _36370_, _36369_);
  or (_36372_, _36362_, _09827_);
  and (_36373_, _36372_, _05669_);
  and (_36375_, _36373_, _36371_);
  and (_36376_, _36375_, _36368_);
  and (_36377_, _15382_, _07681_);
  or (_36378_, _36377_, _36345_);
  and (_36379_, _36378_, _09833_);
  or (_36380_, _36379_, _06019_);
  or (_36381_, _36380_, _36376_);
  and (_36382_, _36381_, _36348_);
  or (_36383_, _36382_, _06112_);
  and (_36384_, _15399_, _07681_);
  or (_36386_, _36384_, _36345_);
  or (_36387_, _36386_, _08751_);
  and (_36388_, _36387_, _08756_);
  and (_36389_, _36388_, _36383_);
  and (_36390_, _10980_, _07681_);
  or (_36391_, _36390_, _36345_);
  and (_36392_, _36391_, _06284_);
  or (_36393_, _36392_, _36389_);
  and (_36394_, _36393_, _07032_);
  or (_36395_, _36345_, _07886_);
  and (_36397_, _36347_, _06108_);
  and (_36398_, _36397_, _36395_);
  or (_36399_, _36398_, _36394_);
  and (_36400_, _36399_, _06278_);
  and (_36401_, _36354_, _06277_);
  and (_36402_, _36401_, _36395_);
  or (_36403_, _36402_, _06130_);
  or (_36404_, _36403_, _36400_);
  and (_36405_, _15396_, _07681_);
  or (_36406_, _36345_, _08777_);
  or (_36408_, _36406_, _36405_);
  and (_36409_, _36408_, _08782_);
  and (_36410_, _36409_, _36404_);
  nor (_36411_, _10979_, _13650_);
  or (_36412_, _36411_, _36345_);
  and (_36413_, _36412_, _06292_);
  or (_36414_, _36413_, _36410_);
  and (_36415_, _36414_, _06718_);
  and (_36416_, _36350_, _06316_);
  or (_36417_, _36416_, _06047_);
  or (_36419_, _36417_, _36415_);
  and (_36420_, _15451_, _07681_);
  or (_36421_, _36345_, _06048_);
  or (_36422_, _36421_, _36420_);
  and (_36423_, _36422_, _01336_);
  and (_36424_, _36423_, _36419_);
  or (_36425_, _36424_, _36344_);
  and (_43508_, _36425_, _42882_);
  not (_36426_, \oc8051_golden_model_1.PSW [0]);
  nor (_36427_, _01336_, _36426_);
  nand (_36429_, _10995_, _07705_);
  nor (_36430_, _07705_, _36426_);
  nor (_36431_, _36430_, _06278_);
  nand (_36432_, _36431_, _36429_);
  and (_36433_, _07705_, _08672_);
  or (_36434_, _36433_, _36430_);
  or (_36435_, _36434_, _06020_);
  and (_36436_, _09120_, _07705_);
  or (_36437_, _36430_, _07012_);
  or (_36438_, _36437_, _36436_);
  nor (_36440_, _08127_, _13745_);
  or (_36441_, _36440_, _36430_);
  or (_36442_, _36441_, _06954_);
  and (_36443_, _07705_, \oc8051_golden_model_1.ACC [0]);
  or (_36444_, _36443_, _36430_);
  and (_36445_, _36444_, _06938_);
  nor (_36446_, _06938_, _36426_);
  or (_36447_, _36446_, _06102_);
  or (_36448_, _36447_, _36445_);
  and (_36449_, _36448_, _06044_);
  and (_36451_, _36449_, _36442_);
  nor (_36452_, _08355_, _36426_);
  and (_36453_, _14102_, _08355_);
  or (_36454_, _36453_, _36452_);
  and (_36455_, _36454_, _06043_);
  or (_36456_, _36455_, _36451_);
  and (_36457_, _36456_, _06848_);
  and (_36458_, _07705_, _06931_);
  or (_36459_, _36458_, _36430_);
  and (_36460_, _36459_, _06239_);
  or (_36462_, _36460_, _06219_);
  or (_36463_, _36462_, _36457_);
  or (_36464_, _36444_, _06220_);
  and (_36465_, _36464_, _06040_);
  and (_36466_, _36465_, _36463_);
  and (_36467_, _36430_, _06039_);
  or (_36468_, _36467_, _06032_);
  or (_36469_, _36468_, _36466_);
  or (_36470_, _36441_, _06033_);
  and (_36471_, _36470_, _06027_);
  and (_36473_, _36471_, _36469_);
  or (_36474_, _36452_, _14131_);
  and (_36475_, _36474_, _06026_);
  and (_36476_, _36475_, _36454_);
  or (_36477_, _36476_, _09818_);
  or (_36478_, _36477_, _36473_);
  or (_36479_, _36459_, _09827_);
  and (_36480_, _36479_, _05669_);
  and (_36481_, _36480_, _36478_);
  and (_36482_, _36481_, _36438_);
  and (_36484_, _14186_, _07705_);
  or (_36485_, _36484_, _36430_);
  and (_36486_, _36485_, _09833_);
  or (_36487_, _36486_, _06019_);
  or (_36488_, _36487_, _36482_);
  and (_36489_, _36488_, _36435_);
  or (_36490_, _36489_, _06112_);
  and (_36491_, _14086_, _07705_);
  or (_36492_, _36491_, _36430_);
  or (_36493_, _36492_, _08751_);
  and (_36495_, _36493_, _08756_);
  and (_36496_, _36495_, _36490_);
  nor (_36497_, _12302_, _13745_);
  or (_36498_, _36497_, _36430_);
  and (_36499_, _36429_, _06284_);
  and (_36500_, _36499_, _36498_);
  or (_36501_, _36500_, _36496_);
  and (_36502_, _36501_, _07032_);
  nand (_36503_, _36434_, _06108_);
  nor (_36504_, _36503_, _36440_);
  or (_36506_, _36504_, _06277_);
  or (_36507_, _36506_, _36502_);
  and (_36508_, _36507_, _36432_);
  or (_36509_, _36508_, _06130_);
  and (_36510_, _14083_, _07705_);
  or (_36511_, _36430_, _08777_);
  or (_36512_, _36511_, _36510_);
  and (_36513_, _36512_, _08782_);
  and (_36514_, _36513_, _36509_);
  and (_36515_, _36498_, _06292_);
  or (_36517_, _36515_, _06316_);
  or (_36518_, _36517_, _36514_);
  or (_36519_, _36441_, _06718_);
  and (_36520_, _36519_, _36518_);
  or (_36521_, _36520_, _05652_);
  or (_36522_, _36430_, _05653_);
  and (_36523_, _36522_, _36521_);
  or (_36524_, _36523_, _06047_);
  or (_36525_, _36441_, _06048_);
  and (_36526_, _36525_, _01336_);
  and (_36528_, _36526_, _36524_);
  or (_36529_, _36528_, _36427_);
  and (_43510_, _36529_, _42882_);
  not (_36530_, \oc8051_golden_model_1.PSW [1]);
  nor (_36531_, _01336_, _36530_);
  nor (_36532_, _07705_, _36530_);
  nor (_36533_, _10993_, _13745_);
  or (_36534_, _36533_, _36532_);
  or (_36535_, _36534_, _08782_);
  or (_36536_, _14367_, _13745_);
  or (_36538_, _07705_, \oc8051_golden_model_1.PSW [1]);
  and (_36539_, _36538_, _09833_);
  and (_36540_, _36539_, _36536_);
  and (_36541_, _09075_, _07705_);
  or (_36542_, _36541_, _36532_);
  and (_36543_, _36542_, _07011_);
  nor (_36544_, _13745_, _07132_);
  or (_36545_, _36544_, _36532_);
  and (_36546_, _36545_, _06239_);
  nor (_36547_, _08355_, _36530_);
  and (_36549_, _14266_, _08355_);
  or (_36550_, _36549_, _36547_);
  or (_36551_, _36550_, _06044_);
  and (_36552_, _14284_, _07705_);
  not (_36553_, _36552_);
  and (_36554_, _36553_, _36538_);
  and (_36555_, _36554_, _06102_);
  nor (_36556_, _06938_, _36530_);
  and (_36557_, _07705_, \oc8051_golden_model_1.ACC [1]);
  or (_36558_, _36557_, _36532_);
  and (_36560_, _36558_, _06938_);
  or (_36561_, _36560_, _36556_);
  and (_36562_, _36561_, _06954_);
  or (_36563_, _36562_, _06043_);
  or (_36564_, _36563_, _36555_);
  and (_36565_, _36564_, _36551_);
  and (_36566_, _36565_, _06848_);
  or (_36567_, _36566_, _36546_);
  or (_36568_, _36567_, _06219_);
  or (_36569_, _36558_, _06220_);
  and (_36571_, _36569_, _06040_);
  and (_36572_, _36571_, _36568_);
  and (_36573_, _14273_, _08355_);
  or (_36574_, _36573_, _36547_);
  and (_36575_, _36574_, _06039_);
  or (_36576_, _36575_, _06032_);
  or (_36577_, _36576_, _36572_);
  or (_36578_, _36547_, _14302_);
  and (_36579_, _36578_, _36550_);
  or (_36580_, _36579_, _06033_);
  and (_36582_, _36580_, _06027_);
  and (_36583_, _36582_, _36577_);
  or (_36584_, _36547_, _14267_);
  and (_36585_, _36584_, _06026_);
  and (_36586_, _36585_, _36550_);
  or (_36587_, _36586_, _09815_);
  or (_36588_, _36587_, _36583_);
  or (_36589_, _36545_, _09827_);
  and (_36590_, _36589_, _07012_);
  and (_36591_, _36590_, _36588_);
  or (_36593_, _36591_, _36543_);
  and (_36594_, _36593_, _05669_);
  or (_36595_, _36594_, _36540_);
  and (_36596_, _36595_, _06020_);
  nand (_36597_, _07705_, _06832_);
  and (_36598_, _36538_, _06019_);
  and (_36599_, _36598_, _36597_);
  or (_36600_, _36599_, _36596_);
  and (_36601_, _36600_, _08751_);
  or (_36602_, _14263_, _13745_);
  and (_36604_, _36538_, _06112_);
  and (_36605_, _36604_, _36602_);
  or (_36606_, _36605_, _06284_);
  or (_36607_, _36606_, _36601_);
  nand (_36608_, _10992_, _07705_);
  and (_36609_, _36608_, _36534_);
  or (_36610_, _36609_, _08756_);
  and (_36611_, _36610_, _07032_);
  and (_36612_, _36611_, _36607_);
  or (_36613_, _14261_, _13745_);
  and (_36615_, _36538_, _06108_);
  and (_36616_, _36615_, _36613_);
  or (_36617_, _36616_, _06277_);
  or (_36618_, _36617_, _36612_);
  nor (_36619_, _36532_, _06278_);
  nand (_36620_, _36619_, _36608_);
  and (_36621_, _36620_, _08777_);
  and (_36622_, _36621_, _36618_);
  or (_36623_, _36597_, _08078_);
  and (_36624_, _36538_, _06130_);
  and (_36626_, _36624_, _36623_);
  or (_36627_, _36626_, _06292_);
  or (_36628_, _36627_, _36622_);
  and (_36629_, _36628_, _36535_);
  or (_36630_, _36629_, _06316_);
  or (_36631_, _36554_, _06718_);
  and (_36632_, _36631_, _05653_);
  and (_36633_, _36632_, _36630_);
  and (_36634_, _36574_, _05652_);
  or (_36635_, _36634_, _06047_);
  or (_36637_, _36635_, _36633_);
  or (_36638_, _36532_, _06048_);
  or (_36639_, _36638_, _36552_);
  and (_36640_, _36639_, _01336_);
  and (_36641_, _36640_, _36637_);
  or (_36642_, _36641_, _36531_);
  and (_43511_, _36642_, _42882_);
  not (_36643_, \oc8051_golden_model_1.PSW [2]);
  nor (_36644_, _01336_, _36643_);
  not (_36645_, _10692_);
  nand (_36647_, _10967_, _36645_);
  or (_36648_, _10967_, _10691_);
  and (_36649_, _36648_, _36647_);
  and (_36650_, _36649_, _06692_);
  nor (_36651_, _10570_, _13739_);
  not (_36652_, _36651_);
  nor (_36653_, _10570_, _06053_);
  or (_36654_, _36653_, \oc8051_golden_model_1.ACC [7]);
  and (_36655_, _36654_, _36652_);
  not (_36656_, _36655_);
  or (_36658_, _36656_, _14017_);
  and (_36659_, _36658_, _10880_);
  or (_36660_, _36659_, _36651_);
  or (_36661_, _36652_, _10877_);
  and (_36662_, _36661_, _10824_);
  and (_36663_, _36662_, _36660_);
  and (_36664_, _09182_, _07705_);
  nor (_36665_, _07705_, _36643_);
  or (_36666_, _36665_, _07012_);
  or (_36667_, _36666_, _36664_);
  nor (_36669_, _13745_, _07530_);
  or (_36670_, _36669_, _36665_);
  or (_36671_, _36670_, _09827_);
  nor (_36672_, _10496_, \oc8051_golden_model_1.ACC [7]);
  nor (_36673_, _10495_, _36645_);
  nor (_36674_, _36673_, _36672_);
  nor (_36675_, _36674_, _10501_);
  nor (_36676_, _13934_, _10497_);
  nor (_36677_, _36676_, _36675_);
  and (_36678_, _36677_, _10556_);
  nor (_36680_, _36677_, _10556_);
  or (_36681_, _36680_, _36678_);
  and (_36682_, _36681_, _12361_);
  nor (_36683_, _08355_, _36643_);
  and (_36684_, _14479_, _08355_);
  or (_36685_, _36684_, _36683_);
  and (_36686_, _36685_, _06039_);
  or (_36687_, _36670_, _06848_);
  and (_36688_, _14493_, _07705_);
  or (_36689_, _36688_, _36665_);
  or (_36691_, _36689_, _06954_);
  and (_36692_, _07705_, \oc8051_golden_model_1.ACC [2]);
  or (_36693_, _36692_, _36665_);
  and (_36694_, _36693_, _06938_);
  nor (_36695_, _06938_, _36643_);
  or (_36696_, _36695_, _06102_);
  or (_36697_, _36696_, _36694_);
  and (_36698_, _36697_, _06044_);
  and (_36699_, _36698_, _36691_);
  and (_36700_, _14497_, _08355_);
  or (_36702_, _36700_, _36683_);
  and (_36703_, _36702_, _06043_);
  or (_36704_, _36703_, _06239_);
  or (_36705_, _36704_, _36699_);
  and (_36706_, _36705_, _36687_);
  or (_36707_, _36706_, _06219_);
  or (_36708_, _36693_, _06220_);
  and (_36709_, _36708_, _06040_);
  and (_36710_, _36709_, _36707_);
  or (_36711_, _36710_, _36686_);
  and (_36713_, _36711_, _06033_);
  and (_36714_, _36700_, _14512_);
  or (_36715_, _36714_, _36683_);
  and (_36716_, _36715_, _06032_);
  or (_36717_, _36716_, _36713_);
  and (_36718_, _36717_, _09800_);
  or (_36719_, _16187_, _09803_);
  or (_36720_, _36719_, _16295_);
  or (_36721_, _36720_, _16411_);
  or (_36722_, _36721_, _16527_);
  or (_36724_, _36722_, _16643_);
  or (_36725_, _36724_, _16757_);
  or (_36726_, _36725_, _16877_);
  and (_36727_, _36726_, _09269_);
  or (_36728_, _36727_, _10468_);
  or (_36729_, _36728_, _36718_);
  nor (_36730_, _10719_, _10240_);
  or (_36731_, _10240_, _07785_);
  and (_36732_, _36731_, _08393_);
  or (_36733_, _36732_, _36730_);
  and (_36735_, _36733_, _13925_);
  nor (_36736_, _36733_, _13925_);
  nor (_36737_, _36736_, _36735_);
  not (_36738_, _36737_);
  nor (_36739_, _36738_, _10490_);
  and (_36740_, _36738_, _10490_);
  or (_36741_, _36740_, _36739_);
  or (_36742_, _36741_, _10469_);
  and (_36743_, _36742_, _13935_);
  and (_36744_, _36743_, _36729_);
  or (_36746_, _36744_, _36682_);
  and (_36747_, _36746_, _06267_);
  nor (_36748_, _10314_, _14043_);
  nor (_36749_, _10315_, \oc8051_golden_model_1.ACC [7]);
  nor (_36750_, _36749_, _36748_);
  nor (_36751_, _36750_, _10320_);
  nor (_36752_, _13761_, _10316_);
  or (_36753_, _36752_, _36751_);
  nand (_36754_, _36753_, _10370_);
  or (_36755_, _36753_, _10370_);
  and (_36757_, _36755_, _06261_);
  and (_36758_, _36757_, _36754_);
  or (_36759_, _36758_, _10306_);
  or (_36760_, _36759_, _36747_);
  nor (_36761_, _36655_, _13947_);
  and (_36762_, _36655_, _13947_);
  nor (_36763_, _36762_, _36761_);
  and (_36764_, _36763_, _10631_);
  nor (_36765_, _36763_, _10631_);
  or (_36766_, _36765_, _36764_);
  or (_36768_, _36766_, _10307_);
  and (_36769_, _36768_, _06027_);
  and (_36770_, _36769_, _36760_);
  or (_36771_, _36683_, _14525_);
  and (_36772_, _36771_, _06026_);
  and (_36773_, _36772_, _36702_);
  or (_36774_, _36773_, _09815_);
  or (_36775_, _36774_, _36770_);
  and (_36776_, _36775_, _36671_);
  or (_36777_, _36776_, _07011_);
  and (_36779_, _36777_, _36667_);
  or (_36780_, _36779_, _09833_);
  and (_36781_, _14580_, _07705_);
  or (_36782_, _36665_, _05669_);
  or (_36783_, _36782_, _36781_);
  and (_36784_, _36783_, _09839_);
  and (_36785_, _36784_, _36780_);
  nor (_36786_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and (_36787_, _36786_, _09832_);
  and (_36788_, _36787_, _09860_);
  or (_36790_, _36788_, _06019_);
  or (_36791_, _36790_, _36785_);
  and (_36792_, _07705_, _08730_);
  or (_36793_, _36792_, _36665_);
  or (_36794_, _36793_, _06020_);
  and (_36795_, _36794_, _36791_);
  or (_36796_, _36795_, _06112_);
  and (_36797_, _14596_, _07705_);
  or (_36798_, _36797_, _36665_);
  or (_36799_, _36798_, _08751_);
  and (_36801_, _36799_, _08756_);
  and (_36802_, _36801_, _36796_);
  and (_36803_, _10991_, _07705_);
  or (_36804_, _36803_, _36665_);
  and (_36805_, _36804_, _06284_);
  or (_36806_, _36805_, _36802_);
  and (_36807_, _36806_, _07032_);
  or (_36808_, _36665_, _08177_);
  and (_36809_, _36793_, _06108_);
  and (_36810_, _36809_, _36808_);
  or (_36812_, _36810_, _36807_);
  and (_36813_, _36812_, _06278_);
  and (_36814_, _36693_, _06277_);
  and (_36815_, _36814_, _36808_);
  or (_36816_, _36815_, _06130_);
  or (_36817_, _36816_, _36813_);
  and (_36818_, _14593_, _07705_);
  or (_36819_, _36665_, _08777_);
  or (_36820_, _36819_, _36818_);
  and (_36821_, _36820_, _08782_);
  and (_36823_, _36821_, _36817_);
  nor (_36824_, _10990_, _13745_);
  or (_36825_, _36824_, _36665_);
  and (_36826_, _36825_, _06292_);
  or (_36827_, _36826_, _10303_);
  or (_36828_, _36827_, _36823_);
  nor (_36829_, _36733_, _13999_);
  nor (_36830_, _36829_, _36730_);
  and (_36831_, _36830_, _10302_);
  and (_36832_, _36730_, _10299_);
  or (_36834_, _36832_, _10304_);
  or (_36835_, _36834_, _36831_);
  and (_36836_, _36835_, _17410_);
  and (_36837_, _36836_, _36828_);
  not (_36838_, _36674_);
  nor (_36839_, _36838_, _14006_);
  nor (_36840_, _36839_, _36673_);
  and (_36841_, _36840_, _10820_);
  and (_36842_, _36673_, _10817_);
  or (_36843_, _36842_, _36841_);
  and (_36845_, _36843_, _17409_);
  or (_36846_, _36845_, _36837_);
  and (_36847_, _36846_, _17423_);
  nand (_36848_, _36843_, _17416_);
  nand (_36849_, _36848_, _06289_);
  or (_36850_, _36849_, _36847_);
  nor (_36851_, _36749_, _14011_);
  nor (_36852_, _36851_, _36748_);
  and (_36853_, _36852_, _10850_);
  and (_36854_, _36748_, _10847_);
  or (_36856_, _36854_, _36853_);
  or (_36857_, _36856_, _06289_);
  and (_36858_, _36857_, _10856_);
  and (_36859_, _36858_, _36850_);
  or (_36860_, _36859_, _36663_);
  and (_36861_, _36860_, _10890_);
  nand (_36862_, _10926_, _10719_);
  and (_36863_, _36862_, _16956_);
  and (_36864_, _36863_, _14027_);
  or (_36865_, _36864_, _17437_);
  or (_36867_, _36865_, _36861_);
  and (_36868_, _36649_, _17443_);
  or (_36869_, _36868_, _10934_);
  and (_36870_, _36869_, _36867_);
  or (_36871_, _36870_, _36650_);
  and (_36872_, _36871_, _10975_);
  or (_36873_, _11008_, _08767_);
  and (_36874_, _14045_, _36873_);
  nand (_36875_, _11048_, _13739_);
  and (_36876_, _36875_, _13741_);
  or (_36878_, _36876_, _06316_);
  or (_36879_, _36878_, _36874_);
  or (_36880_, _36879_, _36872_);
  or (_36881_, _36689_, _06718_);
  and (_36882_, _36881_, _05653_);
  and (_36883_, _36882_, _36880_);
  and (_36884_, _36685_, _05652_);
  or (_36885_, _36884_, _06047_);
  or (_36886_, _36885_, _36883_);
  and (_36887_, _14657_, _07705_);
  or (_36889_, _36665_, _06048_);
  or (_36890_, _36889_, _36887_);
  and (_36891_, _36890_, _01336_);
  and (_36892_, _36891_, _36886_);
  or (_36893_, _36892_, _36644_);
  and (_43512_, _36893_, _42882_);
  nor (_36894_, _01336_, _07369_);
  nor (_36895_, _07705_, _07369_);
  nor (_36896_, _13745_, _07353_);
  or (_36897_, _36896_, _36895_);
  or (_36899_, _36897_, _09827_);
  nor (_36900_, _08355_, _07369_);
  and (_36901_, _14681_, _08355_);
  or (_36902_, _36901_, _36900_);
  and (_36903_, _36902_, _06039_);
  and (_36904_, _14672_, _07705_);
  or (_36905_, _36904_, _36895_);
  or (_36906_, _36905_, _06954_);
  and (_36907_, _07705_, \oc8051_golden_model_1.ACC [3]);
  or (_36908_, _36907_, _36895_);
  and (_36910_, _36908_, _06938_);
  nor (_36911_, _06938_, _07369_);
  or (_36912_, _36911_, _06102_);
  or (_36913_, _36912_, _36910_);
  and (_36914_, _36913_, _06044_);
  and (_36915_, _36914_, _36906_);
  and (_36916_, _14683_, _08355_);
  or (_36917_, _36916_, _36900_);
  and (_36918_, _36917_, _06043_);
  or (_36919_, _36918_, _06239_);
  or (_36921_, _36919_, _36915_);
  or (_36922_, _36897_, _06848_);
  and (_36923_, _36922_, _36921_);
  or (_36924_, _36923_, _06219_);
  or (_36925_, _36908_, _06220_);
  and (_36926_, _36925_, _06040_);
  and (_36927_, _36926_, _36924_);
  or (_36928_, _36927_, _36903_);
  and (_36929_, _36928_, _06033_);
  and (_36930_, _14709_, _08355_);
  or (_36932_, _36930_, _36900_);
  and (_36933_, _36932_, _06032_);
  or (_36934_, _36933_, _36929_);
  and (_36935_, _36934_, _06027_);
  and (_36936_, _14724_, _08355_);
  or (_36937_, _36936_, _36900_);
  and (_36938_, _36937_, _06026_);
  or (_36939_, _36938_, _09815_);
  or (_36940_, _36939_, _36935_);
  and (_36941_, _36940_, _36899_);
  or (_36943_, _36941_, _07011_);
  and (_36944_, _09181_, _07705_);
  or (_36945_, _36895_, _07012_);
  or (_36946_, _36945_, _36944_);
  and (_36947_, _36946_, _36943_);
  or (_36948_, _36947_, _09833_);
  and (_36949_, _14778_, _07705_);
  or (_36950_, _36949_, _36895_);
  or (_36951_, _36950_, _05669_);
  and (_36952_, _36951_, _06020_);
  and (_36954_, _36952_, _36948_);
  and (_36955_, _07705_, _08662_);
  or (_36956_, _36955_, _36895_);
  and (_36957_, _36956_, _06019_);
  or (_36958_, _36957_, _06112_);
  or (_36959_, _36958_, _36954_);
  and (_36960_, _14793_, _07705_);
  or (_36961_, _36960_, _36895_);
  or (_36962_, _36961_, _08751_);
  and (_36963_, _36962_, _08756_);
  and (_36965_, _36963_, _36959_);
  and (_36966_, _12299_, _07705_);
  or (_36967_, _36966_, _36895_);
  and (_36968_, _36967_, _06284_);
  or (_36969_, _36968_, _36965_);
  and (_36970_, _36969_, _07032_);
  or (_36971_, _36895_, _08029_);
  and (_36972_, _36956_, _06108_);
  and (_36973_, _36972_, _36971_);
  or (_36974_, _36973_, _36970_);
  and (_36976_, _36974_, _06278_);
  and (_36977_, _36908_, _06277_);
  and (_36978_, _36977_, _36971_);
  or (_36979_, _36978_, _06130_);
  or (_36980_, _36979_, _36976_);
  and (_36981_, _14792_, _07705_);
  or (_36982_, _36895_, _08777_);
  or (_36983_, _36982_, _36981_);
  and (_36984_, _36983_, _08782_);
  and (_36985_, _36984_, _36980_);
  nor (_36987_, _10988_, _13745_);
  or (_36988_, _36987_, _36895_);
  and (_36989_, _36988_, _06292_);
  or (_36990_, _36989_, _06316_);
  or (_36991_, _36990_, _36985_);
  or (_36992_, _36905_, _06718_);
  and (_36993_, _36992_, _05653_);
  and (_36994_, _36993_, _36991_);
  and (_36995_, _36902_, _05652_);
  or (_36996_, _36995_, _06047_);
  or (_36998_, _36996_, _36994_);
  and (_36999_, _14849_, _07705_);
  or (_37000_, _36895_, _06048_);
  or (_37001_, _37000_, _36999_);
  and (_37002_, _37001_, _01336_);
  and (_37003_, _37002_, _36998_);
  or (_37004_, _37003_, _36894_);
  and (_43513_, _37004_, _42882_);
  not (_37005_, \oc8051_golden_model_1.PSW [4]);
  nor (_37006_, _01336_, _37005_);
  nor (_37008_, _07705_, _37005_);
  nor (_37009_, _08270_, _13745_);
  or (_37010_, _37009_, _37008_);
  or (_37011_, _37010_, _09827_);
  nor (_37012_, _08355_, _37005_);
  and (_37013_, _14882_, _08355_);
  or (_37014_, _37013_, _37012_);
  and (_37015_, _37014_, _06039_);
  and (_37016_, _14887_, _07705_);
  or (_37017_, _37016_, _37008_);
  or (_37019_, _37017_, _06954_);
  and (_37020_, _07705_, \oc8051_golden_model_1.ACC [4]);
  or (_37021_, _37020_, _37008_);
  and (_37022_, _37021_, _06938_);
  nor (_37023_, _06938_, _37005_);
  or (_37024_, _37023_, _06102_);
  or (_37025_, _37024_, _37022_);
  and (_37026_, _37025_, _06044_);
  and (_37027_, _37026_, _37019_);
  and (_37028_, _14878_, _08355_);
  or (_37030_, _37028_, _37012_);
  and (_37031_, _37030_, _06043_);
  or (_37032_, _37031_, _06239_);
  or (_37033_, _37032_, _37027_);
  or (_37034_, _37010_, _06848_);
  and (_37035_, _37034_, _37033_);
  or (_37036_, _37035_, _06219_);
  or (_37037_, _37021_, _06220_);
  and (_37038_, _37037_, _06040_);
  and (_37039_, _37038_, _37036_);
  or (_37041_, _37039_, _37015_);
  and (_37042_, _37041_, _06033_);
  and (_37043_, _14915_, _08355_);
  or (_37044_, _37043_, _37012_);
  and (_37045_, _37044_, _06032_);
  or (_37046_, _37045_, _37042_);
  and (_37047_, _37046_, _06027_);
  or (_37048_, _37012_, _14879_);
  and (_37049_, _37048_, _06026_);
  and (_37050_, _37049_, _37030_);
  or (_37052_, _37050_, _09815_);
  or (_37053_, _37052_, _37047_);
  and (_37054_, _37053_, _37011_);
  or (_37055_, _37054_, _07011_);
  and (_37056_, _09180_, _07705_);
  or (_37057_, _37008_, _07012_);
  or (_37058_, _37057_, _37056_);
  and (_37059_, _37058_, _37055_);
  or (_37060_, _37059_, _09833_);
  and (_37061_, _14983_, _07705_);
  or (_37063_, _37061_, _37008_);
  or (_37064_, _37063_, _05669_);
  and (_37065_, _37064_, _06020_);
  and (_37066_, _37065_, _37060_);
  and (_37067_, _08665_, _07705_);
  or (_37068_, _37067_, _37008_);
  and (_37069_, _37068_, _06019_);
  or (_37070_, _37069_, _06112_);
  or (_37071_, _37070_, _37066_);
  and (_37072_, _14876_, _07705_);
  or (_37074_, _37008_, _08751_);
  or (_37075_, _37074_, _37072_);
  and (_37076_, _37075_, _08756_);
  and (_37077_, _37076_, _37071_);
  and (_37078_, _10986_, _07705_);
  or (_37079_, _37078_, _37008_);
  and (_37080_, _37079_, _06284_);
  or (_37081_, _37080_, _37077_);
  and (_37082_, _37081_, _07032_);
  or (_37083_, _37008_, _08273_);
  and (_37085_, _37068_, _06108_);
  and (_37086_, _37085_, _37083_);
  or (_37087_, _37086_, _37082_);
  and (_37088_, _37087_, _06278_);
  and (_37089_, _37021_, _06277_);
  and (_37090_, _37089_, _37083_);
  or (_37091_, _37090_, _06130_);
  or (_37092_, _37091_, _37088_);
  and (_37093_, _14873_, _07705_);
  or (_37094_, _37008_, _08777_);
  or (_37096_, _37094_, _37093_);
  and (_37097_, _37096_, _08782_);
  and (_37098_, _37097_, _37092_);
  nor (_37099_, _10985_, _13745_);
  or (_37100_, _37099_, _37008_);
  and (_37101_, _37100_, _06292_);
  or (_37102_, _37101_, _06316_);
  or (_37103_, _37102_, _37098_);
  or (_37104_, _37017_, _06718_);
  and (_37105_, _37104_, _05653_);
  and (_37107_, _37105_, _37103_);
  and (_37108_, _37014_, _05652_);
  or (_37109_, _37108_, _06047_);
  or (_37110_, _37109_, _37107_);
  and (_37111_, _15055_, _07705_);
  or (_37112_, _37008_, _06048_);
  or (_37113_, _37112_, _37111_);
  and (_37114_, _37113_, _01336_);
  and (_37115_, _37114_, _37110_);
  or (_37116_, _37115_, _37006_);
  and (_43514_, _37116_, _42882_);
  not (_37118_, \oc8051_golden_model_1.PSW [5]);
  nor (_37119_, _01336_, _37118_);
  nor (_37120_, _07705_, _37118_);
  nor (_37121_, _07977_, _13745_);
  or (_37122_, _37121_, _37120_);
  or (_37123_, _37122_, _09827_);
  and (_37124_, _15093_, _07705_);
  or (_37125_, _37124_, _37120_);
  or (_37126_, _37125_, _06954_);
  and (_37128_, _07705_, \oc8051_golden_model_1.ACC [5]);
  or (_37129_, _37128_, _37120_);
  and (_37130_, _37129_, _06938_);
  nor (_37131_, _06938_, _37118_);
  or (_37132_, _37131_, _06102_);
  or (_37133_, _37132_, _37130_);
  and (_37134_, _37133_, _06044_);
  and (_37135_, _37134_, _37126_);
  nor (_37136_, _08355_, _37118_);
  and (_37137_, _15073_, _08355_);
  or (_37139_, _37137_, _37136_);
  and (_37140_, _37139_, _06043_);
  or (_37141_, _37140_, _06239_);
  or (_37142_, _37141_, _37135_);
  or (_37143_, _37122_, _06848_);
  and (_37144_, _37143_, _37142_);
  or (_37145_, _37144_, _06219_);
  or (_37146_, _37129_, _06220_);
  and (_37147_, _37146_, _06040_);
  and (_37148_, _37147_, _37145_);
  and (_37150_, _15077_, _08355_);
  or (_37151_, _37150_, _37136_);
  and (_37152_, _37151_, _06039_);
  or (_37153_, _37152_, _06032_);
  or (_37154_, _37153_, _37148_);
  or (_37155_, _37136_, _15110_);
  and (_37156_, _37155_, _37139_);
  or (_37157_, _37156_, _06033_);
  and (_37158_, _37157_, _06027_);
  and (_37159_, _37158_, _37154_);
  or (_37161_, _37136_, _15074_);
  and (_37162_, _37161_, _06026_);
  and (_37163_, _37162_, _37139_);
  or (_37164_, _37163_, _09815_);
  or (_37165_, _37164_, _37159_);
  and (_37166_, _37165_, _37123_);
  or (_37167_, _37166_, _07011_);
  and (_37168_, _09179_, _07705_);
  or (_37169_, _37120_, _07012_);
  or (_37170_, _37169_, _37168_);
  and (_37172_, _37170_, _05669_);
  and (_37173_, _37172_, _37167_);
  and (_37174_, _15179_, _07705_);
  or (_37175_, _37174_, _37120_);
  and (_37176_, _37175_, _09833_);
  or (_37177_, _37176_, _06019_);
  or (_37178_, _37177_, _37173_);
  and (_37179_, _08652_, _07705_);
  or (_37180_, _37179_, _37120_);
  or (_37181_, _37180_, _06020_);
  and (_37183_, _37181_, _37178_);
  or (_37184_, _37183_, _06112_);
  and (_37185_, _15195_, _07705_);
  or (_37186_, _37185_, _37120_);
  or (_37187_, _37186_, _08751_);
  and (_37188_, _37187_, _08756_);
  and (_37189_, _37188_, _37184_);
  and (_37190_, _12306_, _07705_);
  or (_37191_, _37190_, _37120_);
  and (_37192_, _37191_, _06284_);
  or (_37194_, _37192_, _37189_);
  and (_37195_, _37194_, _07032_);
  or (_37196_, _37120_, _07980_);
  and (_37197_, _37180_, _06108_);
  and (_37198_, _37197_, _37196_);
  or (_37199_, _37198_, _37195_);
  and (_37200_, _37199_, _06278_);
  and (_37201_, _37129_, _06277_);
  and (_37202_, _37201_, _37196_);
  or (_37203_, _37202_, _06130_);
  or (_37205_, _37203_, _37200_);
  and (_37206_, _15194_, _07705_);
  or (_37207_, _37120_, _08777_);
  or (_37208_, _37207_, _37206_);
  and (_37209_, _37208_, _08782_);
  and (_37210_, _37209_, _37205_);
  nor (_37211_, _10982_, _13745_);
  or (_37212_, _37211_, _37120_);
  and (_37213_, _37212_, _06292_);
  or (_37214_, _37213_, _06316_);
  or (_37216_, _37214_, _37210_);
  or (_37217_, _37125_, _06718_);
  and (_37218_, _37217_, _05653_);
  and (_37219_, _37218_, _37216_);
  and (_37220_, _37151_, _05652_);
  or (_37221_, _37220_, _06047_);
  or (_37222_, _37221_, _37219_);
  and (_37223_, _15253_, _07705_);
  or (_37224_, _37120_, _06048_);
  or (_37225_, _37224_, _37223_);
  and (_37227_, _37225_, _01336_);
  and (_37228_, _37227_, _37222_);
  or (_37229_, _37228_, _37119_);
  and (_43515_, _37229_, _42882_);
  nor (_37230_, _01336_, _17846_);
  or (_37231_, _10871_, _10567_);
  and (_37232_, _37231_, _10824_);
  or (_37233_, _10796_, _10512_);
  or (_37234_, _37233_, _10811_);
  and (_37235_, _06229_, _05731_);
  and (_37237_, _06136_, _05731_);
  and (_37238_, _07005_, _05731_);
  or (_37239_, _10293_, _10237_);
  and (_37240_, _37239_, _37238_);
  and (_37241_, _15396_, _07705_);
  nor (_37242_, _07705_, _17846_);
  or (_37243_, _37242_, _08777_);
  or (_37244_, _37243_, _37241_);
  nor (_37245_, _07883_, _13745_);
  or (_37246_, _37245_, _37242_);
  or (_37248_, _37246_, _09827_);
  and (_37249_, _15293_, _07705_);
  or (_37250_, _37249_, _37242_);
  or (_37251_, _37250_, _06954_);
  and (_37252_, _07705_, \oc8051_golden_model_1.ACC [6]);
  or (_37253_, _37252_, _37242_);
  and (_37254_, _37253_, _06938_);
  nor (_37255_, _06938_, _17846_);
  or (_37256_, _37255_, _06102_);
  or (_37257_, _37256_, _37254_);
  and (_37259_, _37257_, _06044_);
  and (_37260_, _37259_, _37251_);
  nor (_37261_, _08355_, _17846_);
  and (_37262_, _15280_, _08355_);
  or (_37263_, _37262_, _37261_);
  and (_37264_, _37263_, _06043_);
  or (_37265_, _37264_, _06239_);
  or (_37266_, _37265_, _37260_);
  or (_37267_, _37246_, _06848_);
  and (_37268_, _37267_, _37266_);
  or (_37270_, _37268_, _06219_);
  or (_37271_, _37253_, _06220_);
  and (_37272_, _37271_, _06040_);
  and (_37273_, _37272_, _37270_);
  and (_37274_, _15278_, _08355_);
  or (_37275_, _37274_, _37261_);
  and (_37276_, _37275_, _06039_);
  or (_37277_, _37276_, _06032_);
  or (_37278_, _37277_, _37273_);
  or (_37279_, _37261_, _15310_);
  and (_37281_, _37279_, _37263_);
  or (_37282_, _37281_, _06033_);
  and (_37283_, _37282_, _10469_);
  and (_37284_, _37283_, _37278_);
  or (_37285_, _12361_, _10237_);
  or (_37286_, _37285_, _10483_);
  and (_37287_, _37286_, _12368_);
  or (_37288_, _37287_, _37284_);
  or (_37289_, _10512_, _13935_);
  or (_37290_, _37289_, _10549_);
  and (_37292_, _37290_, _37288_);
  or (_37293_, _37292_, _12367_);
  or (_37294_, _10311_, _06267_);
  or (_37295_, _37294_, _10360_);
  or (_37296_, _10567_, _10307_);
  or (_37297_, _37296_, _10621_);
  and (_37298_, _37297_, _06027_);
  and (_37299_, _37298_, _37295_);
  and (_37300_, _37299_, _37293_);
  or (_37301_, _37261_, _15326_);
  and (_37303_, _37301_, _06026_);
  and (_37304_, _37303_, _37263_);
  or (_37305_, _37304_, _09815_);
  or (_37306_, _37305_, _37300_);
  and (_37307_, _37306_, _37248_);
  or (_37308_, _37307_, _07011_);
  and (_37309_, _09178_, _07705_);
  or (_37310_, _37242_, _07012_);
  or (_37311_, _37310_, _37309_);
  and (_37312_, _37311_, _05669_);
  and (_37314_, _37312_, _37308_);
  and (_37315_, _15382_, _07705_);
  or (_37316_, _37315_, _37242_);
  and (_37317_, _37316_, _09833_);
  or (_37318_, _37317_, _06019_);
  or (_37319_, _37318_, _37314_);
  and (_37320_, _15389_, _07705_);
  or (_37321_, _37320_, _37242_);
  or (_37322_, _37321_, _06020_);
  and (_37323_, _37322_, _37319_);
  or (_37325_, _37323_, _06112_);
  and (_37326_, _15399_, _07705_);
  or (_37327_, _37326_, _37242_);
  or (_37328_, _37327_, _08751_);
  and (_37329_, _37328_, _08756_);
  and (_37330_, _37329_, _37325_);
  and (_37331_, _10980_, _07705_);
  or (_37332_, _37331_, _37242_);
  and (_37333_, _37332_, _06284_);
  or (_37334_, _37333_, _37330_);
  and (_37336_, _37334_, _07032_);
  or (_37337_, _37242_, _07886_);
  and (_37338_, _37321_, _06108_);
  and (_37339_, _37338_, _37337_);
  or (_37340_, _37339_, _37336_);
  and (_37341_, _37340_, _06278_);
  and (_37342_, _37253_, _06277_);
  and (_37343_, _37342_, _37337_);
  or (_37344_, _37343_, _06130_);
  or (_37345_, _37344_, _37341_);
  and (_37347_, _37345_, _37244_);
  or (_37348_, _37347_, _06292_);
  nor (_37349_, _10979_, _13745_);
  or (_37350_, _37349_, _37242_);
  nor (_37351_, _37350_, _08782_);
  nor (_37352_, _37351_, _37238_);
  and (_37353_, _37352_, _37348_);
  nor (_37354_, _37353_, _37240_);
  nor (_37355_, _37354_, _37237_);
  and (_37356_, _37239_, _37237_);
  nor (_37358_, _37356_, _37355_);
  nor (_37359_, _37358_, _37235_);
  and (_37360_, _06227_, _05731_);
  and (_37361_, _37239_, _37235_);
  or (_37362_, _37361_, _37360_);
  or (_37363_, _37362_, _37359_);
  and (_37364_, _07002_, _05731_);
  not (_37365_, _37360_);
  nor (_37366_, _37239_, _37365_);
  nor (_37367_, _37366_, _37364_);
  and (_37369_, _37367_, _37363_);
  and (_37370_, _37239_, _37364_);
  or (_37371_, _37370_, _10794_);
  or (_37372_, _37371_, _37369_);
  and (_37373_, _37372_, _37234_);
  or (_37374_, _37373_, _06288_);
  or (_37375_, _10311_, _06289_);
  or (_37376_, _37375_, _10841_);
  and (_37377_, _37376_, _10856_);
  and (_37378_, _37377_, _37374_);
  or (_37380_, _37378_, _37232_);
  and (_37381_, _37380_, _10890_);
  and (_37382_, _10920_, _16956_);
  or (_37383_, _37382_, _10932_);
  or (_37384_, _37383_, _37381_);
  or (_37385_, _10961_, _10934_);
  and (_37386_, _37385_, _06052_);
  and (_37387_, _37386_, _37384_);
  or (_37388_, _11002_, _10974_);
  and (_37389_, _37388_, _10976_);
  or (_37391_, _37389_, _37387_);
  or (_37392_, _11042_, _11050_);
  and (_37393_, _37392_, _37391_);
  or (_37394_, _37393_, _06316_);
  or (_37395_, _37250_, _06718_);
  and (_37396_, _37395_, _05653_);
  and (_37397_, _37396_, _37394_);
  and (_37398_, _37275_, _05652_);
  or (_37399_, _37398_, _06047_);
  or (_37400_, _37399_, _37397_);
  and (_37402_, _15451_, _07705_);
  or (_37403_, _37242_, _06048_);
  or (_37404_, _37403_, _37402_);
  and (_37405_, _37404_, _01336_);
  and (_37406_, _37405_, _37400_);
  or (_37407_, _37406_, _37230_);
  and (_43516_, _37407_, _42882_);
  and (_37408_, _05750_, op0_cnst);
  or (_00001_, _37408_, rst);
  and (_37409_, inst_finished_r, op0_cnst);
  nor (_37411_, word_in[3], word_in[2]);
  not (_37412_, _37411_);
  not (_37413_, word_in[1]);
  and (_37414_, _37413_, word_in[0]);
  and (_37415_, _37414_, \oc8051_golden_model_1.IRAM[1] [1]);
  nor (_37416_, _37413_, word_in[0]);
  and (_37417_, _37416_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor (_37418_, _37417_, _37415_);
  nor (_37419_, word_in[1], word_in[0]);
  and (_37420_, _37419_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_37422_, word_in[1], word_in[0]);
  and (_37423_, _37422_, \oc8051_golden_model_1.IRAM[3] [1]);
  nor (_37424_, _37423_, _37420_);
  and (_37425_, _37424_, _37418_);
  nor (_37426_, _37425_, _37412_);
  and (_37427_, word_in[3], word_in[2]);
  not (_37428_, _37427_);
  and (_37429_, _37414_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_37430_, _37416_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor (_37431_, _37430_, _37429_);
  and (_37433_, _37419_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_37434_, _37422_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor (_37435_, _37434_, _37433_);
  and (_37436_, _37435_, _37431_);
  nor (_37437_, _37436_, _37428_);
  nor (_37438_, _37437_, _37426_);
  not (_37439_, word_in[3]);
  and (_37440_, _37439_, word_in[2]);
  not (_37441_, _37440_);
  and (_37442_, _37414_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_37444_, _37416_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor (_37445_, _37444_, _37442_);
  and (_37446_, _37419_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_37447_, _37422_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor (_37448_, _37447_, _37446_);
  and (_37449_, _37448_, _37445_);
  nor (_37450_, _37449_, _37441_);
  nor (_37451_, _37439_, word_in[2]);
  not (_37452_, _37451_);
  and (_37453_, _37414_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_37455_, _37416_, \oc8051_golden_model_1.IRAM[10] [1]);
  nor (_37456_, _37455_, _37453_);
  and (_37457_, _37419_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_37458_, _37422_, \oc8051_golden_model_1.IRAM[11] [1]);
  nor (_37459_, _37458_, _37457_);
  and (_37460_, _37459_, _37456_);
  nor (_37461_, _37460_, _37452_);
  nor (_37462_, _37461_, _37450_);
  and (_37463_, _37462_, _37438_);
  and (_37464_, _37440_, _37422_);
  and (_37466_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_37467_, _37440_, _37416_);
  and (_37468_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_37469_, _37468_, _37466_);
  and (_37470_, _37427_, _37414_);
  and (_37471_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_37472_, _37427_, _37419_);
  and (_37473_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_37474_, _37473_, _37471_);
  and (_37475_, _37474_, _37469_);
  and (_37477_, _37416_, _37411_);
  and (_37478_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_37479_, _37414_, _37411_);
  and (_37480_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_37481_, _37480_, _37478_);
  and (_37482_, _37427_, _37416_);
  and (_37483_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_37484_, _37451_, _37419_);
  and (_37485_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_37486_, _37485_, _37483_);
  and (_37488_, _37486_, _37481_);
  and (_37489_, _37488_, _37475_);
  and (_37490_, _37451_, _37414_);
  and (_37491_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_37492_, _37419_, _37411_);
  and (_37493_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_37494_, _37493_, _37491_);
  and (_37495_, _37451_, _37416_);
  and (_37496_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_37497_, _37440_, _37414_);
  and (_37499_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_37500_, _37499_, _37496_);
  and (_37501_, _37500_, _37494_);
  and (_37502_, _37427_, _37422_);
  and (_37503_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_37504_, _37440_, _37419_);
  and (_37505_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_37506_, _37505_, _37503_);
  and (_37507_, _37451_, _37422_);
  and (_37508_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_37510_, _37422_, _37411_);
  and (_37511_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_37512_, _37511_, _37508_);
  and (_37513_, _37512_, _37506_);
  and (_37514_, _37513_, _37501_);
  and (_37515_, _37514_, _37489_);
  nand (_37516_, _37515_, _37463_);
  or (_37517_, _37515_, _37463_);
  and (_37518_, _37517_, _37516_);
  and (_37519_, _37414_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_37521_, _37416_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor (_37522_, _37521_, _37519_);
  and (_37523_, _37419_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_37524_, _37422_, \oc8051_golden_model_1.IRAM[3] [0]);
  nor (_37525_, _37524_, _37523_);
  and (_37526_, _37525_, _37522_);
  nor (_37527_, _37526_, _37412_);
  and (_37528_, _37414_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_37529_, _37416_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor (_37530_, _37529_, _37528_);
  and (_37532_, _37419_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_37533_, _37422_, \oc8051_golden_model_1.IRAM[11] [0]);
  nor (_37534_, _37533_, _37532_);
  and (_37535_, _37534_, _37530_);
  nor (_37536_, _37535_, _37452_);
  nor (_37537_, _37536_, _37527_);
  and (_37538_, _37414_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_37539_, _37416_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor (_37540_, _37539_, _37538_);
  and (_37541_, _37419_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_37543_, _37422_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor (_37544_, _37543_, _37541_);
  and (_37545_, _37544_, _37540_);
  nor (_37546_, _37545_, _37441_);
  and (_37547_, _37414_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_37548_, _37416_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor (_37549_, _37548_, _37547_);
  and (_37550_, _37419_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_37551_, _37422_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor (_37552_, _37551_, _37550_);
  and (_37554_, _37552_, _37549_);
  nor (_37555_, _37554_, _37428_);
  nor (_37556_, _37555_, _37546_);
  and (_37557_, _37556_, _37537_);
  and (_37558_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_37559_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_37560_, _37559_, _37558_);
  and (_37561_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_37562_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_37563_, _37562_, _37561_);
  and (_37565_, _37563_, _37560_);
  and (_37566_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_37567_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_37568_, _37567_, _37566_);
  and (_37569_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_37570_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_37571_, _37570_, _37569_);
  and (_37572_, _37571_, _37568_);
  and (_37573_, _37572_, _37565_);
  and (_37574_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_37576_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_37577_, _37576_, _37574_);
  and (_37578_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_37579_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_37580_, _37579_, _37578_);
  and (_37581_, _37580_, _37577_);
  and (_37582_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_37583_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_37584_, _37583_, _37582_);
  and (_37585_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_37587_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_37588_, _37587_, _37585_);
  and (_37589_, _37588_, _37584_);
  and (_37590_, _37589_, _37581_);
  and (_37591_, _37590_, _37573_);
  not (_37592_, _37591_);
  nor (_37593_, _37592_, _37557_);
  and (_37594_, _37592_, _37557_);
  or (_37595_, _37594_, _37593_);
  or (_37596_, _37595_, _37518_);
  and (_37598_, _37414_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_37599_, _37416_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor (_37600_, _37599_, _37598_);
  and (_37601_, _37419_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_37602_, _37422_, \oc8051_golden_model_1.IRAM[3] [3]);
  nor (_37603_, _37602_, _37601_);
  and (_37604_, _37603_, _37600_);
  nor (_37605_, _37604_, _37412_);
  and (_37606_, _37414_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_37607_, _37416_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor (_37609_, _37607_, _37606_);
  and (_37610_, _37419_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_37611_, _37422_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor (_37612_, _37611_, _37610_);
  and (_37613_, _37612_, _37609_);
  nor (_37614_, _37613_, _37428_);
  nor (_37615_, _37614_, _37605_);
  and (_37616_, _37414_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_37617_, _37416_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor (_37618_, _37617_, _37616_);
  and (_37620_, _37419_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_37621_, _37422_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor (_37622_, _37621_, _37620_);
  and (_37623_, _37622_, _37618_);
  nor (_37624_, _37623_, _37441_);
  and (_37625_, _37414_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_37626_, _37416_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor (_37627_, _37626_, _37625_);
  and (_37628_, _37419_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_37629_, _37422_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor (_37631_, _37629_, _37628_);
  and (_37632_, _37631_, _37627_);
  nor (_37633_, _37632_, _37452_);
  nor (_37634_, _37633_, _37624_);
  and (_37635_, _37634_, _37615_);
  and (_37636_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_37637_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_37638_, _37637_, _37636_);
  and (_37639_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_37640_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_37642_, _37640_, _37639_);
  and (_37643_, _37642_, _37638_);
  and (_37644_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_37645_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_37646_, _37645_, _37644_);
  and (_37647_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_37648_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_37649_, _37648_, _37647_);
  and (_37650_, _37649_, _37646_);
  and (_37651_, _37650_, _37643_);
  and (_37653_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_37654_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_37655_, _37654_, _37653_);
  and (_37656_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_37657_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_37658_, _37657_, _37656_);
  and (_37659_, _37658_, _37655_);
  and (_37660_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_37661_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_37662_, _37661_, _37660_);
  and (_37664_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_37665_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_37666_, _37665_, _37664_);
  and (_37667_, _37666_, _37662_);
  and (_37668_, _37667_, _37659_);
  and (_37669_, _37668_, _37651_);
  nand (_37670_, _37669_, _37635_);
  or (_37671_, _37669_, _37635_);
  and (_37672_, _37671_, _37670_);
  and (_37673_, _37414_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_37675_, _37416_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor (_37676_, _37675_, _37673_);
  and (_37677_, _37419_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_37678_, _37422_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor (_37679_, _37678_, _37677_);
  and (_37680_, _37679_, _37676_);
  nor (_37681_, _37680_, _37412_);
  and (_37682_, _37414_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_37683_, _37416_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor (_37684_, _37683_, _37682_);
  and (_37686_, _37419_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_37687_, _37422_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor (_37688_, _37687_, _37686_);
  and (_37689_, _37688_, _37684_);
  nor (_37690_, _37689_, _37452_);
  nor (_37691_, _37690_, _37681_);
  and (_37692_, _37414_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_37693_, _37416_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor (_37694_, _37693_, _37692_);
  and (_37695_, _37419_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_37697_, _37422_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor (_37698_, _37697_, _37695_);
  and (_37699_, _37698_, _37694_);
  nor (_37700_, _37699_, _37441_);
  and (_37701_, _37414_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_37702_, _37416_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor (_37703_, _37702_, _37701_);
  and (_37704_, _37419_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_37705_, _37422_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor (_37706_, _37705_, _37704_);
  and (_37708_, _37706_, _37703_);
  nor (_37709_, _37708_, _37428_);
  nor (_37710_, _37709_, _37700_);
  and (_37711_, _37710_, _37691_);
  and (_37712_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_37713_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_37714_, _37713_, _37712_);
  and (_37715_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_37716_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_37717_, _37716_, _37715_);
  and (_37719_, _37717_, _37714_);
  and (_37720_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_37721_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_37722_, _37721_, _37720_);
  and (_37723_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_37724_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_37725_, _37724_, _37723_);
  and (_37726_, _37725_, _37722_);
  and (_37727_, _37726_, _37719_);
  and (_37728_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_37730_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_37731_, _37730_, _37728_);
  and (_37732_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_37733_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_37734_, _37733_, _37732_);
  and (_37735_, _37734_, _37731_);
  and (_37736_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_37737_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_37738_, _37737_, _37736_);
  and (_37739_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and (_37741_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_37742_, _37741_, _37739_);
  and (_37743_, _37742_, _37738_);
  and (_37744_, _37743_, _37735_);
  and (_37745_, _37744_, _37727_);
  nand (_37746_, _37745_, _37711_);
  or (_37747_, _37745_, _37711_);
  and (_37748_, _37747_, _37746_);
  or (_37749_, _37748_, _37672_);
  or (_37750_, _37749_, _37596_);
  and (_37752_, _37414_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_37753_, _37416_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor (_37754_, _37753_, _37752_);
  and (_37755_, _37419_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_37756_, _37422_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor (_37757_, _37756_, _37755_);
  and (_37758_, _37757_, _37754_);
  nor (_37759_, _37758_, _37441_);
  and (_37760_, _37414_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_37761_, _37416_, \oc8051_golden_model_1.IRAM[10] [4]);
  nor (_37763_, _37761_, _37760_);
  and (_37764_, _37419_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_37765_, _37422_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor (_37766_, _37765_, _37764_);
  and (_37767_, _37766_, _37763_);
  nor (_37768_, _37767_, _37452_);
  nor (_37769_, _37768_, _37759_);
  and (_37770_, _37414_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_37771_, _37416_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor (_37772_, _37771_, _37770_);
  and (_37774_, _37419_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_37775_, _37422_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor (_37776_, _37775_, _37774_);
  and (_37777_, _37776_, _37772_);
  nor (_37778_, _37777_, _37412_);
  and (_37779_, _37414_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_37780_, _37416_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor (_37781_, _37780_, _37779_);
  and (_37782_, _37419_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_37783_, _37422_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor (_37785_, _37783_, _37782_);
  and (_37786_, _37785_, _37781_);
  nor (_37787_, _37786_, _37428_);
  nor (_37788_, _37787_, _37778_);
  and (_37789_, _37788_, _37769_);
  not (_37790_, _37789_);
  and (_37791_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_37792_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_37793_, _37792_, _37791_);
  and (_37794_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_37796_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_37797_, _37796_, _37794_);
  and (_37798_, _37797_, _37793_);
  and (_37799_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_37800_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_37801_, _37800_, _37799_);
  and (_37802_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_37803_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_37804_, _37803_, _37802_);
  and (_37805_, _37804_, _37801_);
  and (_37807_, _37805_, _37798_);
  and (_37808_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_37809_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_37810_, _37809_, _37808_);
  and (_37811_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_37812_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_37813_, _37812_, _37811_);
  and (_37814_, _37813_, _37810_);
  and (_37815_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_37816_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_37818_, _37816_, _37815_);
  and (_37819_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_37820_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_37821_, _37820_, _37819_);
  and (_37822_, _37821_, _37818_);
  and (_37823_, _37822_, _37814_);
  and (_37824_, _37823_, _37807_);
  nor (_37825_, _37824_, _37790_);
  and (_37826_, _37824_, _37790_);
  or (_37827_, _37826_, _37825_);
  and (_37829_, _37414_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_37830_, _37416_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor (_37831_, _37830_, _37829_);
  and (_37832_, _37419_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_37833_, _37422_, \oc8051_golden_model_1.IRAM[3] [5]);
  nor (_37834_, _37833_, _37832_);
  and (_37835_, _37834_, _37831_);
  nor (_37836_, _37835_, _37412_);
  and (_37837_, _37414_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_37838_, _37416_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor (_37840_, _37838_, _37837_);
  and (_37841_, _37419_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_37842_, _37422_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor (_37843_, _37842_, _37841_);
  and (_37844_, _37843_, _37840_);
  nor (_37845_, _37844_, _37428_);
  nor (_37846_, _37845_, _37836_);
  and (_37847_, _37414_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_37848_, _37416_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor (_37849_, _37848_, _37847_);
  and (_37851_, _37419_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_37852_, _37422_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor (_37853_, _37852_, _37851_);
  and (_37854_, _37853_, _37849_);
  nor (_37855_, _37854_, _37441_);
  and (_37856_, _37414_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_37857_, _37416_, \oc8051_golden_model_1.IRAM[10] [5]);
  nor (_37858_, _37857_, _37856_);
  and (_37859_, _37419_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_37860_, _37422_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor (_37862_, _37860_, _37859_);
  and (_37863_, _37862_, _37858_);
  nor (_37864_, _37863_, _37452_);
  nor (_37865_, _37864_, _37855_);
  and (_37866_, _37865_, _37846_);
  and (_37867_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_37868_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_37869_, _37868_, _37867_);
  and (_37870_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_37871_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_37873_, _37871_, _37870_);
  and (_37874_, _37873_, _37869_);
  and (_37875_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_37876_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_37877_, _37876_, _37875_);
  and (_37878_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_37879_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_37880_, _37879_, _37878_);
  and (_37881_, _37880_, _37877_);
  and (_37882_, _37881_, _37874_);
  and (_37884_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_37885_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_37886_, _37885_, _37884_);
  and (_37887_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_37888_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_37889_, _37888_, _37887_);
  and (_37890_, _37889_, _37886_);
  and (_37891_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_37892_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_37893_, _37892_, _37891_);
  and (_37895_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_37896_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_37897_, _37896_, _37895_);
  and (_37898_, _37897_, _37893_);
  and (_37899_, _37898_, _37890_);
  and (_37900_, _37899_, _37882_);
  nand (_37901_, _37900_, _37866_);
  or (_37902_, _37900_, _37866_);
  and (_37903_, _37902_, _37901_);
  or (_37904_, _37903_, _37827_);
  and (_37906_, _37414_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_37907_, _37416_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor (_37908_, _37907_, _37906_);
  and (_37909_, _37419_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_37910_, _37422_, \oc8051_golden_model_1.IRAM[3] [6]);
  nor (_37911_, _37910_, _37909_);
  and (_37912_, _37911_, _37908_);
  nor (_37913_, _37912_, _37412_);
  and (_37914_, _37414_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_37915_, _37416_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor (_37917_, _37915_, _37914_);
  and (_37918_, _37419_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_37919_, _37422_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor (_37920_, _37919_, _37918_);
  and (_37921_, _37920_, _37917_);
  nor (_37922_, _37921_, _37452_);
  nor (_37923_, _37922_, _37913_);
  and (_37924_, _37414_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_37925_, _37416_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor (_37926_, _37925_, _37924_);
  and (_37928_, _37419_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_37929_, _37422_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor (_37930_, _37929_, _37928_);
  and (_37931_, _37930_, _37926_);
  nor (_37932_, _37931_, _37441_);
  and (_37933_, _37414_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_37934_, _37416_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor (_37935_, _37934_, _37933_);
  and (_37936_, _37419_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_37937_, _37422_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor (_37939_, _37937_, _37936_);
  and (_37940_, _37939_, _37935_);
  nor (_37941_, _37940_, _37428_);
  nor (_37942_, _37941_, _37932_);
  and (_37943_, _37942_, _37923_);
  and (_37944_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_37945_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_37946_, _37945_, _37944_);
  and (_37947_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_37948_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_37950_, _37948_, _37947_);
  and (_37951_, _37950_, _37946_);
  and (_37952_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_37953_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_37954_, _37953_, _37952_);
  and (_37955_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_37956_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_37957_, _37956_, _37955_);
  and (_37958_, _37957_, _37954_);
  and (_37959_, _37958_, _37951_);
  and (_37961_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_37962_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_37963_, _37962_, _37961_);
  and (_37964_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_37965_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_37966_, _37965_, _37964_);
  and (_37967_, _37966_, _37963_);
  and (_37968_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_37969_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_37970_, _37969_, _37968_);
  and (_37972_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_37973_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_37974_, _37973_, _37972_);
  and (_37975_, _37974_, _37970_);
  and (_37976_, _37975_, _37967_);
  and (_37977_, _37976_, _37959_);
  nand (_37978_, _37977_, _37943_);
  or (_37979_, _37977_, _37943_);
  and (_37980_, _37979_, _37978_);
  and (_37981_, _37414_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_37983_, _37416_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor (_37984_, _37983_, _37981_);
  and (_37985_, _37419_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_37986_, _37422_, \oc8051_golden_model_1.IRAM[7] [7]);
  nor (_37987_, _37986_, _37985_);
  and (_37988_, _37987_, _37984_);
  nor (_37989_, _37988_, _37441_);
  and (_37990_, _37414_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_37991_, _37416_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_37992_, _37991_, _37990_);
  and (_37994_, _37419_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_37995_, _37422_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor (_37996_, _37995_, _37994_);
  and (_37997_, _37996_, _37992_);
  nor (_37998_, _37997_, _37428_);
  nor (_37999_, _37998_, _37989_);
  and (_38000_, _37414_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_38001_, _37416_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor (_38002_, _38001_, _38000_);
  and (_38003_, _37419_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_38005_, _37422_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor (_38006_, _38005_, _38003_);
  and (_38007_, _38006_, _38002_);
  nor (_38008_, _38007_, _37412_);
  and (_38009_, _37414_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_38010_, _37416_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor (_38011_, _38010_, _38009_);
  and (_38012_, _37419_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_38013_, _37422_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor (_38014_, _38013_, _38012_);
  and (_38016_, _38014_, _38011_);
  nor (_38017_, _38016_, _37452_);
  nor (_38018_, _38017_, _38008_);
  and (_38019_, _38018_, _37999_);
  and (_38020_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_38021_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_38022_, _38021_, _38020_);
  and (_38023_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_38024_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_38025_, _38024_, _38023_);
  and (_38027_, _38025_, _38022_);
  and (_38028_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_38029_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_38030_, _38029_, _38028_);
  and (_38031_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_38032_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_38033_, _38032_, _38031_);
  and (_38034_, _38033_, _38030_);
  and (_38035_, _38034_, _38027_);
  and (_38036_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_38038_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_38039_, _38038_, _38036_);
  and (_38040_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_38041_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_38042_, _38041_, _38040_);
  and (_38043_, _38042_, _38039_);
  and (_38044_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_38045_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_38046_, _38045_, _38044_);
  and (_38047_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_38049_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_38050_, _38049_, _38047_);
  and (_38051_, _38050_, _38046_);
  and (_38052_, _38051_, _38043_);
  and (_38053_, _38052_, _38035_);
  nand (_38054_, _38053_, _38019_);
  or (_38055_, _38053_, _38019_);
  and (_38056_, _38055_, _38054_);
  or (_38057_, _38056_, _37980_);
  or (_38058_, _38057_, _37904_);
  or (_38060_, _38058_, _37750_);
  and (property_invalid_iram, _38060_, _37409_);
  nor (_38061_, _09956_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_38062_, _09956_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_38063_, _38062_, _38061_);
  nand (_38064_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_38065_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38066_, _38065_, _38064_);
  or (_38067_, _38066_, _38063_);
  and (_38068_, _05784_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_38070_, _05784_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_38071_, _38070_, _38068_);
  and (_38072_, _05758_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_38073_, \oc8051_golden_model_1.ACC [0], _39048_);
  or (_38074_, _38073_, _38072_);
  or (_38075_, _38074_, _38071_);
  or (_38076_, _38075_, _38067_);
  or (_38077_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_38078_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_38079_, _38078_, _38077_);
  or (_38081_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_38082_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38083_, _38082_, _38081_);
  or (_38084_, _38083_, _38079_);
  nand (_38085_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_38086_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_38087_, _38086_, _38085_);
  and (_38088_, _08393_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_38089_, _08393_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_38090_, _38089_, _38088_);
  or (_38092_, _38090_, _38087_);
  or (_38093_, _38092_, _38084_);
  or (_38094_, _38093_, _38076_);
  and (property_invalid_acc, _38094_, _37409_);
  and (_38095_, _37408_, _01336_);
  nor (_38096_, _25378_, _01937_);
  and (_38097_, _25378_, _01937_);
  or (_38098_, _38097_, _38096_);
  nor (_38099_, _25728_, _01941_);
  nor (_38100_, _26416_, _01949_);
  or (_38102_, _38100_, _38099_);
  nor (_38103_, _26769_, _01953_);
  and (_38104_, _26416_, _01949_);
  or (_38105_, _38104_, _38103_);
  or (_38106_, _38105_, _38102_);
  nor (_38107_, _26067_, _01945_);
  and (_38108_, _28118_, _38558_);
  nor (_38109_, _28118_, _38558_);
  and (_38110_, _12796_, _38536_);
  nor (_38111_, _12796_, _38536_);
  or (_38113_, _38111_, _38110_);
  and (_38114_, _27796_, _38552_);
  nor (_38115_, _29339_, _38544_);
  or (_38116_, _38115_, _38114_);
  or (_38117_, _38116_, _38113_);
  nand (_38118_, _25007_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_38119_, _25007_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_38120_, _38119_, _38118_);
  nor (_38121_, _29649_, _38540_);
  or (_38122_, _38121_, _38120_);
  nor (_38124_, _28728_, _38548_);
  and (_38125_, _28728_, _38548_);
  and (_38126_, _29649_, _38540_);
  or (_38127_, _38126_, _38125_);
  or (_38128_, _38127_, _38124_);
  or (_38129_, _38128_, _38122_);
  nor (_38130_, _27796_, _38552_);
  and (_38131_, _29339_, _38544_);
  or (_38132_, _38131_, _38130_);
  or (_38133_, _38132_, _38129_);
  or (_38135_, _38133_, _38117_);
  and (_38136_, _28426_, _38563_);
  nor (_38137_, _28426_, _38563_);
  or (_38138_, _38137_, _38136_);
  and (_38139_, _29035_, _38569_);
  nor (_38140_, _29035_, _38569_);
  or (_38141_, _38140_, _38139_);
  or (_38142_, _38141_, _38138_);
  or (_38143_, _38142_, _38135_);
  or (_38144_, _38143_, _38109_);
  or (_38146_, _38144_, _38108_);
  or (_38147_, _38146_, _38107_);
  nor (_38148_, _27474_, _01960_);
  and (_38149_, _27474_, _01960_);
  or (_38150_, _38149_, _38148_);
  and (_38151_, _26067_, _01945_);
  nand (_38152_, _27119_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_38153_, _27119_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_38154_, _38153_, _38152_);
  or (_38155_, _38154_, _38151_);
  or (_38157_, _38155_, _38150_);
  or (_38158_, _38157_, _38147_);
  and (_38159_, _25728_, _01941_);
  and (_38160_, _26769_, _01953_);
  or (_38161_, _38160_, _38159_);
  or (_38162_, _38161_, _38158_);
  or (_38163_, _38162_, _38106_);
  or (_38164_, _38163_, _38098_);
  and (property_invalid_pc, _38164_, _38095_);
  buf (_00543_, _42885_);
  buf (_05103_, _42882_);
  buf (_05155_, _42882_);
  buf (_05206_, _42882_);
  buf (_05258_, _42882_);
  buf (_05309_, _42882_);
  buf (_05362_, _42882_);
  buf (_05415_, _42882_);
  buf (_05468_, _42882_);
  buf (_05521_, _42882_);
  buf (_05574_, _42882_);
  buf (_05627_, _42882_);
  buf (_05680_, _42882_);
  buf (_05733_, _42882_);
  buf (_05786_, _42882_);
  buf (_05839_, _42882_);
  buf (_05892_, _42882_);
  buf (_39058_, _38956_);
  buf (_39060_, _38958_);
  buf (_39073_, _38956_);
  buf (_39074_, _38958_);
  buf (_39386_, _38975_);
  buf (_39387_, _38976_);
  buf (_39388_, _38978_);
  buf (_39389_, _38979_);
  buf (_39390_, _38980_);
  buf (_39391_, _38981_);
  buf (_39392_, _38982_);
  buf (_39393_, _38984_);
  buf (_39394_, _38985_);
  buf (_39396_, _38986_);
  buf (_39397_, _38987_);
  buf (_39398_, _38988_);
  buf (_39399_, _38990_);
  buf (_39400_, _38991_);
  buf (_39451_, _38975_);
  buf (_39452_, _38976_);
  buf (_39453_, _38978_);
  buf (_39454_, _38979_);
  buf (_39455_, _38980_);
  buf (_39456_, _38981_);
  buf (_39457_, _38982_);
  buf (_39458_, _38984_);
  buf (_39459_, _38985_);
  buf (_39461_, _38986_);
  buf (_39462_, _38987_);
  buf (_39463_, _38988_);
  buf (_39464_, _38990_);
  buf (_39465_, _38991_);
  buf (_39855_, _39760_);
  buf (_40018_, _39760_);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _05107_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _05111_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _05115_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _05119_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _05123_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _05126_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _05130_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _05100_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _05103_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _05159_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _05162_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _05166_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _05170_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _05174_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _05178_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _05182_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _05152_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _05155_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _05631_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _05635_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _05639_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _05643_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _05647_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _05651_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _05655_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _05624_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _05627_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _05684_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _05688_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _05692_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _05696_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _05700_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _05704_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _05708_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _05677_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _05680_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _05737_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _05741_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _05745_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _05749_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _05753_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _05757_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _05761_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _05730_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _05733_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _05790_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _05794_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _05798_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _05802_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _05806_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _05810_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _05814_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _05783_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _05786_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _05843_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _05847_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _05851_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _05855_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _05859_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _05863_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _05867_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _05836_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _05839_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _05896_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _05900_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _05904_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _05908_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _05912_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _05916_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _05920_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _05889_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _05892_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _05210_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _05214_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _05218_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _05222_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _05226_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _05230_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _05234_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _05203_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _05206_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _05262_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _05266_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _05270_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _05273_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _05277_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _05281_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _05285_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _05255_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _05258_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _05313_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _05317_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _05321_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _05325_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _05329_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _05333_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _05337_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _05306_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _05309_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _05366_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _05370_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _05374_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _05378_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _05382_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _05386_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _05390_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _05359_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _05362_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _05419_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _05423_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _05427_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _05431_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _05435_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _05439_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _05443_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _05412_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _05415_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _05472_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _05476_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _05480_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _05484_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _05488_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _05492_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _05496_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _05465_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _05468_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _05525_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _05529_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _05533_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _05537_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _05541_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _05545_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _05549_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _05518_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _05521_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _05578_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _05582_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _05586_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _05590_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _05594_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _05598_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _05602_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _05571_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _05574_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _40967_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _40968_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _40969_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _40970_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _40971_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _40972_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _40973_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _40751_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _40956_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _40957_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _40958_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _40959_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _40960_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _40962_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _40963_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _40964_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _40943_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _40945_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _40946_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _40947_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _40948_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _40949_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _40951_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _40952_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _40932_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _40933_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _40934_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _40935_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _40936_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _40937_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _40939_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _40940_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _40919_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _40920_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _40921_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _40924_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _40925_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _40926_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _40927_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _40928_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _40908_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _40909_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _40910_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _40912_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _40913_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _40914_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _40915_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _40916_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _40896_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _40897_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _40898_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _40899_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _40901_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _40902_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _40903_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _40904_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _40884_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _40885_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _40886_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _40887_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _40889_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _40890_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _40891_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _40892_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _40872_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _40873_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _40874_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _40876_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _40877_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _40878_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _40879_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _40880_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _40860_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _40861_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _40862_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _40863_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _40864_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _40865_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _40866_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _40867_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _40848_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _40849_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _40850_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _40851_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _40853_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _40854_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _40855_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _40856_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _40835_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _40836_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _40837_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _40838_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _40841_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _40842_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _40843_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _40844_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _40823_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _40824_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _40825_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _40827_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _40828_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _40829_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _40830_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _40831_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _40813_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _40814_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _40815_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _40816_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _40818_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _40819_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _40820_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _40821_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _40801_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _40802_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _40803_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _40805_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _40806_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _40807_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _40808_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _40809_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _40792_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _40793_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _40794_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _40795_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _40797_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _40798_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _40799_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _40800_);
  dff (\oc8051_golden_model_1.B [0], _43324_);
  dff (\oc8051_golden_model_1.B [1], _43325_);
  dff (\oc8051_golden_model_1.B [2], _43326_);
  dff (\oc8051_golden_model_1.B [3], _43327_);
  dff (\oc8051_golden_model_1.B [4], _43328_);
  dff (\oc8051_golden_model_1.B [5], _43329_);
  dff (\oc8051_golden_model_1.B [6], _43330_);
  dff (\oc8051_golden_model_1.B [7], _40752_);
  dff (\oc8051_golden_model_1.ACC [0], _43332_);
  dff (\oc8051_golden_model_1.ACC [1], _43333_);
  dff (\oc8051_golden_model_1.ACC [2], _43334_);
  dff (\oc8051_golden_model_1.ACC [3], _43335_);
  dff (\oc8051_golden_model_1.ACC [4], _43336_);
  dff (\oc8051_golden_model_1.ACC [5], _43338_);
  dff (\oc8051_golden_model_1.ACC [6], _43339_);
  dff (\oc8051_golden_model_1.ACC [7], _40753_);
  dff (\oc8051_golden_model_1.PCON [0], _43340_);
  dff (\oc8051_golden_model_1.PCON [1], _43342_);
  dff (\oc8051_golden_model_1.PCON [2], _43343_);
  dff (\oc8051_golden_model_1.PCON [3], _43344_);
  dff (\oc8051_golden_model_1.PCON [4], _43345_);
  dff (\oc8051_golden_model_1.PCON [5], _43346_);
  dff (\oc8051_golden_model_1.PCON [6], _43347_);
  dff (\oc8051_golden_model_1.PCON [7], _40756_);
  dff (\oc8051_golden_model_1.TMOD [0], _43349_);
  dff (\oc8051_golden_model_1.TMOD [1], _43350_);
  dff (\oc8051_golden_model_1.TMOD [2], _43351_);
  dff (\oc8051_golden_model_1.TMOD [3], _43352_);
  dff (\oc8051_golden_model_1.TMOD [4], _43353_);
  dff (\oc8051_golden_model_1.TMOD [5], _43354_);
  dff (\oc8051_golden_model_1.TMOD [6], _43355_);
  dff (\oc8051_golden_model_1.TMOD [7], _40757_);
  dff (\oc8051_golden_model_1.DPL [0], _43357_);
  dff (\oc8051_golden_model_1.DPL [1], _43358_);
  dff (\oc8051_golden_model_1.DPL [2], _43359_);
  dff (\oc8051_golden_model_1.DPL [3], _43361_);
  dff (\oc8051_golden_model_1.DPL [4], _43362_);
  dff (\oc8051_golden_model_1.DPL [5], _43363_);
  dff (\oc8051_golden_model_1.DPL [6], _43364_);
  dff (\oc8051_golden_model_1.DPL [7], _40758_);
  dff (\oc8051_golden_model_1.DPH [0], _43366_);
  dff (\oc8051_golden_model_1.DPH [1], _43367_);
  dff (\oc8051_golden_model_1.DPH [2], _43368_);
  dff (\oc8051_golden_model_1.DPH [3], _43369_);
  dff (\oc8051_golden_model_1.DPH [4], _43370_);
  dff (\oc8051_golden_model_1.DPH [5], _43371_);
  dff (\oc8051_golden_model_1.DPH [6], _43372_);
  dff (\oc8051_golden_model_1.DPH [7], _40759_);
  dff (\oc8051_golden_model_1.TL1 [0], _43374_);
  dff (\oc8051_golden_model_1.TL1 [1], _43375_);
  dff (\oc8051_golden_model_1.TL1 [2], _43376_);
  dff (\oc8051_golden_model_1.TL1 [3], _43377_);
  dff (\oc8051_golden_model_1.TL1 [4], _43378_);
  dff (\oc8051_golden_model_1.TL1 [5], _43380_);
  dff (\oc8051_golden_model_1.TL1 [6], _43381_);
  dff (\oc8051_golden_model_1.TL1 [7], _40760_);
  dff (\oc8051_golden_model_1.TL0 [0], _43382_);
  dff (\oc8051_golden_model_1.TL0 [1], _43384_);
  dff (\oc8051_golden_model_1.TL0 [2], _43385_);
  dff (\oc8051_golden_model_1.TL0 [3], _43386_);
  dff (\oc8051_golden_model_1.TL0 [4], _43387_);
  dff (\oc8051_golden_model_1.TL0 [5], _43388_);
  dff (\oc8051_golden_model_1.TL0 [6], _43389_);
  dff (\oc8051_golden_model_1.TL0 [7], _40762_);
  dff (\oc8051_golden_model_1.TCON [0], _43391_);
  dff (\oc8051_golden_model_1.TCON [1], _43392_);
  dff (\oc8051_golden_model_1.TCON [2], _43393_);
  dff (\oc8051_golden_model_1.TCON [3], _43394_);
  dff (\oc8051_golden_model_1.TCON [4], _43395_);
  dff (\oc8051_golden_model_1.TCON [5], _43396_);
  dff (\oc8051_golden_model_1.TCON [6], _43397_);
  dff (\oc8051_golden_model_1.TCON [7], _40763_);
  dff (\oc8051_golden_model_1.TH1 [0], _43399_);
  dff (\oc8051_golden_model_1.TH1 [1], _43400_);
  dff (\oc8051_golden_model_1.TH1 [2], _43401_);
  dff (\oc8051_golden_model_1.TH1 [3], _43403_);
  dff (\oc8051_golden_model_1.TH1 [4], _43404_);
  dff (\oc8051_golden_model_1.TH1 [5], _43405_);
  dff (\oc8051_golden_model_1.TH1 [6], _43406_);
  dff (\oc8051_golden_model_1.TH1 [7], _40764_);
  dff (\oc8051_golden_model_1.TH0 [0], _43408_);
  dff (\oc8051_golden_model_1.TH0 [1], _43409_);
  dff (\oc8051_golden_model_1.TH0 [2], _43410_);
  dff (\oc8051_golden_model_1.TH0 [3], _43411_);
  dff (\oc8051_golden_model_1.TH0 [4], _43412_);
  dff (\oc8051_golden_model_1.TH0 [5], _43413_);
  dff (\oc8051_golden_model_1.TH0 [6], _43414_);
  dff (\oc8051_golden_model_1.TH0 [7], _40765_);
  dff (\oc8051_golden_model_1.PC [0], _43417_);
  dff (\oc8051_golden_model_1.PC [1], _43418_);
  dff (\oc8051_golden_model_1.PC [2], _43419_);
  dff (\oc8051_golden_model_1.PC [3], _43420_);
  dff (\oc8051_golden_model_1.PC [4], _43421_);
  dff (\oc8051_golden_model_1.PC [5], _43422_);
  dff (\oc8051_golden_model_1.PC [6], _43423_);
  dff (\oc8051_golden_model_1.PC [7], _43425_);
  dff (\oc8051_golden_model_1.PC [8], _43426_);
  dff (\oc8051_golden_model_1.PC [9], _43427_);
  dff (\oc8051_golden_model_1.PC [10], _43428_);
  dff (\oc8051_golden_model_1.PC [11], _43429_);
  dff (\oc8051_golden_model_1.PC [12], _43430_);
  dff (\oc8051_golden_model_1.PC [13], _43431_);
  dff (\oc8051_golden_model_1.PC [14], _43432_);
  dff (\oc8051_golden_model_1.PC [15], _40766_);
  dff (\oc8051_golden_model_1.P2 [0], _43434_);
  dff (\oc8051_golden_model_1.P2 [1], _43435_);
  dff (\oc8051_golden_model_1.P2 [2], _43436_);
  dff (\oc8051_golden_model_1.P2 [3], _43437_);
  dff (\oc8051_golden_model_1.P2 [4], _43438_);
  dff (\oc8051_golden_model_1.P2 [5], _43440_);
  dff (\oc8051_golden_model_1.P2 [6], _43441_);
  dff (\oc8051_golden_model_1.P2 [7], _40768_);
  dff (\oc8051_golden_model_1.P3 [0], _43442_);
  dff (\oc8051_golden_model_1.P3 [1], _43444_);
  dff (\oc8051_golden_model_1.P3 [2], _43445_);
  dff (\oc8051_golden_model_1.P3 [3], _43446_);
  dff (\oc8051_golden_model_1.P3 [4], _43447_);
  dff (\oc8051_golden_model_1.P3 [5], _43448_);
  dff (\oc8051_golden_model_1.P3 [6], _43449_);
  dff (\oc8051_golden_model_1.P3 [7], _40769_);
  dff (\oc8051_golden_model_1.P0 [0], _43451_);
  dff (\oc8051_golden_model_1.P0 [1], _43452_);
  dff (\oc8051_golden_model_1.P0 [2], _43453_);
  dff (\oc8051_golden_model_1.P0 [3], _43454_);
  dff (\oc8051_golden_model_1.P0 [4], _43455_);
  dff (\oc8051_golden_model_1.P0 [5], _43456_);
  dff (\oc8051_golden_model_1.P0 [6], _43457_);
  dff (\oc8051_golden_model_1.P0 [7], _40770_);
  dff (\oc8051_golden_model_1.P1 [0], _43459_);
  dff (\oc8051_golden_model_1.P1 [1], _43460_);
  dff (\oc8051_golden_model_1.P1 [2], _43461_);
  dff (\oc8051_golden_model_1.P1 [3], _43463_);
  dff (\oc8051_golden_model_1.P1 [4], _43464_);
  dff (\oc8051_golden_model_1.P1 [5], _43465_);
  dff (\oc8051_golden_model_1.P1 [6], _43466_);
  dff (\oc8051_golden_model_1.P1 [7], _40771_);
  dff (\oc8051_golden_model_1.IP [0], _43468_);
  dff (\oc8051_golden_model_1.IP [1], _43469_);
  dff (\oc8051_golden_model_1.IP [2], _43470_);
  dff (\oc8051_golden_model_1.IP [3], _43471_);
  dff (\oc8051_golden_model_1.IP [4], _43472_);
  dff (\oc8051_golden_model_1.IP [5], _43473_);
  dff (\oc8051_golden_model_1.IP [6], _43474_);
  dff (\oc8051_golden_model_1.IP [7], _40772_);
  dff (\oc8051_golden_model_1.IE [0], _43476_);
  dff (\oc8051_golden_model_1.IE [1], _43477_);
  dff (\oc8051_golden_model_1.IE [2], _43478_);
  dff (\oc8051_golden_model_1.IE [3], _43479_);
  dff (\oc8051_golden_model_1.IE [4], _43480_);
  dff (\oc8051_golden_model_1.IE [5], _43482_);
  dff (\oc8051_golden_model_1.IE [6], _43483_);
  dff (\oc8051_golden_model_1.IE [7], _40774_);
  dff (\oc8051_golden_model_1.SCON [0], _43484_);
  dff (\oc8051_golden_model_1.SCON [1], _43486_);
  dff (\oc8051_golden_model_1.SCON [2], _43487_);
  dff (\oc8051_golden_model_1.SCON [3], _43488_);
  dff (\oc8051_golden_model_1.SCON [4], _43489_);
  dff (\oc8051_golden_model_1.SCON [5], _43490_);
  dff (\oc8051_golden_model_1.SCON [6], _43491_);
  dff (\oc8051_golden_model_1.SCON [7], _40775_);
  dff (\oc8051_golden_model_1.SP [0], _43493_);
  dff (\oc8051_golden_model_1.SP [1], _43494_);
  dff (\oc8051_golden_model_1.SP [2], _43495_);
  dff (\oc8051_golden_model_1.SP [3], _43496_);
  dff (\oc8051_golden_model_1.SP [4], _43497_);
  dff (\oc8051_golden_model_1.SP [5], _43498_);
  dff (\oc8051_golden_model_1.SP [6], _43499_);
  dff (\oc8051_golden_model_1.SP [7], _40776_);
  dff (\oc8051_golden_model_1.SBUF [0], _43501_);
  dff (\oc8051_golden_model_1.SBUF [1], _43502_);
  dff (\oc8051_golden_model_1.SBUF [2], _43503_);
  dff (\oc8051_golden_model_1.SBUF [3], _43505_);
  dff (\oc8051_golden_model_1.SBUF [4], _43506_);
  dff (\oc8051_golden_model_1.SBUF [5], _43507_);
  dff (\oc8051_golden_model_1.SBUF [6], _43508_);
  dff (\oc8051_golden_model_1.SBUF [7], _40777_);
  dff (\oc8051_golden_model_1.PSW [0], _43510_);
  dff (\oc8051_golden_model_1.PSW [1], _43511_);
  dff (\oc8051_golden_model_1.PSW [2], _43512_);
  dff (\oc8051_golden_model_1.PSW [3], _43513_);
  dff (\oc8051_golden_model_1.PSW [4], _43514_);
  dff (\oc8051_golden_model_1.PSW [5], _43515_);
  dff (\oc8051_golden_model_1.PSW [6], _43516_);
  dff (\oc8051_golden_model_1.PSW [7], _40778_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02832_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02844_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02866_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02890_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02914_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00956_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _02924_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00925_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _02936_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _02948_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _02960_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _02971_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _02984_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _02997_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03011_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00976_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02356_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22216_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02542_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02695_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _02877_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03117_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03361_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03562_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03757_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _03954_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04054_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04147_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04246_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04345_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04444_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04542_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04641_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24374_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38968_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38969_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38970_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38971_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38972_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38973_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38974_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38955_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38975_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38976_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38978_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38979_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38980_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38981_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38982_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38956_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38984_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38985_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38986_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38987_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38988_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38990_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38991_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38958_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _34275_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _34278_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _09716_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _34280_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _34282_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _09719_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _34284_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _09722_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _34286_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _34288_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _34290_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _09725_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _34292_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _09728_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _09731_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09790_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09792_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _09695_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09795_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09798_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _09698_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _09801_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _09701_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _09804_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _09807_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _09810_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _09813_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _09816_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _09819_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _09822_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _09704_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _09707_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _34273_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _09713_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _09825_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _09710_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39760_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _39792_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _39793_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _39794_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _39795_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _39796_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _39797_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _39798_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _39762_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _39799_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _39800_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _39801_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _39803_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _39804_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _39805_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _39806_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _39763_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _39807_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _39808_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _39809_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _39810_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _39811_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _39812_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _39814_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _39764_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _39815_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _39816_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _39817_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _39818_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _39819_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _39820_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _39821_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _39765_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39339_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39340_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39341_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39342_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _39056_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _39128_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _39129_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _39130_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _39131_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _39132_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _39134_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _39135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _39136_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _39137_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _39138_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _39139_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _39140_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _39141_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39142_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39143_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _39015_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39148_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39149_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39150_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39151_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39152_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39153_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39154_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39155_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39156_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39157_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39159_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39160_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39161_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39162_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39163_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _39016_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39343_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39344_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39345_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39346_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39348_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39349_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39350_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39351_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39352_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39353_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39354_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39355_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39356_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39357_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39359_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39360_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39361_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39362_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39363_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39364_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39365_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39366_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39367_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39368_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39370_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39371_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39372_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39373_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39374_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39375_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39376_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _39081_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _39054_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39377_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39379_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39380_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39381_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39382_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39383_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39385_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _39057_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39386_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39387_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39388_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39389_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39390_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39391_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39392_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _39058_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39393_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39394_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39396_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39397_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39398_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39399_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39400_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _39060_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _39061_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _39062_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39401_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39402_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39403_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39404_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39405_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39407_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39408_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _39063_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39409_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39410_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39411_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39412_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39413_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39414_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39415_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39416_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39418_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39419_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39420_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39421_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39422_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39423_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39424_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _39064_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39425_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39426_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39427_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39429_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39430_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39431_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39432_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39433_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39434_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39435_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39436_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39437_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39438_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39440_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39441_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _39066_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _39067_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _39069_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _39068_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39442_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39443_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39444_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39445_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39446_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39447_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39448_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _39071_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39449_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39450_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _39072_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39451_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39452_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39453_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39454_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39455_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39456_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39457_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _39073_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39458_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39459_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39461_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39462_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39463_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39464_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39465_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _39074_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _39075_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39466_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39467_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39468_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39469_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39470_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39472_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39473_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _39076_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _39078_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _39079_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39474_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39475_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39476_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _39080_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39477_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39478_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39479_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39480_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39481_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39483_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39484_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39485_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39486_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39487_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39488_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39489_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39490_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39491_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39492_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39494_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39495_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39496_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39497_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39498_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39499_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39500_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39501_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39502_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39503_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39505_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39506_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39507_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39508_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39509_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39510_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _39082_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39511_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39512_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39513_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39514_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39516_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39517_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39518_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _39083_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _39084_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _39086_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39519_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39520_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39521_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39522_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39523_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39524_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39525_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39527_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39528_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39529_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39530_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39531_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39532_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39533_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39534_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _39087_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _39088_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _39089_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _39090_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39535_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39536_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39538_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39539_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39540_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39541_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39542_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39543_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39544_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39545_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39546_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39547_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39549_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39550_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39551_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _39091_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _39092_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _40015_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _40036_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _40037_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _40039_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _40040_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _40041_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _40042_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _40043_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _40016_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _40018_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _40044_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _40045_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _40019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _02796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _02801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _02806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _02811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _02815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _02820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _02825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _02827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _02835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _02838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _02841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _02845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _02849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _02852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _02855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _02858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _02864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _02868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _02871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _02875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _02878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _02882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _02885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _02888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _02926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _02929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _02933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _02937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _02940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _02943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _02947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _02950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _02894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _02898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _02902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _02905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _02909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _02912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _02916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _02919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _02983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _02987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _02991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _02994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _02999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _02954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _02957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _02962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _02965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _02968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _02972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _02976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _02978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _02573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _05083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _05084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _05086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _05090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _05092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02563_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _39849_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _39935_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _39936_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _39937_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _39850_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _39851_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _39853_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39938_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39939_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39940_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39941_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39943_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39944_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39945_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39854_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39855_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19849_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19860_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19872_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19884_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19896_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19908_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19920_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _17998_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08903_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08914_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08925_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08936_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08947_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08958_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08969_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06662_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13668_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13679_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13712_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12713_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13723_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13733_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13744_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13755_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13766_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13777_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13788_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12734_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _42886_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _42885_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _42882_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42880_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _42879_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _42877_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _42875_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _42873_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42872_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42870_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _42840_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _42838_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _42836_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _42834_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _42832_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00171_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _42830_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00176_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00178_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00182_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00185_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _42827_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _40589_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _40591_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _40593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _40595_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _40597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _40599_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _40601_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _31126_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _40603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _40605_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _40607_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _40609_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _40611_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _40612_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _40614_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _31149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _40616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _40618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _40620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _40622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _40624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _40626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _40628_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _31172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _40630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _40632_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _40634_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _40636_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _40638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _40640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _40642_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _31194_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17374_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17385_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17396_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17407_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17418_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17429_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15193_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09519_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10696_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10707_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10718_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10729_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10751_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09540_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _41092_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _41095_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _41601_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _41603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _41605_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _41606_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _41608_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _41610_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _41612_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _41098_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _41614_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _41616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _41618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _41620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _41622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _41623_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _41625_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _41101_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _41104_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _41107_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _41627_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _41629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _41631_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _41633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _41635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _41637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _41638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _41110_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _41640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _41642_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _41644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _41646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _41648_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _41650_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _41652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _41113_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _41116_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _41653_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _41655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _41657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _41659_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _41660_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _41662_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _41664_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _41119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01628_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01631_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01634_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02108_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02109_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02113_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02116_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02118_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02120_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02122_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02123_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02125_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02127_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02129_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02137_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02144_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02146_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02148_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02157_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01658_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01210_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01212_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01214_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01216_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01218_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01220_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01222_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01224_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01226_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01228_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01229_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00567_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00543_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00546_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00548_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00551_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00554_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00556_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01231_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00559_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01233_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01235_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01237_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00562_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01241_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01243_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01249_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01251_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00564_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00570_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00572_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00578_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01253_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01255_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01257_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00583_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01259_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01261_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01263_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01264_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01268_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01270_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01272_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01274_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01276_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00586_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01278_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01280_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01282_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01284_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01286_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01288_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01290_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00588_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01292_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01299_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01301_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01303_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00591_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [0], \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [1], \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [2], \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [3], \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [4], \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [5], \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [6], \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [7], \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [0], \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [1], \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [2], \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [3], \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [4], \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [5], \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [6], \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [7], \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [0], \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [1], \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [2], \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [3], \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [4], \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [5], \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [6], \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [7], \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [0], \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [1], \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [2], \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [3], \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [4], \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [5], \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [6], \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [7], \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0994 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0994 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0994 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0994 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0994 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0994 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0994 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1071 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1071 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1071 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1071 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1073 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1075 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1075 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1076 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1076 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1077 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1077 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1078 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1078 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1079 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1079 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1080 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1080 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1081 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1118 , \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.n1146 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1147 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1147 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1147 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1147 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1147 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1147 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1148 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1148 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1148 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1148 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1148 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1148 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1148 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1149 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1149 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1149 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1149 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1149 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1149 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1149 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1149 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1150 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1151 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1152 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1152 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1152 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1153 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1154 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1154 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1155 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1155 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1155 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1155 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1155 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1155 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1181 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1181 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1181 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1181 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1181 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1181 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1181 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1181 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1181 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1181 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1181 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1181 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1181 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1181 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1181 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1181 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1183 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1183 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1183 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1183 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1183 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1183 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1183 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1183 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1185 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1185 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1185 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1185 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1185 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1185 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1185 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1189 [8], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1190 , \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1191 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1191 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1191 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1191 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1192 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1192 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1192 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1196 [4], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1197 , \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1198 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1198 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1198 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1198 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1198 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1198 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1198 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1198 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1198 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1206 , \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.n1207 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1207 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1207 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1207 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1207 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1211 [8], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1212 , \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1217 [4], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1218 , \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1226 , \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.n1227 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1227 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1227 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1227 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1227 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1229 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1229 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1229 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1229 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1229 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1229 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1229 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1229 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1229 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1231 [8], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1232 , \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1233 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1233 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1233 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1233 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1234 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1234 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1234 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1236 [4], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1237 , \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1238 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1238 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1238 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1238 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1238 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1238 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1238 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1238 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1238 [8], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1245 , \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1246 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1246 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1246 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1246 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1249 [8], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1257 , \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.n1258 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1258 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1258 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1258 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1258 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1260 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1262 [8], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1264 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1267 , \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1268 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1276 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1276 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1276 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1276 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1276 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1276 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1278 [4], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1279 , \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1280 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1280 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1280 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1280 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1280 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1280 [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1282 [8], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1283 , \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1290 , \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1291 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1291 [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1291 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1291 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1291 [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1292 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1292 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1292 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1292 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1292 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1295 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1295 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1295 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1295 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1295 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1295 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1295 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1295 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1295 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1296 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1296 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1296 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1296 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1296 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1296 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1296 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1297 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1297 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1297 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1297 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1297 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1297 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1297 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1297 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1298 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1299 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1299 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1299 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1299 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1299 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1299 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1299 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1299 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1300 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1300 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1303 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1305 [8], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1306 , \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1307 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1307 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1309 [4], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1310 , \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1317 , \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.n1318 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1318 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1318 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1318 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1318 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1322 [8], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1323 , \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1333 , \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.n1334 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1334 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1334 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1334 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1334 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1338 [8], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1339 , \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1342 , \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1350 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1350 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1354 [8], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1355 , \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1357 [4], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1358 , \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1365 , \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.n1366 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1366 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1366 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1366 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1366 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1520 , \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1521 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1521 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1521 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1521 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1521 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1521 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1521 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1553 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1553 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1553 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1553 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.n1555 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1555 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1555 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1555 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1555 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1555 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1555 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1680 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1683 , \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.n1685 , \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.n1691 , \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.n1692 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1692 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1692 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1692 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1692 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1696 , \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.n1698 , \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1709 , \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.n1711 , \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.n1717 , \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.n1718 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1718 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1718 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1718 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1718 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1722 , \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.n1724 , \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.n1730 , \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.n1731 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1731 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1731 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1731 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1731 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1733 , \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.n1734 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1734 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1734 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1734 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1734 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1734 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1734 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1735 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1735 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1735 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1735 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1735 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1735 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1735 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1739 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n1739 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n1739 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n1739 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n1739 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n1739 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n1739 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n1739 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n1739 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [9], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [10], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [11], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [12], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [13], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [14], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1745 , \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.n1746 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1746 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1746 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1746 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1746 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1746 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1746 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1749 , \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.n1750 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1750 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1750 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1750 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1750 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1750 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1750 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1765 , \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.n1766 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1766 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1766 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1766 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1766 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1766 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1766 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1771 , \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.n1772 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1772 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1772 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1772 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1772 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1772 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1772 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1777 , \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.n1778 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1778 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1778 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1778 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1778 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1778 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1778 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1783 , \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.n1784 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1784 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1784 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1784 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1784 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1784 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1784 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1789 , \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.n1790 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1790 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1790 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1790 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1790 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1790 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1790 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1791 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1791 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1791 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1791 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1791 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1791 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1792 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1792 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1792 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1792 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1793 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1793 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1793 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1793 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1793 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1793 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1828 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1828 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1828 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1828 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1828 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1828 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1828 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1828 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1847 , \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.n1848 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1848 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1848 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1848 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1848 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1848 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1848 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1852 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1852 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1852 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1852 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [0], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1853 [1], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1853 [2], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1853 [3], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1854 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1854 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1854 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1854 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
