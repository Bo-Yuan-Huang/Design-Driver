
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pc, property_invalid_acc, property_invalid_iram);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire _44007_;
  wire _44008_;
  wire _44009_;
  wire _44010_;
  wire _44011_;
  wire _44012_;
  wire _44013_;
  wire _44014_;
  wire _44015_;
  wire _44016_;
  wire _44017_;
  wire _44018_;
  wire _44019_;
  wire _44020_;
  wire _44021_;
  wire _44022_;
  wire _44023_;
  wire _44024_;
  wire _44025_;
  wire _44026_;
  wire _44027_;
  wire _44028_;
  wire [7:0] ACC_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [7:0] \oc8051_golden_model_1.n0994 ;
  wire [3:0] \oc8051_golden_model_1.n1090 ;
  wire [3:0] \oc8051_golden_model_1.n1092 ;
  wire [3:0] \oc8051_golden_model_1.n1094 ;
  wire [3:0] \oc8051_golden_model_1.n1095 ;
  wire [3:0] \oc8051_golden_model_1.n1096 ;
  wire [3:0] \oc8051_golden_model_1.n1097 ;
  wire [3:0] \oc8051_golden_model_1.n1098 ;
  wire [3:0] \oc8051_golden_model_1.n1099 ;
  wire [3:0] \oc8051_golden_model_1.n1100 ;
  wire \oc8051_golden_model_1.n1147 ;
  wire \oc8051_golden_model_1.n1175 ;
  wire [8:0] \oc8051_golden_model_1.n1176 ;
  wire [8:0] \oc8051_golden_model_1.n1177 ;
  wire [7:0] \oc8051_golden_model_1.n1178 ;
  wire \oc8051_golden_model_1.n1179 ;
  wire \oc8051_golden_model_1.n1180 ;
  wire [2:0] \oc8051_golden_model_1.n1181 ;
  wire \oc8051_golden_model_1.n1182 ;
  wire [1:0] \oc8051_golden_model_1.n1183 ;
  wire [7:0] \oc8051_golden_model_1.n1184 ;
  wire [15:0] \oc8051_golden_model_1.n1211 ;
  wire [7:0] \oc8051_golden_model_1.n1213 ;
  wire [8:0] \oc8051_golden_model_1.n1215 ;
  wire [8:0] \oc8051_golden_model_1.n1219 ;
  wire \oc8051_golden_model_1.n1220 ;
  wire [3:0] \oc8051_golden_model_1.n1221 ;
  wire [4:0] \oc8051_golden_model_1.n1222 ;
  wire [4:0] \oc8051_golden_model_1.n1226 ;
  wire \oc8051_golden_model_1.n1227 ;
  wire [8:0] \oc8051_golden_model_1.n1228 ;
  wire \oc8051_golden_model_1.n1236 ;
  wire [7:0] \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1241 ;
  wire \oc8051_golden_model_1.n1242 ;
  wire [4:0] \oc8051_golden_model_1.n1247 ;
  wire \oc8051_golden_model_1.n1248 ;
  wire \oc8051_golden_model_1.n1256 ;
  wire [7:0] \oc8051_golden_model_1.n1257 ;
  wire [8:0] \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1261 ;
  wire \oc8051_golden_model_1.n1262 ;
  wire [3:0] \oc8051_golden_model_1.n1263 ;
  wire [4:0] \oc8051_golden_model_1.n1264 ;
  wire [4:0] \oc8051_golden_model_1.n1266 ;
  wire \oc8051_golden_model_1.n1267 ;
  wire [8:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire [7:0] \oc8051_golden_model_1.n1276 ;
  wire [8:0] \oc8051_golden_model_1.n1279 ;
  wire \oc8051_golden_model_1.n1280 ;
  wire \oc8051_golden_model_1.n1287 ;
  wire [7:0] \oc8051_golden_model_1.n1288 ;
  wire [8:0] \oc8051_golden_model_1.n1290 ;
  wire [8:0] \oc8051_golden_model_1.n1292 ;
  wire \oc8051_golden_model_1.n1293 ;
  wire [4:0] \oc8051_golden_model_1.n1294 ;
  wire [4:0] \oc8051_golden_model_1.n1296 ;
  wire \oc8051_golden_model_1.n1297 ;
  wire [8:0] \oc8051_golden_model_1.n1298 ;
  wire \oc8051_golden_model_1.n1305 ;
  wire [7:0] \oc8051_golden_model_1.n1306 ;
  wire [4:0] \oc8051_golden_model_1.n1308 ;
  wire \oc8051_golden_model_1.n1309 ;
  wire [7:0] \oc8051_golden_model_1.n1310 ;
  wire [8:0] \oc8051_golden_model_1.n1312 ;
  wire \oc8051_golden_model_1.n1313 ;
  wire \oc8051_golden_model_1.n1320 ;
  wire [7:0] \oc8051_golden_model_1.n1321 ;
  wire [7:0] \oc8051_golden_model_1.n1322 ;
  wire [8:0] \oc8051_golden_model_1.n1325 ;
  wire [8:0] \oc8051_golden_model_1.n1326 ;
  wire [7:0] \oc8051_golden_model_1.n1327 ;
  wire \oc8051_golden_model_1.n1328 ;
  wire [7:0] \oc8051_golden_model_1.n1329 ;
  wire [7:0] \oc8051_golden_model_1.n1330 ;
  wire [8:0] \oc8051_golden_model_1.n1333 ;
  wire [8:0] \oc8051_golden_model_1.n1335 ;
  wire \oc8051_golden_model_1.n1336 ;
  wire [4:0] \oc8051_golden_model_1.n1337 ;
  wire [4:0] \oc8051_golden_model_1.n1339 ;
  wire \oc8051_golden_model_1.n1340 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire [7:0] \oc8051_golden_model_1.n1348 ;
  wire [8:0] \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire [4:0] \oc8051_golden_model_1.n1355 ;
  wire \oc8051_golden_model_1.n1356 ;
  wire \oc8051_golden_model_1.n1363 ;
  wire [7:0] \oc8051_golden_model_1.n1364 ;
  wire [8:0] \oc8051_golden_model_1.n1368 ;
  wire \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1371 ;
  wire \oc8051_golden_model_1.n1372 ;
  wire \oc8051_golden_model_1.n1379 ;
  wire [7:0] \oc8051_golden_model_1.n1380 ;
  wire [8:0] \oc8051_golden_model_1.n1384 ;
  wire \oc8051_golden_model_1.n1385 ;
  wire [4:0] \oc8051_golden_model_1.n1387 ;
  wire \oc8051_golden_model_1.n1388 ;
  wire \oc8051_golden_model_1.n1395 ;
  wire [7:0] \oc8051_golden_model_1.n1396 ;
  wire \oc8051_golden_model_1.n1556 ;
  wire [6:0] \oc8051_golden_model_1.n1557 ;
  wire [7:0] \oc8051_golden_model_1.n1558 ;
  wire \oc8051_golden_model_1.n1581 ;
  wire [7:0] \oc8051_golden_model_1.n1582 ;
  wire [3:0] \oc8051_golden_model_1.n1589 ;
  wire \oc8051_golden_model_1.n1590 ;
  wire [7:0] \oc8051_golden_model_1.n1591 ;
  wire [7:0] \oc8051_golden_model_1.n1735 ;
  wire \oc8051_golden_model_1.n1738 ;
  wire \oc8051_golden_model_1.n1740 ;
  wire \oc8051_golden_model_1.n1746 ;
  wire [7:0] \oc8051_golden_model_1.n1747 ;
  wire \oc8051_golden_model_1.n1751 ;
  wire \oc8051_golden_model_1.n1753 ;
  wire \oc8051_golden_model_1.n1759 ;
  wire [7:0] \oc8051_golden_model_1.n1760 ;
  wire \oc8051_golden_model_1.n1764 ;
  wire \oc8051_golden_model_1.n1766 ;
  wire \oc8051_golden_model_1.n1772 ;
  wire [7:0] \oc8051_golden_model_1.n1773 ;
  wire \oc8051_golden_model_1.n1777 ;
  wire \oc8051_golden_model_1.n1779 ;
  wire \oc8051_golden_model_1.n1785 ;
  wire [7:0] \oc8051_golden_model_1.n1786 ;
  wire \oc8051_golden_model_1.n1788 ;
  wire [7:0] \oc8051_golden_model_1.n1789 ;
  wire [7:0] \oc8051_golden_model_1.n1790 ;
  wire [15:0] \oc8051_golden_model_1.n1794 ;
  wire \oc8051_golden_model_1.n1800 ;
  wire [7:0] \oc8051_golden_model_1.n1801 ;
  wire \oc8051_golden_model_1.n1804 ;
  wire [7:0] \oc8051_golden_model_1.n1805 ;
  wire \oc8051_golden_model_1.n1825 ;
  wire [7:0] \oc8051_golden_model_1.n1826 ;
  wire \oc8051_golden_model_1.n1831 ;
  wire [7:0] \oc8051_golden_model_1.n1832 ;
  wire \oc8051_golden_model_1.n1837 ;
  wire [7:0] \oc8051_golden_model_1.n1838 ;
  wire \oc8051_golden_model_1.n1843 ;
  wire [7:0] \oc8051_golden_model_1.n1844 ;
  wire \oc8051_golden_model_1.n1849 ;
  wire [7:0] \oc8051_golden_model_1.n1850 ;
  wire [7:0] \oc8051_golden_model_1.n1851 ;
  wire [3:0] \oc8051_golden_model_1.n1852 ;
  wire [7:0] \oc8051_golden_model_1.n1853 ;
  wire [7:0] \oc8051_golden_model_1.n1889 ;
  wire \oc8051_golden_model_1.n1908 ;
  wire [7:0] \oc8051_golden_model_1.n1909 ;
  wire [7:0] \oc8051_golden_model_1.n1913 ;
  wire [3:0] \oc8051_golden_model_1.n1914 ;
  wire [7:0] \oc8051_golden_model_1.n1915 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff0 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff1 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff2 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff3 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_iram;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_43100_, rst);
  not (_18190_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_18201_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_18212_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _18201_);
  and (_18223_, _18212_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_18234_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _18201_);
  and (_18245_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _18201_);
  nor (_18256_, _18245_, _18234_);
  and (_18267_, _18256_, _18223_);
  nor (_18278_, _18267_, _18190_);
  and (_18289_, _18190_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18300_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_18311_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _18300_);
  nor (_18322_, _18311_, _18289_);
  not (_18333_, _18322_);
  and (_18344_, _18333_, _18267_);
  or (_18355_, _18344_, _18278_);
  and (_22218_, _18355_, _43100_);
  nor (_18376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18387_, _18376_);
  and (_18398_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_18409_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_18420_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_18431_, _18420_);
  not (_18442_, _18311_);
  nor (_18453_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_18464_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_18475_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _18464_);
  nor (_18486_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_18497_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_18507_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _18497_);
  nor (_18518_, _18507_, _18486_);
  nor (_18529_, _18518_, _18475_);
  not (_18540_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_18551_, _18475_, _18540_);
  nor (_18562_, _18551_, _18529_);
  and (_18573_, _18562_, _18453_);
  not (_18584_, _18573_);
  and (_18595_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_18606_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_18617_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_18628_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _18617_);
  and (_18639_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_18650_, _18639_, _18606_);
  and (_18671_, _18650_, _18584_);
  nor (_18672_, _18671_, _18442_);
  not (_18683_, _18289_);
  nor (_18704_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_18705_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _18497_);
  nor (_18716_, _18705_, _18704_);
  nor (_18737_, _18716_, _18475_);
  not (_18738_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_18749_, _18475_, _18738_);
  nor (_18770_, _18749_, _18737_);
  and (_18771_, _18770_, _18453_);
  not (_18782_, _18771_);
  and (_18803_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_18804_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_18815_, _18804_, _18803_);
  and (_18836_, _18815_, _18782_);
  nor (_18837_, _18836_, _18683_);
  nor (_18848_, _18837_, _18672_);
  nor (_18868_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_18869_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _18497_);
  nor (_18880_, _18869_, _18868_);
  nor (_18891_, _18880_, _18475_);
  not (_18902_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_18913_, _18475_, _18902_);
  nor (_18924_, _18913_, _18891_);
  and (_18935_, _18924_, _18453_);
  not (_18946_, _18935_);
  and (_18957_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_18968_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_18979_, _18968_, _18957_);
  and (_18990_, _18979_, _18946_);
  nor (_19001_, _18990_, _18333_);
  nor (_19012_, _19001_, _18376_);
  and (_19023_, _19012_, _18848_);
  nor (_19034_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_19045_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _18497_);
  nor (_19056_, _19045_, _19034_);
  nor (_19067_, _19056_, _18475_);
  not (_19078_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_19089_, _18475_, _19078_);
  nor (_19100_, _19089_, _19067_);
  and (_19111_, _19100_, _18453_);
  not (_19122_, _19111_);
  and (_19133_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_19144_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_19155_, _19144_, _19133_);
  and (_19166_, _19155_, _19122_);
  and (_19177_, _19166_, _18376_);
  nor (_19188_, _19177_, _19023_);
  not (_19199_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19210_, _19199_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19220_, _19210_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19231_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_19242_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19253_, _19242_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19264_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_19275_, _19264_, _19231_);
  nor (_19286_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19296_, _19286_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19307_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_19318_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19329_, _19210_, _19318_);
  and (_19340_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_19351_, _19340_, _19307_);
  and (_19362_, _19351_, _19275_);
  and (_19373_, _19286_, _19199_);
  and (_19383_, _19373_, _19100_);
  and (_19394_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19405_, _19394_, _19318_);
  and (_19416_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_19427_, _19394_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19438_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_19449_, _19438_, _19416_);
  not (_19460_, _19449_);
  nor (_19470_, _19460_, _19383_);
  and (_19481_, _19470_, _19362_);
  not (_19492_, _19481_);
  and (_19503_, _19492_, _19188_);
  not (_19514_, _19503_);
  nor (_19525_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_19536_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _18497_);
  nor (_19547_, _19536_, _19525_);
  nor (_19557_, _19547_, _18475_);
  not (_19568_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_19579_, _18475_, _19568_);
  nor (_19590_, _19579_, _19557_);
  and (_19601_, _19590_, _18453_);
  not (_19612_, _19601_);
  and (_19623_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_19634_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_19644_, _19634_, _19623_);
  and (_19655_, _19644_, _19612_);
  nor (_19666_, _19655_, _18442_);
  nor (_19677_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_19688_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _18497_);
  nor (_19699_, _19688_, _19677_);
  nor (_19710_, _19699_, _18475_);
  not (_19720_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_19731_, _18475_, _19720_);
  nor (_19742_, _19731_, _19710_);
  and (_19753_, _19742_, _18453_);
  not (_19764_, _19753_);
  and (_19775_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_19786_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_19797_, _19786_, _19775_);
  and (_19807_, _19797_, _19764_);
  nor (_19818_, _19807_, _18683_);
  nor (_19829_, _19818_, _19666_);
  nor (_19840_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_19862_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _18497_);
  nor (_19874_, _19862_, _19840_);
  nor (_19885_, _19874_, _18475_);
  not (_19897_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_19909_, _18475_, _19897_);
  nor (_19921_, _19909_, _19885_);
  and (_19933_, _19921_, _18453_);
  not (_19934_, _19933_);
  and (_19945_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_19956_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_19967_, _19956_, _19945_);
  and (_19977_, _19967_, _19934_);
  nor (_19988_, _19977_, _18333_);
  nor (_19999_, _19988_, _18376_);
  and (_20010_, _19999_, _19829_);
  nor (_20021_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_20032_, _18497_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_20043_, _20032_, _20021_);
  nor (_20054_, _20043_, _18475_);
  not (_20064_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_20075_, _18475_, _20064_);
  nor (_20086_, _20075_, _20054_);
  and (_20097_, _20086_, _18453_);
  not (_20108_, _20097_);
  and (_20119_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_20130_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_20141_, _20130_, _20119_);
  and (_20151_, _20141_, _20108_);
  and (_20162_, _20151_, _18376_);
  nor (_20173_, _20162_, _20010_);
  and (_20184_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_20195_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_20206_, _20195_, _20184_);
  and (_20217_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_20227_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_20238_, _20227_, _20217_);
  and (_20249_, _20238_, _20206_);
  and (_20260_, _20086_, _19373_);
  and (_20271_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_20282_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_20293_, _20282_, _20271_);
  not (_20304_, _20293_);
  nor (_20314_, _20304_, _20260_);
  and (_20325_, _20314_, _20249_);
  not (_20336_, _20325_);
  and (_20347_, _20336_, _20173_);
  and (_20358_, _20347_, _19514_);
  not (_20369_, _20358_);
  and (_20380_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_20391_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_20401_, _20391_, _20380_);
  and (_20412_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_20423_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_20434_, _20423_, _20412_);
  and (_20445_, _20434_, _20401_);
  and (_20456_, _19742_, _19373_);
  and (_20467_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_20478_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_20488_, _20478_, _20467_);
  not (_20499_, _20488_);
  nor (_20510_, _20499_, _20456_);
  and (_20521_, _20510_, _20445_);
  not (_20532_, _20521_);
  and (_20543_, _20532_, _20173_);
  and (_20554_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_20565_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_20575_, _20565_, _20554_);
  and (_20586_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_20597_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_20608_, _20597_, _20586_);
  and (_20619_, _20608_, _20575_);
  and (_20630_, _19373_, _18770_);
  and (_20641_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_20652_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_20663_, _20652_, _20641_);
  not (_20673_, _20663_);
  nor (_20684_, _20673_, _20630_);
  and (_20695_, _20684_, _20619_);
  not (_20706_, _20695_);
  and (_20717_, _20706_, _19188_);
  and (_20728_, _20543_, _20717_);
  and (_20739_, _19492_, _20728_);
  nor (_20750_, _19503_, _20728_);
  nor (_20770_, _20750_, _20739_);
  and (_20781_, _20770_, _20543_);
  and (_20782_, _20347_, _19503_);
  and (_20793_, _19492_, _20173_);
  and (_20814_, _20336_, _19188_);
  nor (_20825_, _20814_, _20793_);
  nor (_20826_, _20825_, _20782_);
  and (_20847_, _20826_, _20781_);
  nor (_20857_, _20826_, _20781_);
  nor (_20858_, _20857_, _20847_);
  and (_20869_, _20858_, _20739_);
  nor (_20880_, _20869_, _20847_);
  nor (_20891_, _20880_, _20369_);
  and (_20912_, _20173_, _20706_);
  and (_20913_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_20924_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_20935_, _20924_, _20913_);
  and (_20945_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_20956_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_20967_, _20956_, _20945_);
  and (_20978_, _20967_, _20935_);
  and (_20989_, _19590_, _19373_);
  and (_21000_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_21011_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_21022_, _21011_, _21000_);
  not (_21042_, _21022_);
  nor (_21043_, _21042_, _20989_);
  and (_21054_, _21043_, _20978_);
  not (_21065_, _21054_);
  and (_21076_, _21065_, _19188_);
  and (_21087_, _21076_, _20912_);
  and (_21098_, _20532_, _19188_);
  nor (_21109_, _21098_, _20912_);
  nor (_21120_, _21109_, _20728_);
  and (_21130_, _21120_, _21087_);
  nor (_21141_, _19503_, _20543_);
  nor (_21152_, _21141_, _20781_);
  and (_21163_, _21152_, _21130_);
  nor (_21174_, _20858_, _20739_);
  nor (_21185_, _21174_, _20869_);
  and (_21196_, _21185_, _21163_);
  nor (_21216_, _21185_, _21163_);
  nor (_21217_, _21216_, _21196_);
  not (_21228_, _21217_);
  and (_21239_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_21250_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_21261_, _21250_, _21239_);
  and (_21272_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_21283_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_21294_, _21283_, _21272_);
  and (_21305_, _21294_, _21261_);
  and (_21315_, _19921_, _19373_);
  and (_21326_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_21337_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_21348_, _21337_, _21326_);
  not (_21359_, _21348_);
  nor (_21370_, _21359_, _21315_);
  and (_21381_, _21370_, _21305_);
  not (_21392_, _21381_);
  and (_21412_, _21392_, _20173_);
  and (_21413_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_21424_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_21435_, _21424_, _21413_);
  and (_21446_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_21457_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_21468_, _21457_, _21446_);
  and (_21479_, _21468_, _21435_);
  and (_21490_, _19373_, _18562_);
  and (_21500_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_21511_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_21522_, _21511_, _21500_);
  not (_21533_, _21522_);
  nor (_21544_, _21533_, _21490_);
  and (_21555_, _21544_, _21479_);
  not (_21566_, _21555_);
  and (_21577_, _21566_, _19188_);
  and (_21588_, _21577_, _21412_);
  and (_21598_, _21392_, _19188_);
  not (_21609_, _21598_);
  and (_21620_, _21566_, _20173_);
  and (_21631_, _21620_, _21609_);
  and (_21642_, _21631_, _21076_);
  nor (_21653_, _21642_, _21588_);
  and (_21664_, _21065_, _20173_);
  nor (_21675_, _21664_, _20717_);
  nor (_21685_, _21675_, _21087_);
  not (_21696_, _21685_);
  nor (_21707_, _21696_, _21653_);
  nor (_21718_, _21120_, _21087_);
  nor (_21729_, _21718_, _21130_);
  and (_21740_, _21729_, _21707_);
  nor (_21760_, _21152_, _21130_);
  nor (_21761_, _21760_, _21163_);
  and (_21772_, _21761_, _21740_);
  and (_21783_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_21794_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_21805_, _21794_, _21783_);
  and (_21816_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_21827_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_21838_, _21827_, _21816_);
  and (_21848_, _21838_, _21805_);
  and (_21869_, _19373_, _18924_);
  and (_21870_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_21881_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_21892_, _21881_, _21870_);
  not (_21903_, _21892_);
  nor (_21914_, _21903_, _21869_);
  and (_21925_, _21914_, _21848_);
  not (_21935_, _21925_);
  and (_21946_, _21935_, _20173_);
  and (_21957_, _21946_, _21598_);
  nor (_21968_, _21577_, _21412_);
  nor (_21979_, _21968_, _21588_);
  and (_21990_, _21979_, _21957_);
  nor (_22001_, _21631_, _21076_);
  nor (_22012_, _22001_, _21642_);
  and (_22022_, _22012_, _21990_);
  and (_22033_, _21696_, _21653_);
  nor (_22044_, _22033_, _21707_);
  and (_22055_, _22044_, _22022_);
  nor (_22066_, _21729_, _21707_);
  nor (_22077_, _22066_, _21740_);
  and (_22088_, _22077_, _22055_);
  nor (_22098_, _21761_, _21740_);
  nor (_22109_, _22098_, _21772_);
  and (_22120_, _22109_, _22088_);
  nor (_22131_, _22120_, _21772_);
  nor (_22142_, _22131_, _21228_);
  nor (_22153_, _22142_, _21196_);
  and (_22164_, _20880_, _20369_);
  nor (_22175_, _22164_, _20891_);
  not (_22185_, _22175_);
  nor (_22196_, _22185_, _22153_);
  or (_22207_, _22196_, _20782_);
  nor (_22219_, _22207_, _20891_);
  nor (_22230_, _22219_, _18431_);
  and (_22241_, _22219_, _18431_);
  nor (_22252_, _22241_, _22230_);
  not (_22263_, _22252_);
  and (_22273_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_22284_, _22185_, _22153_);
  nor (_22295_, _22284_, _22196_);
  and (_22316_, _22295_, _22273_);
  and (_22317_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_22328_, _22131_, _21228_);
  nor (_22339_, _22328_, _22142_);
  and (_22349_, _22339_, _22317_);
  nor (_22360_, _22339_, _22317_);
  nor (_22371_, _22360_, _22349_);
  not (_22382_, _22371_);
  and (_22393_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_22404_, _22109_, _22088_);
  nor (_22415_, _22404_, _22120_);
  and (_22426_, _22415_, _22393_);
  nor (_22436_, _22415_, _22393_);
  nor (_22447_, _22436_, _22426_);
  not (_22458_, _22447_);
  and (_22469_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_22480_, _22077_, _22055_);
  nor (_22491_, _22480_, _22088_);
  and (_22502_, _22491_, _22469_);
  nor (_22513_, _22491_, _22469_);
  nor (_22523_, _22513_, _22502_);
  not (_22534_, _22523_);
  and (_22545_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_22556_, _22044_, _22022_);
  nor (_22567_, _22556_, _22055_);
  and (_22578_, _22567_, _22545_);
  and (_22589_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_22609_, _22012_, _21990_);
  nor (_22610_, _22609_, _22022_);
  and (_22621_, _22610_, _22589_);
  and (_22632_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_22643_, _21979_, _21957_);
  nor (_22654_, _22643_, _21990_);
  and (_22665_, _22654_, _22632_);
  nor (_22676_, _22610_, _22589_);
  nor (_22686_, _22676_, _22621_);
  and (_22697_, _22686_, _22665_);
  nor (_22718_, _22697_, _22621_);
  not (_22719_, _22718_);
  nor (_22730_, _22567_, _22545_);
  nor (_22741_, _22730_, _22578_);
  and (_22752_, _22741_, _22719_);
  nor (_22763_, _22752_, _22578_);
  nor (_22773_, _22763_, _22534_);
  nor (_22784_, _22773_, _22502_);
  nor (_22795_, _22784_, _22458_);
  nor (_22806_, _22795_, _22426_);
  nor (_22817_, _22806_, _22382_);
  nor (_22828_, _22817_, _22349_);
  nor (_22839_, _22295_, _22273_);
  nor (_22850_, _22839_, _22316_);
  not (_22860_, _22850_);
  nor (_22871_, _22860_, _22828_);
  nor (_22882_, _22871_, _22316_);
  nor (_22893_, _22882_, _22263_);
  nor (_22904_, _22893_, _22230_);
  not (_22915_, _22904_);
  and (_22936_, _22915_, _18409_);
  and (_22937_, _22936_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_22948_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_22958_, _22948_, _22937_);
  and (_22969_, _22958_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_22980_, _22969_, _18398_);
  not (_22991_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_23002_, _18376_, _22991_);
  or (_23013_, _23002_, _22980_);
  nand (_23024_, _22980_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  and (_23035_, _23024_, _23013_);
  and (_24376_, _23035_, _43100_);
  nor (_23056_, _18267_, _18300_);
  and (_23066_, _18267_, _18300_);
  or (_23077_, _23066_, _23056_);
  and (_02359_, _23077_, _43100_);
  and (_23098_, _21935_, _19188_);
  and (_02546_, _23098_, _43100_);
  nor (_23119_, _21946_, _21598_);
  nor (_23130_, _23119_, _21957_);
  and (_02703_, _23130_, _43100_);
  nor (_23151_, _22654_, _22632_);
  nor (_23162_, _23151_, _22665_);
  and (_02884_, _23162_, _43100_);
  nor (_23192_, _22686_, _22665_);
  nor (_23193_, _23192_, _22697_);
  and (_03126_, _23193_, _43100_);
  nor (_23214_, _22741_, _22719_);
  nor (_23225_, _23214_, _22752_);
  and (_03363_, _23225_, _43100_);
  and (_23246_, _22763_, _22534_);
  nor (_23257_, _23246_, _22773_);
  and (_03564_, _23257_, _43100_);
  and (_23277_, _22784_, _22458_);
  nor (_23288_, _23277_, _22795_);
  and (_03763_, _23288_, _43100_);
  and (_23309_, _22806_, _22382_);
  nor (_23320_, _23309_, _22817_);
  and (_03958_, _23320_, _43100_);
  and (_23341_, _22860_, _22828_);
  nor (_23352_, _23341_, _22871_);
  and (_04057_, _23352_, _43100_);
  and (_23373_, _22882_, _22263_);
  nor (_23384_, _23373_, _22893_);
  and (_04156_, _23384_, _43100_);
  nor (_23404_, _22915_, _18409_);
  nor (_23415_, _23404_, _22936_);
  and (_04250_, _23415_, _43100_);
  and (_23436_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_23447_, _23436_, _22936_);
  nor (_23468_, _23447_, _22937_);
  and (_04349_, _23468_, _43100_);
  nor (_23479_, _22948_, _22937_);
  nor (_23490_, _23479_, _22958_);
  and (_04447_, _23490_, _43100_);
  and (_23510_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_23521_, _23510_, _22958_);
  nor (_23532_, _23521_, _22969_);
  and (_04546_, _23532_, _43100_);
  nor (_23553_, _22969_, _18398_);
  nor (_23564_, _23553_, _22980_);
  and (_04645_, _23564_, _43100_);
  and (_23585_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _18201_);
  nor (_23596_, _23585_, _18212_);
  not (_23606_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_23617_, _18234_, _23606_);
  and (_23628_, _23617_, _23596_);
  and (_23639_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_23650_, _23639_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_23661_, _23639_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_23672_, _23661_, _23650_);
  and (_00927_, _23672_, _43100_);
  and (_00957_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _43100_);
  not (_23702_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_23713_, _19977_, _23702_);
  and (_23724_, _19655_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23735_, _23724_, _23713_);
  nor (_23746_, _23735_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_23757_, _19807_, _23702_);
  and (_23767_, _20151_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_23778_, _23767_, _23757_);
  and (_23789_, _23778_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_23800_, _23789_, _23746_);
  nor (_23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_23822_, _23811_, _20325_);
  nor (_23833_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor (_23844_, _23833_, _23822_);
  not (_23854_, _23844_);
  and (_23865_, _18990_, _23702_);
  and (_23876_, _18671_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23897_, _23876_, _23865_);
  nor (_23898_, _23897_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_23909_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_23920_, _18836_, _23702_);
  and (_23930_, _19166_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23941_, _23930_, _23920_);
  nor (_23952_, _23941_, _23909_);
  nor (_23963_, _23952_, _23898_);
  nor (_23974_, _23963_, _23854_);
  and (_23985_, _23963_, _23854_);
  nor (_23996_, _23985_, _23974_);
  and (_24007_, _23811_, _19481_);
  nor (_24017_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor (_24028_, _24017_, _24007_);
  not (_24039_, _24028_);
  nor (_24050_, _19977_, _23702_);
  nor (_24061_, _24050_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24082_, _19655_, _23702_);
  and (_24083_, _19807_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24094_, _24083_, _24082_);
  nor (_24104_, _24094_, _23909_);
  nor (_24115_, _24104_, _24061_);
  nor (_24126_, _24115_, _24039_);
  and (_24137_, _24115_, _24039_);
  nor (_24148_, _24137_, _24126_);
  not (_24159_, _24148_);
  nor (_24170_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and (_24181_, _23811_, _20521_);
  nor (_24191_, _24181_, _24170_);
  not (_24202_, _24191_);
  nor (_24213_, _18990_, _23702_);
  nor (_24224_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24235_, _18671_, _23702_);
  and (_24246_, _18836_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24257_, _24246_, _24235_);
  nor (_24267_, _24257_, _23909_);
  nor (_24278_, _24267_, _24224_);
  nor (_24289_, _24278_, _24202_);
  and (_24300_, _24278_, _24202_);
  and (_24311_, _23735_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24322_, _24311_);
  nor (_24333_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_24344_, _23811_, _20695_);
  nor (_24354_, _24344_, _24333_);
  and (_24365_, _24354_, _24322_);
  and (_24377_, _23897_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24388_, _24377_);
  and (_24399_, _23811_, _21054_);
  nor (_24410_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_24421_, _24410_, _24399_);
  and (_24431_, _24421_, _24388_);
  nor (_24442_, _24421_, _24388_);
  nor (_24453_, _24442_, _24431_);
  not (_24464_, _24453_);
  and (_24475_, _24050_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24486_, _24475_);
  and (_24497_, _23811_, _21555_);
  nor (_24508_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_24518_, _24508_, _24497_);
  and (_24529_, _24518_, _24486_);
  and (_24540_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24551_, _24540_);
  and (_24562_, _23811_, _21381_);
  nor (_24573_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  nor (_24584_, _24573_, _24562_);
  nor (_24595_, _24584_, _24551_);
  not (_24615_, _24595_);
  nor (_24616_, _24518_, _24486_);
  nor (_24627_, _24616_, _24529_);
  and (_24638_, _24627_, _24615_);
  nor (_24649_, _24638_, _24529_);
  nor (_24660_, _24649_, _24464_);
  nor (_24671_, _24660_, _24431_);
  nor (_24681_, _24354_, _24322_);
  nor (_24692_, _24681_, _24365_);
  not (_24703_, _24692_);
  nor (_24714_, _24703_, _24671_);
  nor (_24725_, _24714_, _24365_);
  nor (_24736_, _24725_, _24300_);
  nor (_24747_, _24736_, _24289_);
  nor (_24758_, _24747_, _24159_);
  nor (_24768_, _24758_, _24126_);
  not (_24779_, _24768_);
  and (_24790_, _24779_, _23996_);
  or (_24801_, _24790_, _23974_);
  and (_24812_, _20151_, _19166_);
  or (_24823_, _24812_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_24834_, _23941_);
  and (_24845_, _23778_, _24834_);
  nor (_24856_, _24257_, _24094_);
  and (_24867_, _24856_, _24845_);
  or (_24878_, _24867_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24889_, _24878_, _24823_);
  and (_24900_, _24889_, _24801_);
  and (_24911_, _24900_, _23800_);
  nor (_24922_, _24779_, _23996_);
  or (_24933_, _24922_, _24790_);
  and (_24944_, _24933_, _24911_);
  nor (_24955_, _24911_, _23844_);
  nor (_24966_, _24955_, _24944_);
  not (_24977_, _24966_);
  and (_24988_, _24966_, _23800_);
  not (_24999_, _23963_);
  nor (_25010_, _24911_, _24039_);
  and (_25021_, _24747_, _24159_);
  nor (_25031_, _25021_, _24758_);
  and (_25042_, _25031_, _24911_);
  or (_25053_, _25042_, _25010_);
  and (_25064_, _25053_, _24999_);
  nor (_25075_, _25053_, _24999_);
  nor (_25086_, _25075_, _25064_);
  not (_25097_, _25086_);
  not (_25108_, _24115_);
  nor (_25119_, _24911_, _24202_);
  nor (_25130_, _24300_, _24289_);
  nor (_25141_, _25130_, _24725_);
  and (_25162_, _25130_, _24725_);
  or (_25163_, _25162_, _25141_);
  and (_25174_, _25163_, _24911_);
  or (_25185_, _25174_, _25119_);
  and (_25196_, _25185_, _25108_);
  nor (_25207_, _25185_, _25108_);
  not (_25218_, _24278_);
  and (_25229_, _24703_, _24671_);
  or (_25240_, _25229_, _24714_);
  and (_25251_, _25240_, _24911_);
  nor (_25262_, _24911_, _24354_);
  nor (_25273_, _25262_, _25251_);
  and (_25284_, _25273_, _25218_);
  and (_25295_, _24649_, _24464_);
  nor (_25306_, _25295_, _24660_);
  not (_25317_, _25306_);
  and (_25328_, _25317_, _24911_);
  nor (_25339_, _24911_, _24421_);
  nor (_25350_, _25339_, _25328_);
  and (_25361_, _25350_, _24322_);
  nor (_25372_, _25350_, _24322_);
  nor (_25383_, _25372_, _25361_);
  not (_25394_, _25383_);
  nor (_25404_, _24627_, _24615_);
  nor (_25425_, _25404_, _24638_);
  not (_25426_, _25425_);
  and (_25437_, _25426_, _24911_);
  nor (_25448_, _24911_, _24518_);
  nor (_25459_, _25448_, _25437_);
  and (_25470_, _25459_, _24388_);
  and (_25481_, _24911_, _24540_);
  nor (_25492_, _25481_, _24584_);
  and (_25503_, _25481_, _24584_);
  nor (_25514_, _25503_, _25492_);
  and (_25525_, _25514_, _24486_);
  nor (_25536_, _25514_, _24486_);
  nor (_25547_, _25536_, _25525_);
  and (_25558_, _23811_, _21925_);
  nor (_25569_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_25580_, _25569_, _25558_);
  nor (_25591_, _25580_, _24551_);
  not (_25602_, _25591_);
  and (_25613_, _25602_, _25547_);
  nor (_25624_, _25613_, _25525_);
  nor (_25635_, _25459_, _24388_);
  nor (_25646_, _25635_, _25470_);
  not (_25657_, _25646_);
  nor (_25668_, _25657_, _25624_);
  nor (_25679_, _25668_, _25470_);
  nor (_25690_, _25679_, _25394_);
  nor (_25701_, _25690_, _25361_);
  nor (_25712_, _25273_, _25218_);
  nor (_25733_, _25712_, _25284_);
  not (_25734_, _25733_);
  nor (_25745_, _25734_, _25701_);
  nor (_25755_, _25745_, _25284_);
  nor (_25766_, _25755_, _25207_);
  nor (_25777_, _25766_, _25196_);
  nor (_25788_, _25777_, _25097_);
  or (_25799_, _25788_, _25064_);
  or (_25810_, _25799_, _24988_);
  and (_25821_, _25810_, _24889_);
  nor (_25832_, _25821_, _24977_);
  and (_25843_, _24988_, _24889_);
  and (_25854_, _25843_, _25799_);
  or (_25865_, _25854_, _25832_);
  and (_00976_, _25865_, _43100_);
  or (_25886_, _24966_, _23800_);
  and (_25897_, _25886_, _25821_);
  and (_02839_, _25897_, _43100_);
  and (_02851_, _24911_, _43100_);
  and (_02873_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _43100_);
  and (_02897_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _43100_);
  and (_02919_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _43100_);
  or (_25958_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_25969_, _23639_, rst);
  and (_02931_, _25969_, _25958_);
  and (_25990_, _25897_, _24540_);
  or (_26001_, _25990_, _25580_);
  nand (_26012_, _25990_, _25580_);
  and (_26023_, _26012_, _26001_);
  and (_02944_, _26023_, _43100_);
  nor (_26054_, _25602_, _25547_);
  or (_26055_, _26054_, _25613_);
  nand (_26066_, _26055_, _25897_);
  or (_26077_, _25897_, _25514_);
  and (_26088_, _26077_, _26066_);
  and (_02957_, _26088_, _43100_);
  and (_26108_, _25657_, _25624_);
  or (_26119_, _26108_, _25668_);
  nand (_26130_, _26119_, _25897_);
  or (_26141_, _25897_, _25459_);
  and (_26152_, _26141_, _26130_);
  and (_02969_, _26152_, _43100_);
  and (_26173_, _25679_, _25394_);
  or (_26184_, _26173_, _25690_);
  nand (_26195_, _26184_, _25897_);
  or (_26206_, _25897_, _25350_);
  and (_26217_, _26206_, _26195_);
  and (_02980_, _26217_, _43100_);
  and (_26238_, _25734_, _25701_);
  or (_26249_, _26238_, _25745_);
  nand (_26260_, _26249_, _25897_);
  or (_26271_, _25897_, _25273_);
  and (_26282_, _26271_, _26260_);
  and (_02994_, _26282_, _43100_);
  or (_26303_, _25207_, _25196_);
  and (_26314_, _26303_, _25755_);
  nor (_26325_, _26303_, _25755_);
  or (_26336_, _26325_, _26314_);
  nand (_26347_, _26336_, _25897_);
  or (_26358_, _25897_, _25185_);
  and (_26369_, _26358_, _26347_);
  and (_03006_, _26369_, _43100_);
  and (_26390_, _25777_, _25097_);
  or (_26401_, _26390_, _25788_);
  nand (_26412_, _26401_, _25897_);
  or (_26423_, _25897_, _25053_);
  and (_26433_, _26423_, _26412_);
  and (_03020_, _26433_, _43100_);
  not (_26454_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_26465_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _18201_);
  and (_26476_, _26465_, _26454_);
  and (_26487_, _26476_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_26498_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_26509_, _26498_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_26530_, _26498_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_26531_, _26530_, _26509_);
  and (_26542_, _26531_, _26487_);
  not (_26553_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_26564_, _26476_, _26553_);
  and (_26575_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_26586_, _26575_, _26542_);
  not (_26597_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_26608_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _18201_);
  and (_26619_, _26608_, _26597_);
  and (_26630_, _26619_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_26641_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_26652_, _26619_, _26454_);
  and (_26663_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or (_26674_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_26685_, _26674_, _18201_);
  nor (_26696_, _26685_, _26608_);
  and (_26707_, _26696_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_26718_, _26707_, _26663_);
  nor (_26729_, _26718_, _26641_);
  and (_26740_, _26729_, _26586_);
  and (_26761_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor (_26762_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_26773_, _26762_, _26498_);
  and (_26784_, _26773_, _26487_);
  nor (_26794_, _26784_, _26761_);
  and (_26805_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_26816_, _26696_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_26827_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_26838_, _26827_, _26816_);
  nor (_26849_, _26838_, _26805_);
  and (_26860_, _26849_, _26794_);
  and (_26871_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_26882_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_26893_, _26882_, _26871_);
  and (_26904_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not (_26915_, _26904_);
  not (_26926_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_26937_, _26487_, _26926_);
  and (_26948_, _26696_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_26959_, _26948_, _26937_);
  and (_26970_, _26959_, _26915_);
  and (_26981_, _26970_, _26893_);
  and (_26992_, _26981_, _26860_);
  and (_27003_, _26992_, _26740_);
  and (_27014_, _26509_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_27025_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_27036_, _27025_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_27047_, _27036_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_27058_, _27047_);
  not (_27069_, _26487_);
  nor (_27080_, _27036_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_27091_, _27080_, _27069_);
  and (_27102_, _27091_, _27058_);
  not (_27113_, _27102_);
  and (_27124_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27134_, _27124_, _26465_);
  and (_27145_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_27156_, _27145_, _27134_);
  and (_27167_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_27178_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_27189_, _27178_, _27167_);
  and (_27200_, _27189_, _27156_);
  and (_27211_, _27200_, _27113_);
  nor (_27222_, _27025_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_27233_, _27222_);
  nor (_27244_, _27036_, _27069_);
  and (_27255_, _27244_, _27233_);
  not (_27266_, _27255_);
  and (_27277_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_27288_, _27277_, _27134_);
  and (_27299_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_27310_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_27321_, _27310_, _27299_);
  and (_27342_, _27321_, _27288_);
  and (_27343_, _27342_, _27266_);
  nor (_27354_, _27343_, _27211_);
  not (_27365_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_27376_, _27047_, _27365_);
  and (_27387_, _27047_, _27365_);
  nor (_27398_, _27387_, _27376_);
  nor (_27409_, _27398_, _27069_);
  not (_27420_, _27409_);
  and (_27431_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_27442_, _27431_, _27134_);
  and (_27453_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_27464_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_27475_, _27464_, _27453_);
  and (_27485_, _27475_, _27442_);
  and (_27496_, _27485_, _27420_);
  not (_27507_, _27496_);
  and (_27518_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_27529_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_27540_, _27529_, _27518_);
  not (_27551_, _27014_);
  nor (_27562_, _26509_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_27573_, _27562_, _27069_);
  and (_27584_, _27573_, _27551_);
  and (_27595_, _26696_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_27606_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_27617_, _27606_, _27595_);
  not (_27628_, _27617_);
  nor (_27639_, _27628_, _27584_);
  and (_27650_, _27639_, _27540_);
  not (_27661_, _27650_);
  and (_27672_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_27683_, _27672_, _27134_);
  and (_27694_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_27705_, _27694_);
  and (_27716_, _27705_, _27683_);
  nor (_27727_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_27738_, _27727_);
  nor (_27749_, _27025_, _27069_);
  and (_27760_, _27749_, _27738_);
  and (_27771_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and (_27782_, _26696_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_27793_, _27782_, _27771_);
  not (_27804_, _27793_);
  nor (_27814_, _27804_, _27760_);
  and (_27825_, _27814_, _27716_);
  nor (_27836_, _27825_, _27661_);
  and (_27847_, _27836_, _27507_);
  and (_27858_, _27847_, _27354_);
  nand (_27869_, _27858_, _27003_);
  and (_27880_, _25865_, _23628_);
  not (_27891_, _27880_);
  and (_27902_, _23035_, _18267_);
  not (_27913_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_27924_, _18212_, _27913_);
  and (_27935_, _27924_, _18256_);
  not (_27946_, _27935_);
  nor (_27957_, _20325_, _20151_);
  and (_27978_, _20325_, _20151_);
  nor (_27979_, _27978_, _27957_);
  not (_27990_, _19166_);
  nor (_28001_, _19481_, _27990_);
  nor (_28012_, _19481_, _19166_);
  and (_28023_, _19481_, _19166_);
  nor (_28034_, _28023_, _28012_);
  not (_28045_, _19807_);
  nor (_28056_, _20521_, _28045_);
  nor (_28067_, _20521_, _19807_);
  and (_28078_, _20521_, _19807_);
  nor (_28089_, _28078_, _28067_);
  not (_28100_, _18836_);
  and (_28111_, _20695_, _28100_);
  nor (_28122_, _28111_, _28089_);
  nor (_28132_, _28122_, _28056_);
  nor (_28143_, _28132_, _28034_);
  nor (_28154_, _28143_, _28001_);
  and (_28165_, _28132_, _28034_);
  nor (_28176_, _28165_, _28143_);
  not (_28187_, _28176_);
  and (_28198_, _28111_, _28089_);
  nor (_28209_, _28198_, _28122_);
  not (_28220_, _28209_);
  nor (_28231_, _20695_, _18836_);
  and (_28242_, _20695_, _18836_);
  nor (_28253_, _28242_, _28231_);
  not (_28264_, _28253_);
  and (_28285_, _21054_, _19655_);
  nor (_28286_, _21054_, _19655_);
  nor (_28297_, _28286_, _28285_);
  nor (_28308_, _21555_, _18671_);
  and (_28319_, _21555_, _18671_);
  nor (_28330_, _28319_, _28308_);
  nor (_28341_, _21381_, _19977_);
  and (_28352_, _21381_, _19977_);
  nor (_28363_, _28352_, _28341_);
  not (_28374_, _18990_);
  and (_28385_, _21925_, _28374_);
  nor (_28396_, _28385_, _28363_);
  not (_28407_, _19977_);
  nor (_28418_, _21381_, _28407_);
  nor (_28429_, _28418_, _28396_);
  nor (_28440_, _28429_, _28330_);
  not (_28450_, _18671_);
  nor (_28461_, _21555_, _28450_);
  nor (_28472_, _28461_, _28440_);
  nor (_28483_, _28472_, _28297_);
  and (_28494_, _28472_, _28297_);
  nor (_28505_, _28494_, _28483_);
  not (_28516_, _28505_);
  and (_28527_, _28429_, _28330_);
  nor (_28538_, _28527_, _28440_);
  not (_28549_, _28538_);
  and (_28560_, _28385_, _28363_);
  nor (_28571_, _28560_, _28396_);
  not (_28582_, _28571_);
  nor (_28593_, _21925_, _18990_);
  and (_28604_, _21925_, _18990_);
  nor (_28615_, _28604_, _28593_);
  not (_28636_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_28637_, _18475_, _28636_);
  not (_28648_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_28659_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28670_, _28659_, _20043_);
  nor (_28681_, _28670_, _28648_);
  nor (_28692_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28703_, _28692_, _18716_);
  not (_28714_, _28703_);
  not (_28725_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28736_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _28725_);
  and (_28746_, _28736_, _19699_);
  not (_28757_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_28768_, _28757_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28779_, _28768_, _19056_);
  nor (_28790_, _28779_, _28746_);
  and (_28801_, _28790_, _28714_);
  and (_28812_, _28801_, _28681_);
  and (_28823_, _28659_, _19547_);
  nor (_28834_, _28823_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_28845_, _28768_, _18518_);
  not (_28856_, _28845_);
  and (_28867_, _28736_, _19874_);
  and (_28878_, _28692_, _18880_);
  nor (_28889_, _28878_, _28867_);
  and (_28900_, _28889_, _28856_);
  and (_28911_, _28900_, _28834_);
  nor (_28922_, _28911_, _28812_);
  nor (_28933_, _28922_, _18475_);
  nor (_28944_, _28933_, _28637_);
  and (_28955_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_28966_, _28955_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_28977_, _28966_);
  and (_28988_, _28977_, _28944_);
  and (_29009_, _28977_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_29010_, _29009_, _28988_);
  nor (_29021_, _29010_, _28615_);
  and (_29032_, _29021_, _28582_);
  and (_29043_, _29032_, _28549_);
  and (_29054_, _29043_, _28516_);
  not (_29064_, _19655_);
  or (_29075_, _21054_, _29064_);
  and (_29086_, _21054_, _29064_);
  or (_29097_, _28472_, _29086_);
  and (_29108_, _29097_, _29075_);
  or (_29119_, _29108_, _29054_);
  and (_29130_, _29119_, _28264_);
  and (_29141_, _29130_, _28220_);
  and (_29152_, _29141_, _28187_);
  nor (_29163_, _29152_, _28154_);
  nor (_29174_, _29163_, _27979_);
  and (_29185_, _29163_, _27979_);
  nor (_29196_, _29185_, _29174_);
  nor (_29207_, _29196_, _27946_);
  not (_29218_, _29207_);
  not (_29229_, _27979_);
  not (_29240_, _28034_);
  and (_29251_, _28231_, _28089_);
  nor (_29262_, _29251_, _28067_);
  nor (_29273_, _29262_, _29240_);
  not (_29284_, _28330_);
  and (_29295_, _28593_, _28363_);
  nor (_29306_, _29295_, _28341_);
  nor (_29317_, _29306_, _29284_);
  nor (_29328_, _29317_, _28308_);
  nor (_29339_, _29328_, _28297_);
  and (_29350_, _29328_, _28297_);
  nor (_29361_, _29350_, _29339_);
  not (_29371_, _28615_);
  nor (_29382_, _29010_, _29371_);
  and (_29393_, _29382_, _28363_);
  and (_29404_, _29306_, _29284_);
  nor (_29415_, _29404_, _29317_);
  and (_29426_, _29415_, _29393_);
  not (_29437_, _29426_);
  nor (_29448_, _29437_, _29361_);
  nor (_29459_, _29328_, _28285_);
  or (_29470_, _29459_, _28286_);
  or (_29481_, _29470_, _29448_);
  and (_29492_, _29481_, _28253_);
  and (_29503_, _29492_, _28089_);
  and (_29514_, _29262_, _29240_);
  nor (_29535_, _29514_, _29273_);
  and (_29536_, _29535_, _29503_);
  or (_29547_, _29536_, _29273_);
  nor (_29558_, _29547_, _28012_);
  and (_29569_, _29558_, _29229_);
  nor (_29580_, _29558_, _29229_);
  not (_29591_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_29602_, _23585_, _29591_);
  and (_29613_, _29602_, _18256_);
  not (_29624_, _29613_);
  or (_29635_, _29624_, _29580_);
  nor (_29646_, _29635_, _29569_);
  and (_29657_, _18245_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_29668_, _29657_, _27924_);
  nor (_29678_, _21925_, _21381_);
  and (_29689_, _29678_, _21566_);
  and (_29700_, _29689_, _21065_);
  and (_29711_, _29700_, _20706_);
  and (_29722_, _29711_, _20532_);
  and (_29733_, _29722_, _19492_);
  and (_29744_, _29733_, _29010_);
  not (_29755_, _29010_);
  and (_29766_, _19481_, _20521_);
  and (_29777_, _21555_, _21381_);
  and (_29788_, _29777_, _21925_);
  and (_29808_, _29788_, _21054_);
  and (_29809_, _29808_, _20695_);
  and (_29820_, _29809_, _29766_);
  and (_29831_, _29820_, _29755_);
  nor (_29842_, _29831_, _29744_);
  and (_29853_, _29842_, _20325_);
  nor (_29864_, _29842_, _20325_);
  nor (_29875_, _29864_, _29853_);
  and (_29886_, _29875_, _29668_);
  not (_29897_, _20151_);
  nor (_29908_, _29010_, _29897_);
  not (_29919_, _29908_);
  and (_29930_, _29010_, _20325_);
  and (_29941_, _29657_, _18223_);
  not (_29951_, _29941_);
  nor (_29962_, _29951_, _29930_);
  and (_29973_, _29962_, _29919_);
  nor (_29984_, _29973_, _29886_);
  and (_29995_, _29602_, _23617_);
  nor (_30006_, _29777_, _21054_);
  and (_30017_, _30006_, _29995_);
  and (_30028_, _30017_, _20706_);
  nor (_30039_, _30028_, _20532_);
  and (_30050_, _30039_, _19481_);
  nor (_30061_, _29766_, _20325_);
  nor (_30072_, _30061_, _30017_);
  and (_30083_, _30072_, _29010_);
  nor (_30093_, _30083_, _30050_);
  nor (_30104_, _30093_, _20336_);
  and (_30115_, _30093_, _20336_);
  nor (_30126_, _30115_, _30104_);
  and (_30137_, _30126_, _29995_);
  and (_30148_, _29657_, _29602_);
  not (_30159_, _30148_);
  nor (_30170_, _30159_, _29010_);
  not (_30181_, _30170_);
  not (_30192_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_30203_, _18245_, _30192_);
  and (_30214_, _30203_, _29602_);
  not (_30225_, _30214_);
  nor (_30235_, _30225_, _27978_);
  and (_30246_, _30203_, _23596_);
  and (_30257_, _30246_, _27979_);
  nor (_30268_, _30257_, _30235_);
  and (_30279_, _23617_, _18223_);
  and (_30290_, _30279_, _27957_);
  and (_30301_, _27924_, _23617_);
  and (_30312_, _30301_, _20325_);
  nor (_30323_, _30312_, _30290_);
  and (_30334_, _30203_, _18212_);
  not (_30345_, _30334_);
  nor (_30356_, _30345_, _19481_);
  not (_30367_, _30356_);
  and (_30377_, _23596_, _18256_);
  not (_30388_, _30377_);
  nor (_30399_, _30388_, _20325_);
  and (_30410_, _29657_, _23596_);
  and (_30431_, _30410_, _21935_);
  nor (_30432_, _30431_, _30399_);
  and (_30443_, _30432_, _30367_);
  and (_30454_, _30443_, _30323_);
  and (_30465_, _30454_, _30268_);
  and (_30476_, _30465_, _30181_);
  not (_30487_, _30476_);
  nor (_30498_, _30487_, _30137_);
  and (_30509_, _30498_, _29984_);
  not (_30519_, _30509_);
  nor (_30530_, _30519_, _29646_);
  and (_30541_, _30530_, _29218_);
  not (_30552_, _30541_);
  nor (_30563_, _30552_, _27902_);
  and (_30574_, _30563_, _27891_);
  not (_30585_, _30574_);
  or (_30596_, _30585_, _27869_);
  not (_30607_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_30618_, \oc8051_top_1.oc8051_decoder1.wr , _18201_);
  not (_30629_, _30618_);
  nor (_30640_, _30629_, _26476_);
  and (_30651_, _30640_, _30607_);
  not (_30661_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_30672_, _27869_, _30661_);
  and (_30683_, _30672_, _30651_);
  and (_30694_, _30683_, _30596_);
  nor (_30705_, _30640_, _30661_);
  nor (_30716_, _29580_, _27957_);
  nor (_30727_, _30716_, _29624_);
  not (_30738_, _30727_);
  and (_30749_, _20325_, _29897_);
  nor (_30759_, _30749_, _29174_);
  nor (_30770_, _30759_, _27946_);
  and (_30781_, _29010_, _19481_);
  and (_30792_, _30781_, _30039_);
  nor (_30803_, _30792_, _29930_);
  not (_30814_, _29995_);
  nor (_30825_, _29010_, _20325_);
  not (_30836_, _30825_);
  nor (_30847_, _30836_, _30050_);
  nor (_30858_, _30847_, _30814_);
  and (_30869_, _30858_, _30803_);
  not (_30879_, _30869_);
  nor (_30890_, _29009_, _28944_);
  not (_30901_, _30246_);
  nor (_30912_, _30901_, _28988_);
  nor (_30923_, _30912_, _30214_);
  nor (_30934_, _30923_, _30890_);
  not (_30945_, _30934_);
  nor (_30956_, _30388_, _29010_);
  not (_30967_, _30956_);
  and (_30978_, _28966_, _28944_);
  and (_30988_, _30203_, _27924_);
  and (_30999_, _30279_, _28944_);
  nor (_31010_, _30999_, _30988_);
  nor (_31021_, _31010_, _30978_);
  not (_31032_, _31021_);
  not (_31043_, _29009_);
  and (_31054_, _30301_, _31043_);
  and (_31065_, _30410_, _29009_);
  nor (_31076_, _31065_, _31054_);
  nor (_31087_, _31076_, _28988_);
  not (_31097_, _31087_);
  nor (_31108_, _30159_, _21925_);
  and (_31119_, _30203_, _18223_);
  not (_31141_, _31119_);
  nor (_31142_, _31141_, _20325_);
  nor (_31164_, _31142_, _31108_);
  not (_31165_, _31164_);
  nor (_31187_, _31165_, _30017_);
  and (_31188_, _31187_, _31097_);
  and (_31210_, _31188_, _31032_);
  and (_31211_, _31210_, _30967_);
  and (_31221_, _31211_, _30945_);
  and (_31232_, _31221_, _30879_);
  not (_31243_, _31232_);
  nor (_31264_, _31243_, _30770_);
  and (_31265_, _31264_, _30738_);
  not (_31286_, _26740_);
  nor (_31287_, _26981_, _26860_);
  and (_31308_, _31287_, _31286_);
  and (_31309_, _31308_, _27858_);
  nand (_31329_, _31309_, _31265_);
  or (_31330_, _31309_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_31351_, _30640_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_31352_, _31351_, _31330_);
  and (_31373_, _31352_, _31329_);
  or (_31374_, _31373_, _30705_);
  or (_31395_, _31374_, _30694_);
  and (_06664_, _31395_, _43100_);
  and (_31416_, _26023_, _23628_);
  not (_31417_, _31416_);
  and (_31437_, _23352_, _18267_);
  and (_31438_, _29010_, _29371_);
  nor (_31459_, _31438_, _29382_);
  not (_31460_, _31459_);
  nor (_31481_, _29613_, _27935_);
  nor (_31482_, _31481_, _31460_);
  nor (_31503_, _31141_, _29010_);
  not (_31504_, _31503_);
  nor (_31525_, _30901_, _28593_);
  nor (_31526_, _31525_, _30214_);
  or (_31546_, _31526_, _28604_);
  and (_31547_, _29657_, _29591_);
  not (_31568_, _31547_);
  nor (_31569_, _31568_, _21381_);
  and (_31590_, _30988_, _20336_);
  nor (_31591_, _31590_, _31569_);
  and (_31612_, _30279_, _28593_);
  and (_31613_, _30301_, _21925_);
  nor (_31634_, _31613_, _31612_);
  nor (_31635_, _29951_, _18990_);
  and (_31655_, _29668_, _21925_);
  nor (_31656_, _31655_, _31635_);
  nor (_31677_, _30377_, _29995_);
  nor (_31678_, _31677_, _21925_);
  not (_31699_, _31678_);
  and (_31700_, _31699_, _31656_);
  and (_31721_, _31700_, _31634_);
  and (_31722_, _31721_, _31591_);
  and (_31743_, _31722_, _31546_);
  and (_31744_, _31743_, _31504_);
  not (_31764_, _31744_);
  nor (_31765_, _31764_, _31482_);
  not (_31786_, _31765_);
  nor (_31787_, _31786_, _31437_);
  and (_31808_, _31787_, _31417_);
  not (_31809_, _31808_);
  or (_31830_, _31809_, _27869_);
  not (_31831_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_31852_, _27869_, _31831_);
  and (_31853_, _31852_, _30651_);
  and (_31864_, _31853_, _31830_);
  nor (_31874_, _30640_, _31831_);
  not (_31885_, _31265_);
  or (_31896_, _31885_, _27869_);
  and (_31907_, _31852_, _31351_);
  and (_31918_, _31907_, _31896_);
  or (_31929_, _31918_, _31874_);
  or (_31940_, _31929_, _31864_);
  and (_08905_, _31940_, _43100_);
  and (_31961_, _23384_, _18267_);
  not (_31972_, _31961_);
  and (_31982_, _26088_, _23628_);
  nor (_31993_, _28593_, _28363_);
  or (_32004_, _31993_, _29295_);
  and (_32015_, _32004_, _29382_);
  nor (_32026_, _32004_, _29382_);
  or (_32037_, _32026_, _32015_);
  and (_32048_, _32037_, _29613_);
  nor (_32059_, _29021_, _28582_);
  nor (_32070_, _32059_, _29032_);
  nor (_32081_, _32070_, _27946_);
  not (_32091_, _32081_);
  nor (_32102_, _30006_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_32113_, _32102_, _21392_);
  nor (_32124_, _32102_, _21392_);
  nor (_32135_, _32124_, _32113_);
  nor (_32146_, _32135_, _30814_);
  not (_32157_, _32146_);
  and (_32168_, _30246_, _28363_);
  nor (_32179_, _30225_, _28352_);
  not (_32190_, _32179_);
  and (_32200_, _30279_, _28341_);
  and (_32211_, _30301_, _21381_);
  nor (_32222_, _32211_, _32200_);
  nand (_32233_, _32222_, _32190_);
  nor (_32244_, _32233_, _32168_);
  nor (_32255_, _30345_, _21925_);
  not (_32266_, _32255_);
  nor (_32277_, _30388_, _21381_);
  nor (_32288_, _31568_, _21555_);
  nor (_32299_, _32288_, _32277_);
  and (_32309_, _32299_, _32266_);
  and (_32320_, _32309_, _32244_);
  and (_32331_, _32320_, _32157_);
  and (_32342_, _32331_, _32091_);
  nor (_32353_, _29951_, _19977_);
  and (_32364_, _21925_, _21381_);
  nor (_32375_, _32364_, _29678_);
  not (_32386_, _32375_);
  nor (_32397_, _32386_, _29010_);
  and (_32408_, _32386_, _29010_);
  nor (_32418_, _32408_, _32397_);
  and (_32429_, _32418_, _29668_);
  nor (_32440_, _32429_, _32353_);
  nand (_32451_, _32440_, _32342_);
  nor (_32462_, _32451_, _32048_);
  not (_32473_, _32462_);
  nor (_32484_, _32473_, _31982_);
  and (_32495_, _32484_, _31972_);
  not (_32506_, _32495_);
  or (_32517_, _32506_, _27869_);
  not (_32527_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_32538_, _27869_, _32527_);
  and (_32549_, _32538_, _30651_);
  and (_32560_, _32549_, _32517_);
  nor (_32571_, _30640_, _32527_);
  not (_32582_, _26981_);
  and (_32593_, _32582_, _26860_);
  and (_32604_, _32593_, _26740_);
  and (_32615_, _32604_, _27858_);
  nand (_32626_, _32615_, _31265_);
  or (_32636_, _32615_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_32647_, _32636_, _31351_);
  and (_32658_, _32647_, _32626_);
  or (_32669_, _32658_, _32571_);
  or (_32680_, _32669_, _32560_);
  and (_08916_, _32680_, _43100_);
  and (_32701_, _26152_, _23628_);
  not (_32712_, _32701_);
  and (_32723_, _23415_, _18267_);
  nor (_32734_, _29951_, _18671_);
  nor (_32744_, _32364_, _29010_);
  nor (_32755_, _29678_, _29755_);
  nor (_32766_, _32755_, _32744_);
  and (_32777_, _32766_, _21566_);
  not (_32788_, _32777_);
  not (_32799_, _29668_);
  nor (_32810_, _32766_, _21566_);
  nor (_32821_, _32810_, _32799_);
  and (_32832_, _32821_, _32788_);
  nor (_32843_, _32832_, _32734_);
  nor (_32854_, _29032_, _28549_);
  nor (_32864_, _32854_, _29043_);
  nor (_32875_, _32864_, _27946_);
  and (_32886_, _30246_, _28330_);
  nor (_32897_, _30225_, _28319_);
  not (_32908_, _32897_);
  and (_32919_, _30279_, _28308_);
  and (_32930_, _30301_, _21555_);
  nor (_32941_, _32930_, _32919_);
  nand (_32952_, _32941_, _32908_);
  nor (_32963_, _32952_, _32886_);
  nor (_32973_, _30345_, _21381_);
  not (_32984_, _32973_);
  nor (_32995_, _30388_, _21555_);
  nor (_33006_, _31568_, _21054_);
  nor (_33017_, _33006_, _32995_);
  and (_33028_, _33017_, _32984_);
  and (_33039_, _33028_, _32963_);
  not (_33050_, _33039_);
  nor (_33061_, _33050_, _32875_);
  nor (_33071_, _29415_, _29393_);
  nor (_33082_, _33071_, _29624_);
  and (_33093_, _33082_, _29437_);
  and (_33104_, _29777_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_33115_, _32124_, _21555_);
  nor (_33126_, _33115_, _33104_);
  nor (_33137_, _33126_, _30814_);
  nor (_33148_, _33137_, _33093_);
  and (_33159_, _33148_, _33061_);
  and (_33170_, _33159_, _32843_);
  not (_33180_, _33170_);
  nor (_33191_, _33180_, _32723_);
  and (_33202_, _33191_, _32712_);
  not (_33213_, _33202_);
  or (_33224_, _33213_, _27869_);
  not (_33235_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_33246_, _27869_, _33235_);
  and (_33257_, _33246_, _30651_);
  and (_33268_, _33257_, _33224_);
  nor (_33279_, _30640_, _33235_);
  nand (_33289_, _27858_, _26740_);
  or (_33300_, _31287_, _33289_);
  and (_33311_, _33300_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_33322_, _26860_);
  and (_33333_, _26740_, _26981_);
  and (_33344_, _33333_, _33322_);
  not (_33355_, _33344_);
  nor (_33366_, _33355_, _31265_);
  and (_33377_, _26740_, _26860_);
  and (_33388_, _33377_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_33399_, _33388_, _33366_);
  and (_33409_, _33399_, _27858_);
  or (_33420_, _33409_, _33311_);
  and (_33431_, _33420_, _31351_);
  or (_33442_, _33431_, _33279_);
  or (_33453_, _33442_, _33268_);
  and (_08927_, _33453_, _43100_);
  and (_33474_, _26217_, _23628_);
  not (_33485_, _33474_);
  not (_33496_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_33507_, _29777_, _33496_);
  nor (_33517_, _33507_, _21065_);
  nor (_33528_, _30388_, _21054_);
  nor (_33539_, _30006_, _30814_);
  nor (_33550_, _33539_, _33528_);
  nor (_33561_, _33550_, _33517_);
  not (_33572_, _33561_);
  nor (_33583_, _30225_, _28285_);
  and (_33594_, _30246_, _28297_);
  nor (_33605_, _33594_, _33583_);
  and (_33616_, _30279_, _28286_);
  and (_33626_, _30301_, _21054_);
  nor (_33637_, _33626_, _33616_);
  nor (_33648_, _31568_, _20695_);
  nor (_33659_, _30345_, _21555_);
  nor (_33670_, _33659_, _33648_);
  and (_33681_, _33670_, _33637_);
  and (_33692_, _33681_, _33605_);
  and (_33703_, _33692_, _33572_);
  nor (_33714_, _29043_, _28516_);
  nor (_33725_, _33714_, _29054_);
  nor (_33735_, _33725_, _27946_);
  and (_33746_, _29437_, _29361_);
  or (_33757_, _33746_, _29624_);
  nor (_33768_, _33757_, _29448_);
  nor (_33779_, _33768_, _33735_);
  and (_33790_, _33779_, _33703_);
  and (_33801_, _23468_, _18267_);
  not (_33812_, _33801_);
  nor (_33823_, _29951_, _19655_);
  and (_33833_, _29689_, _29010_);
  and (_33844_, _29788_, _29755_);
  nor (_33855_, _33844_, _33833_);
  nor (_33866_, _33855_, _21054_);
  not (_33877_, _33866_);
  and (_33888_, _33855_, _21054_);
  nor (_33899_, _33888_, _32799_);
  and (_33910_, _33899_, _33877_);
  nor (_33921_, _33910_, _33823_);
  and (_33932_, _33921_, _33812_);
  and (_33943_, _33932_, _33790_);
  and (_33953_, _33943_, _33485_);
  not (_33964_, _33953_);
  or (_33975_, _33964_, _27869_);
  not (_33986_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_33997_, _27869_, _33986_);
  and (_34008_, _33997_, _30651_);
  and (_34019_, _34008_, _33975_);
  nor (_34030_, _30640_, _33986_);
  and (_34041_, _33289_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_34052_, _31287_, _26740_);
  and (_34062_, _34052_, _31885_);
  nor (_34073_, _33377_, _33333_);
  nor (_34084_, _34073_, _33986_);
  or (_34095_, _34084_, _34062_);
  and (_34106_, _34095_, _27858_);
  or (_34117_, _34106_, _34041_);
  and (_34128_, _34117_, _31351_);
  or (_34139_, _34128_, _34030_);
  or (_34150_, _34139_, _34019_);
  and (_08938_, _34150_, _43100_);
  and (_34170_, _23490_, _18267_);
  not (_34181_, _34170_);
  and (_34192_, _26282_, _23628_);
  nor (_34203_, _29010_, _18836_);
  and (_34214_, _29010_, _20706_);
  nor (_34225_, _34214_, _34203_);
  nor (_34236_, _34225_, _29951_);
  and (_34247_, _29700_, _29010_);
  and (_34258_, _29808_, _29755_);
  nor (_34269_, _34258_, _34247_);
  and (_34281_, _34269_, _20695_);
  nor (_34300_, _34269_, _20695_);
  nor (_34311_, _34300_, _34281_);
  and (_34322_, _34311_, _29668_);
  nor (_34333_, _34322_, _34236_);
  and (_34344_, _30279_, _28231_);
  and (_34355_, _30301_, _20695_);
  nor (_34366_, _34355_, _34344_);
  nor (_34377_, _31568_, _20521_);
  not (_34388_, _34377_);
  and (_34398_, _34388_, _34366_);
  nor (_34409_, _30017_, _20706_);
  not (_34420_, _34409_);
  nor (_34431_, _30028_, _30814_);
  and (_34442_, _34431_, _34420_);
  nor (_34453_, _30225_, _28242_);
  and (_34464_, _30246_, _28253_);
  nor (_34475_, _34464_, _34453_);
  nor (_34486_, _30345_, _21054_);
  nor (_34497_, _30388_, _20695_);
  nor (_34507_, _34497_, _34486_);
  nand (_34518_, _34507_, _34475_);
  nor (_34529_, _34518_, _34442_);
  and (_34540_, _34529_, _34398_);
  nor (_34551_, _29119_, _28253_);
  and (_34562_, _29119_, _28253_);
  nor (_34573_, _34562_, _34551_);
  and (_34584_, _34573_, _27935_);
  nor (_34595_, _29481_, _28253_);
  not (_34606_, _34595_);
  nor (_34616_, _29624_, _29492_);
  and (_34627_, _34616_, _34606_);
  nor (_34638_, _34627_, _34584_);
  and (_34649_, _34638_, _34540_);
  and (_34660_, _34649_, _34333_);
  not (_34671_, _34660_);
  nor (_34682_, _34671_, _34192_);
  and (_34693_, _34682_, _34181_);
  not (_34704_, _34693_);
  or (_34715_, _34704_, _27869_);
  not (_34725_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_34736_, _27869_, _34725_);
  and (_34747_, _34736_, _30651_);
  and (_34758_, _34747_, _34715_);
  nor (_34769_, _30640_, _34725_);
  not (_34780_, _27858_);
  and (_34791_, _26992_, _31286_);
  nor (_34802_, _26992_, _31286_);
  nor (_34813_, _34802_, _34791_);
  or (_34824_, _34813_, _34780_);
  and (_34834_, _34824_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_34845_, _34791_, _31885_);
  and (_34856_, _34802_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_34867_, _34856_, _34845_);
  and (_34878_, _34867_, _27858_);
  or (_34889_, _34878_, _34834_);
  and (_34900_, _34889_, _31351_);
  or (_34911_, _34900_, _34769_);
  or (_34922_, _34911_, _34758_);
  and (_08949_, _34922_, _43100_);
  and (_34942_, _26369_, _23628_);
  not (_34953_, _34942_);
  and (_34964_, _23532_, _18267_);
  nor (_34975_, _28231_, _28089_);
  nor (_34986_, _34975_, _29251_);
  nor (_34997_, _34986_, _29492_);
  nor (_35008_, _34997_, _29503_);
  and (_35019_, _35008_, _29613_);
  not (_35030_, _35019_);
  nor (_35041_, _29130_, _28220_);
  nor (_35051_, _35041_, _29141_);
  nor (_35062_, _35051_, _27946_);
  nor (_35073_, _29010_, _19807_);
  and (_35084_, _29010_, _20532_);
  nor (_35095_, _35084_, _35073_);
  nor (_35106_, _35095_, _29951_);
  and (_35117_, _29711_, _29010_);
  and (_35128_, _29809_, _29755_);
  nor (_35139_, _35128_, _35117_);
  nor (_35150_, _35139_, _20521_);
  and (_35160_, _35139_, _20521_);
  or (_35171_, _35160_, _32799_);
  nor (_35182_, _35171_, _35150_);
  nor (_35193_, _35182_, _35106_);
  not (_35204_, _30083_);
  and (_35215_, _35204_, _30039_);
  nor (_35226_, _30083_, _30028_);
  nor (_35237_, _35226_, _20521_);
  nor (_35248_, _35237_, _35215_);
  nor (_35259_, _35248_, _30814_);
  and (_35269_, _30246_, _28089_);
  nor (_35280_, _30225_, _28078_);
  not (_35291_, _35280_);
  and (_35302_, _30279_, _28067_);
  and (_35313_, _30301_, _20521_);
  nor (_35324_, _35313_, _35302_);
  nand (_35335_, _35324_, _35291_);
  nor (_35346_, _35335_, _35269_);
  nor (_35356_, _30388_, _20521_);
  not (_35367_, _35356_);
  nor (_35378_, _31568_, _19481_);
  nor (_35389_, _30345_, _20695_);
  nor (_35400_, _35389_, _35378_);
  and (_35411_, _35400_, _35367_);
  and (_35422_, _35411_, _35346_);
  not (_35433_, _35422_);
  nor (_35444_, _35433_, _35259_);
  and (_35455_, _35444_, _35193_);
  not (_35465_, _35455_);
  nor (_35476_, _35465_, _35062_);
  and (_35487_, _35476_, _35030_);
  not (_35498_, _35487_);
  nor (_35509_, _35498_, _34964_);
  and (_35520_, _35509_, _34953_);
  not (_35531_, _35520_);
  or (_35542_, _35531_, _27869_);
  not (_35553_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_35564_, _27869_, _35553_);
  and (_35575_, _35564_, _30651_);
  and (_35585_, _35575_, _35542_);
  nor (_35596_, _30640_, _35553_);
  and (_35607_, _32593_, _31286_);
  and (_35618_, _35607_, _27858_);
  nand (_35629_, _35618_, _31265_);
  or (_35640_, _35618_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_35651_, _35640_, _31351_);
  and (_35662_, _35651_, _35629_);
  or (_35673_, _35662_, _35596_);
  or (_35684_, _35673_, _35585_);
  and (_08960_, _35684_, _43100_);
  and (_35704_, _26433_, _23628_);
  not (_35715_, _35704_);
  and (_35726_, _23564_, _18267_);
  nor (_35737_, _29141_, _28187_);
  nor (_35748_, _35737_, _29152_);
  nor (_35759_, _35748_, _27946_);
  not (_35770_, _35759_);
  nor (_35781_, _29535_, _29503_);
  not (_35792_, _35781_);
  nor (_35803_, _29624_, _29536_);
  and (_35814_, _35803_, _35792_);
  nor (_35825_, _29010_, _27990_);
  or (_35835_, _35825_, _29951_);
  nor (_35846_, _35835_, _30781_);
  or (_35857_, _29010_, _20521_);
  or (_35868_, _35128_, _29722_);
  and (_35879_, _35868_, _35857_);
  nor (_35890_, _35879_, _19492_);
  and (_35901_, _35879_, _19492_);
  or (_35912_, _35901_, _32799_);
  nor (_35923_, _35912_, _35890_);
  nor (_35934_, _35923_, _35846_);
  nor (_35945_, _35215_, _19481_);
  and (_35955_, _35215_, _19481_);
  nor (_35966_, _35955_, _35945_);
  nor (_35977_, _35966_, _30814_);
  and (_35988_, _30246_, _28034_);
  nor (_35999_, _30225_, _28023_);
  not (_36010_, _35999_);
  and (_36021_, _30279_, _28012_);
  and (_36032_, _30301_, _19481_);
  nor (_36043_, _36032_, _36021_);
  nand (_36054_, _36043_, _36010_);
  nor (_36065_, _36054_, _35988_);
  nor (_36076_, _31568_, _20325_);
  not (_36086_, _36076_);
  nor (_36097_, _30388_, _19481_);
  nor (_36108_, _30345_, _20521_);
  nor (_36119_, _36108_, _36097_);
  and (_36130_, _36119_, _36086_);
  and (_36141_, _36130_, _36065_);
  not (_36152_, _36141_);
  nor (_36162_, _36152_, _35977_);
  and (_36173_, _36162_, _35934_);
  not (_36184_, _36173_);
  nor (_36195_, _36184_, _35814_);
  and (_36206_, _36195_, _35770_);
  not (_36217_, _36206_);
  nor (_36228_, _36217_, _35726_);
  and (_36239_, _36228_, _35715_);
  not (_36249_, _36239_);
  or (_36260_, _36249_, _27869_);
  not (_36271_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_36282_, _27869_, _36271_);
  and (_36293_, _36282_, _30651_);
  and (_36304_, _36293_, _36260_);
  nor (_36315_, _30640_, _36271_);
  nor (_36326_, _26740_, _26860_);
  and (_36336_, _36326_, _26981_);
  and (_36347_, _36336_, _27858_);
  nand (_36358_, _36347_, _31265_);
  or (_36369_, _36347_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_36380_, _36369_, _31351_);
  and (_36391_, _36380_, _36358_);
  or (_36402_, _36391_, _36315_);
  or (_36413_, _36402_, _36304_);
  and (_08971_, _36413_, _43100_);
  and (_36433_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36444_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_36455_, _36444_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_36466_, _36455_);
  not (_36477_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_36488_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_36498_, _36488_, _36477_);
  and (_36509_, _36444_, _18201_);
  and (_36520_, _36509_, _36498_);
  not (_36531_, _36520_);
  not (_36542_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_36553_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_36564_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_36575_, _36564_, _36553_);
  and (_36585_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_36596_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_36607_, _36596_, _36553_);
  and (_36618_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not (_36629_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_36640_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _36629_);
  and (_36651_, _36640_, _36553_);
  and (_36662_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_36672_, _36662_, _36618_);
  or (_36683_, _36672_, _36585_);
  and (_36694_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_36705_, _36596_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_36716_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_36727_, _36716_, _36694_);
  nor (_36738_, _36596_, _36553_);
  and (_36749_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  not (_36760_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_36770_, _36760_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_36781_, _36770_, _36553_);
  and (_36792_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_36803_, _36792_, _36749_);
  or (_36814_, _36803_, _36727_);
  nor (_36825_, _36814_, _36683_);
  and (_36836_, _36825_, _36542_);
  nor (_36847_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _36542_);
  or (_36858_, _36847_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_36869_, _36858_, _36836_);
  and (_36880_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_36890_, _36880_, _36869_);
  nor (_36901_, _36890_, _36531_);
  not (_36912_, _36901_);
  not (_36923_, _36498_);
  nor (_36934_, _36509_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_36945_, _36934_, _36923_);
  and (_36956_, _36945_, _36912_);
  not (_36967_, _36956_);
  and (_36978_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_36989_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37000_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_37011_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_37022_, _37011_, _37000_);
  and (_37033_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_37044_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_37055_, _37044_, _37033_);
  and (_37066_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_37077_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_37088_, _37077_, _37066_);
  and (_37099_, _37088_, _37055_);
  and (_37110_, _37099_, _37022_);
  nor (_37121_, _37110_, _36694_);
  and (_37132_, _37121_, _36542_);
  nor (_37142_, _37132_, _36989_);
  nor (_37153_, _37142_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37164_, _37153_, _36978_);
  and (_37175_, _37164_, _36520_);
  not (_37186_, _37175_);
  nor (_37197_, _36509_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_37208_, _37197_, _36923_);
  and (_37219_, _37208_, _37186_);
  and (_37230_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  not (_37241_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37251_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  or (_37262_, _36694_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37273_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_37284_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_37295_, _37284_, _37273_);
  and (_37306_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_37317_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_37328_, _37317_, _37306_);
  and (_37339_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_37350_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_37361_, _37350_, _37339_);
  and (_37371_, _37361_, _37328_);
  and (_37382_, _37371_, _37295_);
  nor (_37393_, _37382_, _37262_);
  or (_37404_, _37393_, _37251_);
  and (_37415_, _37404_, _37241_);
  nor (_37426_, _37415_, _37230_);
  nor (_37437_, _37426_, _36531_);
  and (_37448_, _36531_, \oc8051_top_1.oc8051_decoder1.op [7]);
  or (_37459_, _37448_, _37437_);
  and (_37470_, _37459_, _36498_);
  and (_37480_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37491_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37502_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_37513_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_37524_, _37513_, _37502_);
  and (_37535_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_37546_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_37557_, _37546_, _37535_);
  and (_37568_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_37579_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_37590_, _37579_, _37568_);
  and (_37601_, _37590_, _37557_);
  and (_37612_, _37601_, _37524_);
  nor (_37623_, _37612_, _37262_);
  or (_37634_, _37623_, _37491_);
  and (_37645_, _37634_, _37241_);
  nor (_37654_, _37645_, _37480_);
  and (_37665_, _37654_, _36520_);
  not (_37676_, _37665_);
  nor (_37687_, _36509_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_37698_, _37687_, _36923_);
  and (_37709_, _37698_, _37676_);
  not (_37720_, _37709_);
  and (_37731_, _37720_, _37470_);
  and (_37742_, _37731_, _37219_);
  and (_37753_, _37742_, _36967_);
  and (_37764_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37775_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37786_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_37797_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_37808_, _37797_, _37786_);
  and (_37819_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_37830_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_37841_, _37830_, _37819_);
  and (_37852_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_37863_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_37874_, _37863_, _37852_);
  and (_37885_, _37874_, _37841_);
  and (_37896_, _37885_, _37808_);
  nor (_37907_, _37896_, _36694_);
  and (_37918_, _37907_, _36542_);
  nor (_37929_, _37918_, _37775_);
  nor (_37940_, _37929_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37951_, _37940_, _37764_);
  and (_37962_, _37951_, _36520_);
  not (_37973_, _37962_);
  nor (_37984_, _36509_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_37995_, _37984_, _36923_);
  and (_38006_, _37995_, _37973_);
  not (_38017_, _36694_);
  and (_38028_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_38039_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_38050_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_38061_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_38072_, _38061_, _38050_);
  and (_38083_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_38094_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_38105_, _38094_, _38083_);
  nand (_38116_, _38105_, _38072_);
  or (_38127_, _38116_, _38039_);
  nor (_38138_, _38127_, _38028_);
  and (_38149_, _38138_, _38017_);
  and (_38160_, _38149_, _36542_);
  nor (_38171_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _36542_);
  nor (_38182_, _38171_, _38160_);
  nor (_38193_, _38182_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_38204_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _37241_);
  nor (_38215_, _38204_, _38193_);
  nor (_38226_, _38215_, _36531_);
  not (_38237_, _38226_);
  nor (_38248_, _36509_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_38259_, _38248_, _36923_);
  and (_38270_, _38259_, _38237_);
  and (_38281_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_38292_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_38302_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_38313_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_38324_, _38313_, _38302_);
  and (_38335_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_38345_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_38356_, _38345_, _38335_);
  and (_38367_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_38378_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_38389_, _38378_, _38367_);
  and (_38400_, _38389_, _38356_);
  and (_38406_, _38400_, _38324_);
  nor (_38407_, _38406_, _37262_);
  nor (_38408_, _38407_, _38292_);
  nor (_38409_, _38408_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_38410_, _38409_, _38281_);
  nor (_38411_, _38410_, _36531_);
  and (_38412_, _36531_, \oc8051_top_1.oc8051_decoder1.op [2]);
  or (_38413_, _38412_, _38411_);
  and (_38414_, _38413_, _36498_);
  and (_38415_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_38416_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_38417_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_38418_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_38419_, _38418_, _38417_);
  and (_38420_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_38421_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_38422_, _38421_, _38420_);
  and (_38423_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_38424_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_38425_, _38424_, _38423_);
  and (_38426_, _38425_, _38422_);
  and (_38427_, _38426_, _38419_);
  nor (_38428_, _38427_, _36694_);
  and (_38429_, _38428_, _36542_);
  or (_38430_, _38429_, _38416_);
  and (_38431_, _38430_, _37241_);
  nor (_38432_, _38431_, _38415_);
  and (_38433_, _38432_, _36520_);
  not (_38434_, _38433_);
  nor (_38435_, _36509_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_38436_, _38435_, _36923_);
  and (_38437_, _38436_, _38434_);
  nor (_38438_, _38437_, _38414_);
  and (_38439_, _38438_, _38270_);
  and (_38440_, _38439_, _38006_);
  and (_38441_, _38440_, _37753_);
  not (_38442_, _38441_);
  nor (_38443_, _37720_, _37470_);
  and (_38444_, _38443_, _37219_);
  and (_38445_, _38444_, _36956_);
  and (_38446_, _38440_, _38445_);
  nor (_38447_, _37219_, _37709_);
  and (_38448_, _38447_, _37470_);
  and (_38449_, _38448_, _36956_);
  and (_38450_, _38440_, _38449_);
  nor (_38451_, _38450_, _38446_);
  and (_38452_, _38451_, _38442_);
  and (_38453_, _38448_, _36967_);
  not (_38454_, _38437_);
  and (_38455_, _38454_, _38414_);
  nor (_38456_, _38006_, _38270_);
  and (_38457_, _38456_, _38455_);
  and (_38458_, _38457_, _38453_);
  and (_38459_, _38457_, _37753_);
  nor (_38460_, _38459_, _38458_);
  and (_38461_, _38460_, _38452_);
  nor (_38462_, _38461_, _36466_);
  not (_38463_, _38462_);
  not (_38464_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_38465_, _18201_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_38466_, _38465_, _38464_);
  and (_38467_, _38456_, _38438_);
  and (_38468_, _38467_, _38443_);
  and (_38469_, _38468_, _38466_);
  and (_38470_, _38459_, _18201_);
  and (_38471_, _38458_, _18201_);
  nor (_38472_, _38471_, _38470_);
  nor (_38473_, _38472_, _36444_);
  nor (_38474_, _38473_, _38469_);
  and (_38475_, _38474_, _38463_);
  nor (_38476_, _38475_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38477_, _38476_, _36433_);
  and (_38478_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_38479_, _38006_);
  nor (_38480_, _38479_, _38270_);
  and (_38481_, _38480_, _38455_);
  and (_38482_, _37709_, _37470_);
  and (_38483_, _38482_, _37219_);
  and (_38484_, _38483_, _36967_);
  and (_38485_, _38484_, _38481_);
  not (_38486_, _38485_);
  and (_38487_, _38270_, _38455_);
  and (_38488_, _38487_, _36967_);
  and (_38489_, _38488_, _37742_);
  not (_38490_, _38481_);
  and (_38491_, _37742_, _36956_);
  nor (_38492_, _38491_, _38449_);
  nor (_38493_, _38492_, _38490_);
  nor (_38494_, _38493_, _38489_);
  and (_38495_, _38494_, _38486_);
  nor (_38496_, _37709_, _37470_);
  and (_38497_, _38496_, _37219_);
  not (_38498_, _37219_);
  and (_38499_, _38443_, _38498_);
  and (_38500_, _38499_, _36956_);
  nor (_38501_, _38500_, _38497_);
  nor (_38502_, _38501_, _38490_);
  not (_38503_, _38502_);
  and (_38504_, _38439_, _38479_);
  and (_38505_, _38504_, _38497_);
  not (_38506_, _38505_);
  and (_38507_, _38496_, _38498_);
  and (_38508_, _38507_, _36967_);
  and (_38509_, _38508_, _38481_);
  and (_38510_, _37753_, _38437_);
  nor (_38511_, _38510_, _38509_);
  and (_38512_, _38511_, _38506_);
  and (_38513_, _38512_, _38503_);
  and (_38514_, _38444_, _36967_);
  and (_38515_, _38514_, _38481_);
  and (_38516_, _38482_, _38498_);
  and (_38517_, _38516_, _36967_);
  and (_38518_, _38517_, _38481_);
  nor (_38519_, _38518_, _38515_);
  and (_38520_, _38516_, _36956_);
  and (_38521_, _38520_, _38504_);
  and (_38522_, _37753_, _38504_);
  nor (_38523_, _38522_, _38521_);
  and (_38524_, _38523_, _38519_);
  and (_38525_, _38524_, _38513_);
  and (_38526_, _38525_, _38495_);
  and (_38527_, _38499_, _36967_);
  and (_38528_, _38527_, _38439_);
  not (_38529_, _38528_);
  and (_38530_, _38507_, _36956_);
  and (_38531_, _38530_, _38481_);
  and (_38532_, _38467_, _38491_);
  nor (_38533_, _38532_, _38531_);
  and (_38534_, _38533_, _38529_);
  and (_38535_, _38445_, _38504_);
  and (_38536_, _38520_, _38481_);
  nor (_38537_, _38536_, _38535_);
  and (_38538_, _38537_, _38534_);
  and (_38539_, _38467_, _37753_);
  and (_38540_, _38527_, _38481_);
  nor (_38541_, _38540_, _38539_);
  and (_38542_, _38504_, _38491_);
  and (_38543_, _38517_, _38504_);
  nor (_38544_, _38543_, _38542_);
  and (_38545_, _38544_, _38541_);
  and (_38546_, _38545_, _38538_);
  and (_38547_, _38453_, _38504_);
  and (_38548_, _38439_, _38500_);
  nor (_38549_, _38548_, _38547_);
  and (_38550_, _38504_, _38449_);
  and (_38551_, _38453_, _38481_);
  nor (_38552_, _38551_, _38550_);
  and (_38553_, _38552_, _38549_);
  and (_38554_, _38497_, _36956_);
  and (_38555_, _38554_, _38467_);
  not (_38556_, _38555_);
  and (_38557_, _38497_, _36967_);
  and (_38558_, _38557_, _38467_);
  and (_38559_, _38467_, _38530_);
  nor (_38560_, _38559_, _38558_);
  and (_38561_, _38560_, _38556_);
  and (_38562_, _38467_, _38516_);
  and (_38563_, _38514_, _38439_);
  nor (_38564_, _38563_, _38562_);
  and (_38565_, _38564_, _38561_);
  and (_38566_, _38565_, _38553_);
  and (_38567_, _38566_, _38546_);
  and (_38568_, _38567_, _38526_);
  nor (_38569_, _38568_, _36466_);
  and (_38570_, \oc8051_top_1.oc8051_decoder1.state [0], _18201_);
  and (_38571_, _38570_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_38572_, _38571_, _38505_);
  nor (_38573_, _38572_, _38469_);
  not (_38574_, _38573_);
  nor (_38575_, _38574_, _38569_);
  nor (_38576_, _38575_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38577_, _38576_, _38478_);
  and (_38578_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_38579_, _38270_, _38414_);
  nor (_38580_, _36967_, _38437_);
  and (_38581_, _38580_, _38579_);
  and (_38582_, _38581_, _38499_);
  and (_38583_, _38497_, _38487_);
  or (_38584_, _38583_, _38582_);
  not (_38585_, _38584_);
  and (_38586_, _38453_, _38487_);
  nor (_38587_, _38586_, _38505_);
  and (_38588_, _38581_, _37742_);
  and (_38589_, _38507_, _38487_);
  nor (_38590_, _38589_, _38588_);
  not (_38591_, _38590_);
  or (_38592_, _38499_, _38483_);
  and (_38593_, _38592_, _38488_);
  nor (_38594_, _38593_, _38591_);
  and (_38595_, _38594_, _38587_);
  and (_38596_, _38595_, _38585_);
  and (_38597_, _38562_, _36956_);
  not (_38598_, _38597_);
  and (_38599_, _38516_, _38487_);
  and (_38600_, _38581_, _38448_);
  nor (_38601_, _38600_, _38599_);
  not (_38602_, _38601_);
  and (_38603_, _38514_, _38487_);
  nor (_38604_, _38603_, _38602_);
  and (_38605_, _38604_, _38598_);
  and (_38606_, _38605_, _38452_);
  and (_38607_, _38606_, _38596_);
  nor (_38608_, _38607_, _36466_);
  and (_38609_, _38466_, _38444_);
  and (_38610_, _38609_, _38467_);
  or (_38611_, _38610_, _38572_);
  nor (_38612_, _38611_, _38608_);
  nor (_38613_, _38612_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38614_, _38613_, _38578_);
  nor (_38615_, _38614_, _38577_);
  and (_38616_, _38615_, _38477_);
  and (_09521_, _38616_, _43100_);
  and (_38617_, _30651_, _27650_);
  and (_38618_, _27825_, _27343_);
  and (_38619_, _27211_, _27507_);
  and (_38620_, _38619_, _38618_);
  and (_38621_, _38620_, _32593_);
  and (_38622_, _38621_, _26740_);
  and (_38623_, _38622_, _38617_);
  not (_38624_, _38623_);
  and (_38625_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_38626_, _23628_, _18267_);
  and (_38627_, _29602_, _23606_);
  nor (_38628_, _30377_, _38627_);
  and (_38629_, _38628_, _30345_);
  and (_38630_, _38629_, _38626_);
  and (_38631_, _38630_, _31568_);
  nor (_38632_, _38631_, _19481_);
  not (_38633_, _38632_);
  and (_38634_, _38633_, _36065_);
  and (_38635_, _38634_, _35934_);
  nor (_38636_, _38635_, _38624_);
  nor (_38637_, _38636_, _38625_);
  and (_38638_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_38639_, _38631_, _20521_);
  not (_38640_, _38639_);
  and (_38641_, _38640_, _35346_);
  and (_38642_, _38641_, _35193_);
  nor (_38643_, _38642_, _38624_);
  nor (_38644_, _38643_, _38638_);
  and (_38645_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_38646_, _38631_, _20695_);
  not (_38647_, _38646_);
  and (_38648_, _38647_, _34366_);
  and (_38649_, _38648_, _34475_);
  and (_38650_, _38649_, _34333_);
  nor (_38651_, _38650_, _38624_);
  nor (_38652_, _38651_, _38645_);
  and (_38653_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_38654_, _38631_, _21054_);
  not (_38655_, _38654_);
  and (_38656_, _38655_, _33637_);
  and (_38657_, _38656_, _33605_);
  and (_38658_, _38657_, _33921_);
  nor (_38659_, _38658_, _38624_);
  nor (_38660_, _38659_, _38653_);
  and (_38661_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_38662_, _38631_, _21555_);
  not (_38663_, _38662_);
  and (_38664_, _38663_, _32963_);
  and (_38665_, _38664_, _32843_);
  nor (_38666_, _38665_, _38624_);
  nor (_38667_, _38666_, _38661_);
  and (_38668_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_38669_, _38631_, _21381_);
  not (_38670_, _38669_);
  and (_38671_, _38670_, _32244_);
  and (_38672_, _38671_, _32440_);
  nor (_38673_, _38672_, _38624_);
  nor (_38674_, _38673_, _38668_);
  and (_38675_, _38617_, _26740_);
  and (_38676_, _38675_, _38621_);
  nor (_38677_, _38676_, _26926_);
  nor (_38678_, _38631_, _21925_);
  not (_38679_, _38678_);
  and (_38680_, _38679_, _31656_);
  and (_38681_, _38680_, _31634_);
  and (_38682_, _38681_, _31546_);
  not (_38683_, _38682_);
  and (_38684_, _38683_, _38623_);
  nor (_38685_, _38684_, _38677_);
  and (_38686_, _38685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38687_, _38686_, _38674_);
  and (_38688_, _38687_, _38667_);
  and (_38689_, _38688_, _38660_);
  and (_38690_, _38689_, _38652_);
  and (_38691_, _38690_, _38644_);
  and (_38692_, _38691_, _38637_);
  nor (_38693_, _38676_, _27365_);
  nand (_38694_, _38693_, _38692_);
  or (_38695_, _38693_, _38692_);
  and (_38696_, _38695_, _27069_);
  and (_38697_, _38696_, _38694_);
  or (_38698_, _38676_, _27409_);
  or (_38699_, _38698_, _38697_);
  nor (_38700_, _38631_, _20325_);
  not (_38701_, _38700_);
  and (_38702_, _38701_, _30323_);
  and (_38703_, _38702_, _30268_);
  and (_38704_, _38703_, _29984_);
  nand (_38705_, _38704_, _38676_);
  and (_38706_, _38705_, _38699_);
  and (_09542_, _38706_, _43100_);
  not (_38707_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38708_, _38685_, _38707_);
  nor (_38709_, _38685_, _38707_);
  nor (_38710_, _38709_, _38708_);
  and (_38711_, _38710_, _27069_);
  nor (_38712_, _38711_, _26937_);
  nor (_38713_, _38712_, _38623_);
  nor (_38714_, _38713_, _38684_);
  nand (_10698_, _38714_, _43100_);
  nor (_38715_, _38686_, _38674_);
  nor (_38716_, _38715_, _38687_);
  nor (_38717_, _38716_, _26487_);
  nor (_38718_, _38717_, _26784_);
  nor (_38719_, _38718_, _38623_);
  nor (_38720_, _38719_, _38673_);
  nand (_10709_, _38720_, _43100_);
  nor (_38721_, _38687_, _38667_);
  nor (_38722_, _38721_, _38688_);
  nor (_38723_, _38722_, _26487_);
  nor (_38724_, _38723_, _26542_);
  nor (_38725_, _38724_, _38623_);
  nor (_38726_, _38725_, _38666_);
  nand (_10720_, _38726_, _43100_);
  nor (_38727_, _38688_, _38660_);
  nor (_38728_, _38727_, _38689_);
  nor (_38729_, _38728_, _26487_);
  nor (_38730_, _38729_, _27584_);
  nor (_38731_, _38730_, _38623_);
  nor (_38732_, _38731_, _38659_);
  nor (_10731_, _38732_, rst);
  nor (_38733_, _38689_, _38652_);
  nor (_38734_, _38733_, _38690_);
  nor (_38735_, _38734_, _26487_);
  nor (_38736_, _38735_, _27760_);
  nor (_38737_, _38736_, _38623_);
  nor (_38738_, _38737_, _38651_);
  nor (_10742_, _38738_, rst);
  nor (_38739_, _38690_, _38644_);
  nor (_38740_, _38739_, _38691_);
  nor (_38741_, _38740_, _26487_);
  nor (_38742_, _38741_, _27255_);
  nor (_38743_, _38742_, _38623_);
  nor (_38744_, _38743_, _38643_);
  nor (_10753_, _38744_, rst);
  nor (_38745_, _38691_, _38637_);
  nor (_38746_, _38745_, _38692_);
  nor (_38747_, _38746_, _26487_);
  nor (_38748_, _38747_, _27102_);
  nor (_38749_, _38748_, _38623_);
  nor (_38750_, _38749_, _38636_);
  nor (_10764_, _38750_, rst);
  and (_38751_, _38620_, _34052_);
  nand (_38752_, _38751_, _38617_);
  nor (_38753_, _38752_, _30574_);
  and (_38754_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18201_);
  and (_38755_, _38754_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38756_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38757_, _38756_, _38755_);
  or (_38758_, _38757_, _38753_);
  nor (_38759_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38760_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38761_, _38760_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38762_, _38761_, _38759_);
  nor (_38763_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38764_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38765_, _38764_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38766_, _38765_, _38763_);
  nor (_38767_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38768_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38769_, _38768_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38770_, _38769_, _38767_);
  nor (_38771_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38772_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38773_, _38772_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38774_, _38773_, _38771_);
  nor (_38775_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38776_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38777_, _38776_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38778_, _38777_, _38775_);
  not (_38779_, _38778_);
  nor (_38780_, _38779_, _30716_);
  nor (_38781_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38782_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38783_, _38782_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38784_, _38783_, _38781_);
  and (_38785_, _38784_, _38780_);
  nor (_38786_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38787_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38788_, _38787_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38789_, _38788_, _38786_);
  and (_38790_, _38789_, _38785_);
  and (_38791_, _38790_, _38774_);
  nor (_38792_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38793_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38794_, _38793_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38795_, _38794_, _38792_);
  and (_38796_, _38795_, _38791_);
  and (_38797_, _38796_, _38770_);
  and (_38798_, _38797_, _38766_);
  or (_38799_, _38798_, _38762_);
  nand (_38800_, _38798_, _38762_);
  and (_38801_, _38800_, _38799_);
  and (_38802_, _38801_, _29613_);
  not (_38803_, _38802_);
  and (_38804_, _23320_, _18267_);
  and (_38805_, _29733_, _20336_);
  and (_38806_, _38805_, _28374_);
  and (_38807_, _38806_, _28407_);
  and (_38808_, _38807_, _28450_);
  and (_38809_, _38808_, _29064_);
  nor (_38810_, _38809_, _29755_);
  and (_38811_, _29010_, _18836_);
  nor (_38812_, _38811_, _38810_);
  and (_38813_, _29820_, _20325_);
  and (_38814_, _19655_, _18671_);
  and (_38815_, _19977_, _18990_);
  and (_38816_, _38815_, _38814_);
  and (_38817_, _38816_, _38813_);
  and (_38818_, _19807_, _18836_);
  and (_38819_, _38818_, _38817_);
  nor (_38820_, _38819_, _29010_);
  and (_38821_, _29010_, _19807_);
  nor (_38822_, _38821_, _38820_);
  and (_38823_, _38822_, _38812_);
  nor (_38824_, _29010_, _19166_);
  and (_38825_, _29010_, _19166_);
  nor (_38826_, _38825_, _38824_);
  and (_38827_, _38826_, _38823_);
  and (_38828_, _38827_, _29897_);
  nor (_38829_, _38827_, _29897_);
  nor (_38830_, _38829_, _38828_);
  and (_38831_, _38830_, _29668_);
  and (_38832_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_38833_, _29010_, _29897_);
  nor (_38834_, _38833_, _30825_);
  nor (_38835_, _38834_, _29951_);
  nor (_38836_, _31141_, _21054_);
  nor (_38837_, _30388_, _20151_);
  or (_38838_, _38837_, _38836_);
  or (_38839_, _38838_, _38835_);
  nor (_38840_, _38839_, _38832_);
  not (_38841_, _38840_);
  nor (_38842_, _38841_, _38831_);
  not (_38843_, _38842_);
  nor (_38844_, _38843_, _38804_);
  and (_38845_, _38844_, _38803_);
  nand (_38846_, _38845_, _38755_);
  and (_38847_, _38846_, _43100_);
  and (_12715_, _38847_, _38758_);
  and (_38848_, _38620_, _33344_);
  and (_38849_, _38848_, _38617_);
  nor (_38850_, _38849_, _38755_);
  not (_38851_, _38850_);
  nand (_38852_, _38851_, _30574_);
  or (_38853_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38854_, _38853_, _43100_);
  and (_12736_, _38854_, _38852_);
  nor (_38855_, _38752_, _31808_);
  and (_38856_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38857_, _38856_, _38755_);
  or (_38858_, _38857_, _38855_);
  and (_38859_, _25897_, _23628_);
  not (_38860_, _38859_);
  and (_38861_, _38779_, _30716_);
  nor (_38862_, _38861_, _38780_);
  and (_38863_, _38862_, _29613_);
  nor (_38864_, _30825_, _29930_);
  not (_38865_, _38864_);
  nor (_38866_, _38865_, _29842_);
  nor (_38867_, _38866_, _28374_);
  and (_38868_, _38866_, _28374_);
  or (_38869_, _38868_, _32799_);
  nor (_38870_, _38869_, _38867_);
  nor (_38871_, _30388_, _18990_);
  and (_38872_, _23098_, _18267_);
  nor (_38873_, _31141_, _20695_);
  nor (_38874_, _29951_, _21925_);
  or (_38875_, _38874_, _38873_);
  or (_38876_, _38875_, _38872_);
  nor (_38877_, _38876_, _38871_);
  not (_38878_, _38877_);
  nor (_38879_, _38878_, _38870_);
  not (_38880_, _38879_);
  nor (_38881_, _38880_, _38863_);
  and (_38882_, _38881_, _38860_);
  nand (_38883_, _38882_, _38755_);
  and (_38884_, _38883_, _43100_);
  and (_13649_, _38884_, _38858_);
  nor (_38885_, _38752_, _32495_);
  and (_38886_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38887_, _38886_, _38755_);
  or (_38888_, _38887_, _38885_);
  nor (_38889_, _38784_, _38780_);
  not (_38890_, _38889_);
  nor (_38891_, _38785_, _29624_);
  and (_38892_, _38891_, _38890_);
  not (_38893_, _38892_);
  and (_38894_, _24911_, _23628_);
  nor (_38895_, _20325_, _18990_);
  and (_38896_, _38895_, _29733_);
  and (_38897_, _38896_, _29010_);
  and (_38898_, _38813_, _18990_);
  and (_38899_, _38898_, _29755_);
  nor (_38900_, _38899_, _38897_);
  nor (_38901_, _38900_, _28407_);
  and (_38902_, _38900_, _28407_);
  nor (_38903_, _38902_, _38901_);
  nor (_38904_, _38903_, _32799_);
  nor (_38905_, _30388_, _19977_);
  and (_38906_, _23130_, _18267_);
  nor (_38907_, _31141_, _20521_);
  nor (_38908_, _29951_, _21381_);
  or (_38909_, _38908_, _38907_);
  or (_38910_, _38909_, _38906_);
  nor (_38911_, _38910_, _38905_);
  not (_38912_, _38911_);
  nor (_38913_, _38912_, _38904_);
  not (_38914_, _38913_);
  nor (_38915_, _38914_, _38894_);
  and (_38916_, _38915_, _38893_);
  nand (_38917_, _38916_, _38755_);
  and (_38918_, _38917_, _43100_);
  and (_13660_, _38918_, _38888_);
  nor (_38919_, _38752_, _33202_);
  and (_38920_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38921_, _38920_, _38755_);
  or (_38922_, _38921_, _38919_);
  nor (_38923_, _38789_, _38785_);
  nor (_38924_, _38923_, _38790_);
  and (_38925_, _38924_, _29613_);
  not (_38926_, _38925_);
  and (_38927_, _38898_, _19977_);
  and (_38928_, _38927_, _29755_);
  and (_38929_, _38896_, _28407_);
  and (_38930_, _38929_, _29010_);
  nor (_38931_, _38930_, _38928_);
  and (_38932_, _38931_, _18671_);
  nor (_38933_, _38931_, _18671_);
  nor (_38934_, _38933_, _38932_);
  and (_38935_, _38934_, _29668_);
  not (_38936_, _38935_);
  nor (_38937_, _29951_, _21555_);
  and (_38938_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38939_, _38938_, _38937_);
  and (_38940_, _23162_, _18267_);
  nor (_38941_, _31141_, _19481_);
  nor (_38942_, _30388_, _18671_);
  or (_38943_, _38942_, _38941_);
  nor (_38944_, _38943_, _38940_);
  and (_38945_, _38944_, _38939_);
  and (_38946_, _38945_, _38936_);
  and (_38947_, _38946_, _38926_);
  nand (_38948_, _38947_, _38755_);
  and (_38949_, _38948_, _43100_);
  and (_13671_, _38949_, _38922_);
  nor (_38950_, _38752_, _33953_);
  and (_38951_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38952_, _38951_, _38755_);
  or (_38953_, _38952_, _38950_);
  nor (_38954_, _38790_, _38774_);
  nor (_38955_, _38954_, _38791_);
  and (_38956_, _38955_, _29613_);
  not (_38957_, _38956_);
  nor (_38958_, _38808_, _29064_);
  not (_38959_, _38958_);
  and (_38960_, _38959_, _38810_);
  and (_38961_, _38927_, _18671_);
  nor (_38962_, _38961_, _19655_);
  nor (_38963_, _38962_, _38817_);
  nor (_38964_, _38963_, _29010_);
  nor (_38965_, _38964_, _38960_);
  nor (_38966_, _38965_, _32799_);
  nor (_38967_, _30388_, _19655_);
  or (_38968_, _38967_, _31142_);
  nor (_38969_, _38968_, _38966_);
  and (_38970_, _23193_, _18267_);
  nor (_38971_, _29951_, _21054_);
  and (_38972_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_38973_, _38972_, _38971_);
  nor (_38974_, _38973_, _38970_);
  and (_38975_, _38974_, _38969_);
  and (_38976_, _38975_, _38957_);
  nand (_38977_, _38976_, _38755_);
  and (_38978_, _38977_, _43100_);
  and (_13682_, _38978_, _38953_);
  nor (_38979_, _38752_, _34693_);
  and (_38980_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_38981_, _38980_, _38755_);
  or (_38982_, _38981_, _38979_);
  nor (_38983_, _38795_, _38791_);
  nor (_38984_, _38983_, _38796_);
  and (_38985_, _38984_, _29613_);
  not (_38986_, _38985_);
  and (_38987_, _23225_, _18267_);
  nor (_38988_, _38817_, _29010_);
  nor (_38989_, _38988_, _38810_);
  nor (_38990_, _38989_, _28100_);
  and (_38991_, _38989_, _28100_);
  nor (_38992_, _38991_, _38990_);
  and (_38993_, _38992_, _29668_);
  and (_38994_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_38995_, _29010_, _20706_);
  or (_38996_, _38995_, _29951_);
  nor (_38997_, _38996_, _38811_);
  nor (_38998_, _31141_, _21925_);
  nor (_38999_, _30388_, _18836_);
  or (_39000_, _38999_, _38998_);
  or (_39001_, _39000_, _38997_);
  nor (_39002_, _39001_, _38994_);
  not (_39003_, _39002_);
  nor (_39004_, _39003_, _38993_);
  not (_39005_, _39004_);
  nor (_39006_, _39005_, _38987_);
  and (_39007_, _39006_, _38986_);
  nand (_39008_, _39007_, _38755_);
  and (_39009_, _39008_, _43100_);
  and (_13693_, _39009_, _38982_);
  nor (_39010_, _38752_, _35520_);
  and (_39011_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_39012_, _39011_, _38755_);
  or (_39013_, _39012_, _39010_);
  nor (_39014_, _38796_, _38770_);
  not (_39015_, _39014_);
  nor (_39016_, _38797_, _29624_);
  and (_39017_, _39016_, _39015_);
  not (_39018_, _39017_);
  and (_39019_, _23257_, _18267_);
  and (_39020_, _38817_, _18836_);
  nor (_39021_, _39020_, _29010_);
  not (_39022_, _39021_);
  and (_39023_, _39022_, _38812_);
  and (_39024_, _39023_, _19807_);
  nor (_39025_, _39023_, _19807_);
  nor (_39026_, _39025_, _39024_);
  nor (_39027_, _39026_, _32799_);
  and (_39028_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_39029_, _29010_, _20532_);
  or (_39030_, _39029_, _29951_);
  nor (_39031_, _39030_, _38821_);
  nor (_39032_, _31141_, _21381_);
  nor (_39033_, _30388_, _19807_);
  or (_39034_, _39033_, _39032_);
  or (_39035_, _39034_, _39031_);
  nor (_39036_, _39035_, _39028_);
  not (_39037_, _39036_);
  nor (_39038_, _39037_, _39027_);
  not (_39039_, _39038_);
  nor (_39040_, _39039_, _39019_);
  and (_39041_, _39040_, _39018_);
  nand (_39042_, _39041_, _38755_);
  and (_39043_, _39042_, _43100_);
  and (_13704_, _39043_, _39013_);
  nor (_39044_, _38752_, _36239_);
  and (_39045_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_39046_, _39045_, _38755_);
  or (_39047_, _39046_, _39044_);
  nor (_39048_, _38797_, _38766_);
  not (_39049_, _39048_);
  nor (_39050_, _38798_, _29624_);
  and (_39051_, _39050_, _39049_);
  not (_39052_, _39051_);
  and (_39053_, _23288_, _18267_);
  and (_39054_, _38823_, _19166_);
  nor (_39055_, _38823_, _19166_);
  nor (_39056_, _39055_, _39054_);
  nor (_39057_, _39056_, _32799_);
  and (_39058_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_39059_, _29010_, _19492_);
  or (_39060_, _39059_, _29951_);
  nor (_39061_, _39060_, _38825_);
  nor (_39062_, _31141_, _21555_);
  nor (_39063_, _30388_, _19166_);
  or (_39064_, _39063_, _39062_);
  or (_39065_, _39064_, _39061_);
  nor (_39066_, _39065_, _39058_);
  not (_39067_, _39066_);
  nor (_39068_, _39067_, _39057_);
  not (_39069_, _39068_);
  nor (_39070_, _39069_, _39053_);
  and (_39071_, _39070_, _39052_);
  nand (_39072_, _39071_, _38755_);
  and (_39073_, _39072_, _43100_);
  and (_13715_, _39073_, _39047_);
  nand (_39074_, _38851_, _31808_);
  or (_39075_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_39076_, _39075_, _43100_);
  and (_13726_, _39076_, _39074_);
  nand (_39077_, _38851_, _32495_);
  or (_39078_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_39079_, _39078_, _43100_);
  and (_13737_, _39079_, _39077_);
  nand (_39080_, _38851_, _33202_);
  or (_39081_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_39082_, _39081_, _43100_);
  and (_13748_, _39082_, _39080_);
  nand (_39083_, _38851_, _33953_);
  or (_39084_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_39085_, _39084_, _43100_);
  and (_13758_, _39085_, _39083_);
  nand (_39086_, _38851_, _34693_);
  or (_39087_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_39088_, _39087_, _43100_);
  and (_13769_, _39088_, _39086_);
  nand (_39089_, _38851_, _35520_);
  or (_39090_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_39091_, _39090_, _43100_);
  and (_13780_, _39091_, _39089_);
  nand (_39092_, _38851_, _36239_);
  or (_39093_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_39094_, _39093_, _43100_);
  and (_13791_, _39094_, _39092_);
  not (_39095_, _27343_);
  nor (_39096_, _39095_, _27211_);
  and (_39097_, _39096_, _31351_);
  and (_39098_, _39097_, _27847_);
  not (_39099_, _31308_);
  nor (_39100_, _39099_, _31265_);
  not (_39101_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_39102_, _31308_, _39101_);
  or (_39103_, _39102_, _39100_);
  and (_39104_, _39103_, _39098_);
  nor (_39105_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_39106_, _39105_);
  nand (_39107_, _39106_, _31265_);
  and (_39108_, _39105_, _39101_);
  nor (_39109_, _39108_, _39098_);
  and (_39110_, _39109_, _39107_);
  nor (_39111_, _27825_, _39095_);
  nor (_39112_, _27211_, _27496_);
  and (_39113_, _38617_, _27003_);
  and (_39114_, _39113_, _39112_);
  and (_39115_, _39114_, _39111_);
  or (_39116_, _39115_, _39110_);
  or (_39117_, _39116_, _39104_);
  nand (_39118_, _39115_, _38704_);
  and (_39119_, _39118_, _43100_);
  and (_15195_, _39119_, _39117_);
  and (_39120_, _39098_, _32604_);
  nand (_39121_, _39120_, _31265_);
  not (_39122_, _39115_);
  or (_39123_, _39120_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_39124_, _39123_, _39122_);
  and (_39125_, _39124_, _39121_);
  nor (_39126_, _39122_, _38672_);
  or (_39127_, _39126_, _39125_);
  and (_17376_, _39127_, _43100_);
  or (_39128_, _23384_, _23352_);
  or (_39129_, _39128_, _23415_);
  or (_39130_, _39129_, _23468_);
  or (_39131_, _39130_, _23490_);
  or (_39132_, _39131_, _23532_);
  and (_39133_, _39132_, _18267_);
  or (_39134_, _30759_, _29163_);
  not (_39135_, _30749_);
  nand (_39136_, _39135_, _29163_);
  and (_39137_, _39136_, _27935_);
  and (_39138_, _39137_, _39134_);
  not (_39139_, _27957_);
  nand (_39140_, _29558_, _39139_);
  or (_39141_, _29558_, _27978_);
  and (_39142_, _29613_, _39141_);
  and (_39143_, _39142_, _39140_);
  and (_39144_, _38818_, _24812_);
  and (_39145_, _38816_, _23628_);
  nand (_39146_, _39145_, _39144_);
  nand (_39147_, _39146_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_39148_, _39147_, _39143_);
  or (_39149_, _39148_, _39138_);
  or (_39150_, _39149_, _35726_);
  or (_39151_, _39150_, _39133_);
  or (_39152_, _39151_, _27902_);
  nor (_39153_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_39154_, _39153_, _39098_);
  and (_39155_, _39154_, _39152_);
  and (_39156_, _33355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_39157_, _39156_, _33366_);
  and (_39158_, _39157_, _39098_);
  or (_39159_, _39158_, _39115_);
  or (_39160_, _39159_, _39155_);
  nand (_39161_, _39115_, _38665_);
  and (_39162_, _39161_, _43100_);
  and (_17387_, _39162_, _39160_);
  and (_39163_, _39098_, _34052_);
  nand (_39164_, _39163_, _31265_);
  or (_39165_, _39163_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_39166_, _39165_, _39122_);
  and (_39167_, _39166_, _39164_);
  nor (_39168_, _39122_, _38658_);
  or (_39169_, _39168_, _39167_);
  and (_17398_, _39169_, _43100_);
  not (_39170_, _39098_);
  or (_39171_, _39170_, _34813_);
  and (_39172_, _39171_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_39175_, _34802_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_39177_, _39175_, _34845_);
  and (_39178_, _39177_, _39098_);
  or (_39179_, _39178_, _39172_);
  and (_39180_, _39179_, _39122_);
  nor (_39181_, _39122_, _38650_);
  or (_39182_, _39181_, _39180_);
  and (_17409_, _39182_, _43100_);
  and (_39183_, _39098_, _35607_);
  nand (_39184_, _39183_, _31265_);
  or (_39185_, _39183_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_39187_, _39185_, _39122_);
  and (_39196_, _39187_, _39184_);
  nor (_39202_, _39122_, _38642_);
  or (_39208_, _39202_, _39196_);
  and (_17420_, _39208_, _43100_);
  and (_39211_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_39212_, _39211_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_39213_, _29119_, _27935_);
  and (_39214_, _29613_, _29481_);
  nand (_39215_, _30377_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_39216_, _39215_, _39211_);
  or (_39217_, _39216_, _39214_);
  or (_39218_, _39217_, _39213_);
  and (_39219_, _39218_, _39212_);
  or (_39220_, _39219_, _39098_);
  not (_39221_, _36336_);
  nor (_39222_, _39221_, _31265_);
  or (_39223_, _36336_, _33496_);
  nand (_39224_, _39223_, _39098_);
  or (_39225_, _39224_, _39222_);
  and (_39226_, _39225_, _39220_);
  or (_39227_, _39226_, _39115_);
  nand (_39228_, _39115_, _38635_);
  and (_39229_, _39228_, _43100_);
  and (_17431_, _39229_, _39227_);
  not (_39230_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39231_, _38754_, _39230_);
  not (_39232_, _39231_);
  nor (_39233_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_39236_, _39233_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39237_, _27003_, _27650_);
  and (_39238_, _27825_, _39095_);
  and (_39239_, _39238_, _39112_);
  and (_39240_, _39239_, _39237_);
  and (_39241_, _39240_, _30651_);
  nor (_39242_, _39241_, _39236_);
  nor (_39243_, _39242_, _30574_);
  and (_39244_, _27825_, _27650_);
  and (_39245_, _39244_, _27354_);
  not (_39246_, _31351_);
  nor (_39247_, _39246_, _27496_);
  and (_39248_, _39247_, _39245_);
  and (_39249_, _39248_, _31308_);
  and (_39250_, _39249_, _31265_);
  nor (_39251_, _39249_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_39252_, _39251_);
  and (_39253_, _39242_, _39232_);
  and (_39254_, _39253_, _39252_);
  not (_39255_, _39254_);
  nor (_39256_, _39255_, _39250_);
  or (_39257_, _39256_, _39243_);
  and (_39258_, _39257_, _39232_);
  nor (_39259_, _39232_, _38845_);
  or (_39260_, _39259_, _39258_);
  and (_18000_, _39260_, _43100_);
  nor (_39261_, _39232_, _38882_);
  not (_39262_, _39242_);
  and (_39263_, _39262_, _31808_);
  not (_39264_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_39265_, _39248_, _39264_);
  nor (_39266_, _39265_, _39262_);
  not (_39267_, _39266_);
  and (_39268_, _31885_, _27003_);
  nor (_39269_, _27003_, _39264_);
  nor (_39270_, _39269_, _39268_);
  and (_39271_, _39244_, _27507_);
  and (_39272_, _31351_, _27354_);
  and (_39274_, _39272_, _39271_);
  and (_39278_, _39253_, _39274_);
  not (_39284_, _39278_);
  nor (_39289_, _39284_, _39270_);
  nor (_39296_, _39289_, _39267_);
  nor (_39304_, _39296_, _39231_);
  not (_39312_, _39304_);
  nor (_39313_, _39312_, _39263_);
  nor (_39314_, _39313_, _39261_);
  nor (_19851_, _39314_, rst);
  nor (_39315_, _39242_, _32495_);
  and (_39316_, _39248_, _32604_);
  and (_39317_, _39316_, _31265_);
  nor (_39318_, _39316_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not (_39319_, _39318_);
  and (_39320_, _39319_, _39253_);
  not (_39321_, _39320_);
  nor (_39322_, _39321_, _39317_);
  or (_39323_, _39322_, _39315_);
  and (_39324_, _39323_, _39232_);
  nor (_39325_, _39232_, _38916_);
  or (_39326_, _39325_, _39324_);
  and (_19863_, _39326_, _43100_);
  nor (_39327_, _39242_, _33202_);
  and (_39328_, _39248_, _33344_);
  and (_39329_, _39328_, _31265_);
  nor (_39330_, _39328_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_39331_, _39330_);
  and (_39332_, _39331_, _39253_);
  not (_39333_, _39332_);
  nor (_39334_, _39333_, _39329_);
  or (_39335_, _39334_, _39327_);
  and (_39336_, _39335_, _39232_);
  nor (_39337_, _39232_, _38947_);
  or (_39338_, _39337_, _39336_);
  and (_19875_, _39338_, _43100_);
  nor (_39339_, _39232_, _38976_);
  and (_39340_, _39262_, _33953_);
  not (_39341_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_39342_, _39248_, _39341_);
  not (_39343_, _39342_);
  not (_39344_, _39248_);
  nor (_39345_, _34052_, _39341_);
  nor (_39346_, _39345_, _34062_);
  or (_39352_, _39346_, _39344_);
  and (_39363_, _39352_, _39242_);
  and (_39364_, _39363_, _39343_);
  nor (_39365_, _39364_, _39231_);
  not (_39366_, _39365_);
  nor (_39377_, _39366_, _39340_);
  nor (_39383_, _39377_, _39339_);
  nor (_19886_, _39383_, rst);
  nor (_39384_, _39242_, _34693_);
  and (_39385_, _39248_, _34791_);
  and (_39386_, _39385_, _31265_);
  nor (_39387_, _39385_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_39388_, _39387_);
  and (_39389_, _39388_, _39253_);
  not (_39390_, _39389_);
  nor (_39391_, _39390_, _39386_);
  or (_39392_, _39391_, _39384_);
  and (_39393_, _39392_, _39232_);
  nor (_39394_, _39232_, _39007_);
  or (_39395_, _39394_, _39393_);
  and (_19898_, _39395_, _43100_);
  nor (_39396_, _39242_, _35520_);
  and (_39397_, _39248_, _35607_);
  and (_39398_, _39397_, _31265_);
  nor (_39399_, _39397_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not (_39400_, _39399_);
  and (_39401_, _39400_, _39253_);
  not (_39402_, _39401_);
  nor (_39403_, _39402_, _39398_);
  or (_39404_, _39403_, _39396_);
  and (_39405_, _39404_, _39232_);
  nor (_39406_, _39232_, _39041_);
  or (_39407_, _39406_, _39405_);
  and (_19910_, _39407_, _43100_);
  nor (_39408_, _39242_, _36239_);
  and (_39409_, _39253_, _39344_);
  and (_39410_, _39409_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_39411_, _39221_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_39412_, _39411_, _39222_);
  nor (_39413_, _39412_, _39284_);
  nor (_39414_, _39413_, _39410_);
  and (_39415_, _39414_, _39232_);
  not (_39416_, _39415_);
  nor (_39417_, _39416_, _39408_);
  and (_39418_, _39231_, _39071_);
  or (_39419_, _39418_, _39417_);
  nor (_19922_, _39419_, rst);
  and (_39420_, _27343_, _27211_);
  and (_39421_, _39271_, _39420_);
  and (_39422_, _39421_, _31308_);
  nand (_39423_, _39422_, _31265_);
  or (_39424_, _39422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39425_, _39424_, _31351_);
  and (_39426_, _39425_, _39423_);
  and (_39427_, _38620_, _39237_);
  nand (_39428_, _39427_, _38704_);
  or (_39429_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39430_, _39429_, _30651_);
  and (_39431_, _39430_, _39428_);
  not (_39432_, _30640_);
  and (_39433_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_39434_, _39433_, rst);
  or (_39435_, _39434_, _39431_);
  or (_31130_, _39435_, _39426_);
  and (_39436_, _39420_, _27847_);
  and (_39437_, _39436_, _31308_);
  nand (_39438_, _39437_, _31265_);
  or (_39439_, _39437_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39440_, _39439_, _31351_);
  and (_39441_, _39440_, _39438_);
  and (_39442_, _39111_, _38619_);
  and (_39443_, _39442_, _39237_);
  nand (_39444_, _39443_, _38704_);
  or (_39445_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39446_, _39445_, _30651_);
  and (_39447_, _39446_, _39444_);
  and (_39448_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_39449_, _39448_, rst);
  or (_39450_, _39449_, _39447_);
  or (_31153_, _39450_, _39441_);
  and (_39451_, _39095_, _27211_);
  and (_39452_, _39451_, _39271_);
  and (_39453_, _39452_, _31308_);
  nand (_39454_, _39453_, _31265_);
  or (_39455_, _39453_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_39456_, _39455_, _31351_);
  and (_39457_, _39456_, _39454_);
  and (_39458_, _39238_, _38619_);
  and (_39459_, _39458_, _39237_);
  not (_39460_, _39459_);
  nor (_39461_, _39460_, _38704_);
  and (_39462_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_39463_, _39462_, _39461_);
  and (_39464_, _39463_, _30651_);
  and (_39465_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_39466_, _39465_, rst);
  or (_39467_, _39466_, _39464_);
  or (_31176_, _39467_, _39457_);
  and (_39468_, _39451_, _27847_);
  and (_39469_, _39468_, _31308_);
  nand (_39470_, _39469_, _31265_);
  or (_39471_, _39469_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_39472_, _39471_, _31351_);
  and (_39473_, _39472_, _39470_);
  nor (_39474_, _27825_, _27343_);
  and (_39475_, _38619_, _39474_);
  and (_39476_, _39475_, _39237_);
  not (_39477_, _39476_);
  nor (_39478_, _39477_, _38704_);
  and (_39479_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_39480_, _39479_, _39478_);
  and (_39481_, _39480_, _30651_);
  and (_39482_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_39483_, _39482_, rst);
  or (_39484_, _39483_, _39481_);
  or (_31199_, _39484_, _39473_);
  or (_39485_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_39486_, _39485_, _31351_);
  and (_39487_, _39421_, _27003_);
  nand (_39488_, _39487_, _31265_);
  and (_39489_, _39488_, _39486_);
  nand (_39490_, _39427_, _38682_);
  and (_39491_, _39490_, _30651_);
  and (_39492_, _39491_, _39485_);
  not (_39493_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_39494_, _30640_, _39493_);
  or (_39495_, _39494_, rst);
  or (_39496_, _39495_, _39492_);
  or (_40808_, _39496_, _39489_);
  and (_39497_, _32604_, _27650_);
  and (_39498_, _39497_, _38620_);
  nand (_39499_, _39498_, _31265_);
  or (_39500_, _39498_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39501_, _39500_, _31351_);
  and (_39502_, _39501_, _39499_);
  nand (_39503_, _39427_, _38672_);
  or (_39504_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39505_, _39504_, _30651_);
  and (_39506_, _39505_, _39503_);
  and (_39507_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_39508_, _39507_, rst);
  or (_39509_, _39508_, _39506_);
  or (_40810_, _39509_, _39502_);
  not (_39510_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  not (_39511_, _34073_);
  and (_39512_, _39421_, _39511_);
  nor (_39513_, _39512_, _39510_);
  and (_39514_, _33377_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39515_, _39514_, _33366_);
  and (_39516_, _39515_, _39421_);
  or (_39517_, _39516_, _39513_);
  and (_39518_, _39517_, _31351_);
  nand (_39519_, _39427_, _38665_);
  or (_39520_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39521_, _39520_, _30651_);
  and (_39522_, _39521_, _39519_);
  nor (_39523_, _30640_, _39510_);
  or (_39524_, _39523_, rst);
  or (_39525_, _39524_, _39522_);
  or (_40812_, _39525_, _39518_);
  and (_39526_, _39421_, _34052_);
  nand (_39527_, _39526_, _31265_);
  or (_39528_, _39526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39529_, _39528_, _31351_);
  and (_39530_, _39529_, _39527_);
  nand (_39531_, _39427_, _38658_);
  or (_39532_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39533_, _39532_, _30651_);
  and (_39534_, _39533_, _39531_);
  and (_39535_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_39536_, _39535_, rst);
  or (_39537_, _39536_, _39534_);
  or (_40814_, _39537_, _39530_);
  not (_39538_, _39421_);
  or (_39539_, _39538_, _34813_);
  and (_39540_, _39539_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39541_, _34802_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39542_, _39541_, _34845_);
  and (_39543_, _39542_, _39421_);
  or (_39544_, _39543_, _39540_);
  and (_39545_, _39544_, _31351_);
  nand (_39546_, _39427_, _38650_);
  or (_39547_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39548_, _39547_, _30651_);
  and (_39549_, _39548_, _39546_);
  and (_39550_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39551_, _39550_, rst);
  or (_39552_, _39551_, _39549_);
  or (_40816_, _39552_, _39545_);
  and (_39553_, _39421_, _35607_);
  nand (_39554_, _39553_, _31265_);
  or (_39555_, _39553_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39556_, _39555_, _31351_);
  and (_39557_, _39556_, _39554_);
  nand (_39566_, _39427_, _38642_);
  or (_39577_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39588_, _39577_, _30651_);
  and (_39597_, _39588_, _39566_);
  and (_39603_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39614_, _39603_, rst);
  or (_39625_, _39614_, _39597_);
  or (_40818_, _39625_, _39557_);
  and (_39646_, _39421_, _36336_);
  nand (_39657_, _39646_, _31265_);
  or (_39668_, _39646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39679_, _39668_, _31351_);
  and (_39690_, _39679_, _39657_);
  nand (_39701_, _39427_, _38635_);
  or (_39712_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39723_, _39712_, _30651_);
  and (_39734_, _39723_, _39701_);
  and (_39745_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_39756_, _39745_, rst);
  or (_39767_, _39756_, _39734_);
  or (_40820_, _39767_, _39690_);
  and (_39771_, _39436_, _27003_);
  nand (_39772_, _39771_, _31265_);
  or (_39773_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39774_, _39773_, _31351_);
  and (_39775_, _39774_, _39772_);
  nand (_39776_, _39443_, _38682_);
  and (_39777_, _39776_, _30651_);
  and (_39778_, _39777_, _39773_);
  not (_39779_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_39780_, _30640_, _39779_);
  or (_39781_, _39780_, rst);
  or (_39782_, _39781_, _39778_);
  or (_40821_, _39782_, _39775_);
  and (_39783_, _39436_, _32604_);
  nand (_39784_, _39783_, _31265_);
  or (_39785_, _39783_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39786_, _39785_, _31351_);
  and (_39787_, _39786_, _39784_);
  nand (_39788_, _39443_, _38672_);
  or (_39789_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39790_, _39789_, _30651_);
  and (_39791_, _39790_, _39788_);
  and (_39792_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39793_, _39792_, rst);
  or (_39794_, _39793_, _39791_);
  or (_40823_, _39794_, _39787_);
  and (_39795_, _39436_, _33344_);
  nand (_39796_, _39795_, _31265_);
  or (_39797_, _39795_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39798_, _39797_, _31351_);
  and (_39799_, _39798_, _39796_);
  nand (_39800_, _39443_, _38665_);
  or (_39801_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39802_, _39801_, _30651_);
  and (_39803_, _39802_, _39800_);
  and (_39804_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_39805_, _39804_, rst);
  or (_39806_, _39805_, _39803_);
  or (_40825_, _39806_, _39799_);
  and (_39807_, _39436_, _34052_);
  nand (_39808_, _39807_, _31265_);
  or (_39809_, _39807_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39810_, _39809_, _31351_);
  and (_39811_, _39810_, _39808_);
  nand (_39812_, _39443_, _38658_);
  or (_39813_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39814_, _39813_, _30651_);
  and (_39815_, _39814_, _39812_);
  and (_39816_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39817_, _39816_, rst);
  or (_39818_, _39817_, _39815_);
  or (_40827_, _39818_, _39811_);
  and (_39819_, _39436_, _34791_);
  nand (_39820_, _39819_, _31265_);
  or (_39821_, _39819_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39822_, _39821_, _31351_);
  and (_39823_, _39822_, _39820_);
  nand (_39824_, _39443_, _38650_);
  or (_39825_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39826_, _39825_, _30651_);
  and (_39827_, _39826_, _39824_);
  and (_39828_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39829_, _39828_, rst);
  or (_39830_, _39829_, _39827_);
  or (_40829_, _39830_, _39823_);
  and (_39831_, _39436_, _35607_);
  nand (_39832_, _39831_, _31265_);
  or (_39833_, _39831_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39834_, _39833_, _31351_);
  and (_39835_, _39834_, _39832_);
  nand (_39836_, _39443_, _38642_);
  or (_39837_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39838_, _39837_, _30651_);
  and (_39839_, _39838_, _39836_);
  and (_39840_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39841_, _39840_, rst);
  or (_39842_, _39841_, _39839_);
  or (_40831_, _39842_, _39835_);
  and (_39843_, _39436_, _36336_);
  nand (_39844_, _39843_, _31265_);
  or (_39845_, _39843_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39846_, _39845_, _31351_);
  and (_39847_, _39846_, _39844_);
  nand (_39848_, _39443_, _38635_);
  or (_39849_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39850_, _39849_, _30651_);
  and (_39851_, _39850_, _39848_);
  and (_39852_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39853_, _39852_, rst);
  or (_39854_, _39853_, _39851_);
  or (_40833_, _39854_, _39847_);
  nand (_39855_, _39459_, _31265_);
  or (_39856_, _39459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39857_, _39856_, _31351_);
  and (_39858_, _39857_, _39855_);
  and (_39859_, _39459_, _38683_);
  not (_39860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_39861_, _39459_, _39860_);
  or (_39862_, _39861_, _39859_);
  and (_39863_, _39862_, _30651_);
  nor (_39864_, _30640_, _39860_);
  or (_39865_, _39864_, rst);
  or (_39866_, _39865_, _39863_);
  or (_40835_, _39866_, _39858_);
  and (_39867_, _39452_, _32604_);
  nand (_39868_, _39867_, _31265_);
  or (_39869_, _39867_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39870_, _39869_, _31351_);
  and (_39871_, _39870_, _39868_);
  nor (_39872_, _39460_, _38672_);
  and (_39873_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39874_, _39873_, _39872_);
  and (_39875_, _39874_, _30651_);
  and (_39876_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39877_, _39876_, rst);
  or (_39878_, _39877_, _39875_);
  or (_40837_, _39878_, _39871_);
  and (_39879_, _39452_, _33344_);
  nand (_39880_, _39879_, _31265_);
  or (_39881_, _39879_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39882_, _39881_, _31351_);
  and (_39883_, _39882_, _39880_);
  nor (_39884_, _39460_, _38665_);
  and (_39885_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39886_, _39885_, _39884_);
  and (_39887_, _39886_, _30651_);
  and (_39888_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39889_, _39888_, rst);
  or (_39890_, _39889_, _39887_);
  or (_40839_, _39890_, _39883_);
  and (_39891_, _39452_, _34052_);
  nand (_39892_, _39891_, _31265_);
  or (_39893_, _39891_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39894_, _39893_, _31351_);
  and (_39895_, _39894_, _39892_);
  nor (_39896_, _39460_, _38658_);
  and (_39897_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39898_, _39897_, _39896_);
  and (_39899_, _39898_, _30651_);
  and (_39900_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39901_, _39900_, rst);
  or (_39902_, _39901_, _39899_);
  or (_40841_, _39902_, _39895_);
  and (_39903_, _39452_, _34791_);
  nand (_39904_, _39903_, _31265_);
  or (_39905_, _39903_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39906_, _39905_, _31351_);
  and (_39907_, _39906_, _39904_);
  nor (_39908_, _39460_, _38650_);
  and (_39909_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39910_, _39909_, _39908_);
  and (_39911_, _39910_, _30651_);
  and (_39912_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39913_, _39912_, rst);
  or (_39914_, _39913_, _39911_);
  or (_40843_, _39914_, _39907_);
  and (_39915_, _39452_, _35607_);
  nand (_39916_, _39915_, _31265_);
  or (_39917_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39918_, _39917_, _31351_);
  and (_39919_, _39918_, _39916_);
  nor (_39920_, _39460_, _38642_);
  and (_39921_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39922_, _39921_, _39920_);
  and (_39923_, _39922_, _30651_);
  and (_39924_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39925_, _39924_, rst);
  or (_39926_, _39925_, _39923_);
  or (_40845_, _39926_, _39919_);
  and (_39927_, _39452_, _36336_);
  nand (_39928_, _39927_, _31265_);
  or (_39929_, _39927_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39930_, _39929_, _31351_);
  and (_39931_, _39930_, _39928_);
  nor (_39932_, _39460_, _38635_);
  and (_39933_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39934_, _39933_, _39932_);
  and (_39935_, _39934_, _30651_);
  and (_39936_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39937_, _39936_, rst);
  or (_39938_, _39937_, _39935_);
  or (_40847_, _39938_, _39931_);
  and (_39939_, _39468_, _27003_);
  nand (_39940_, _39939_, _31265_);
  or (_39941_, _39476_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39942_, _39941_, _31351_);
  and (_39943_, _39942_, _39940_);
  nand (_39944_, _39476_, _38682_);
  and (_39945_, _39941_, _30651_);
  and (_39946_, _39945_, _39944_);
  not (_39947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_39948_, _30640_, _39947_);
  or (_39949_, _39948_, rst);
  or (_39950_, _39949_, _39946_);
  or (_40849_, _39950_, _39943_);
  and (_39951_, _39468_, _32604_);
  nand (_39952_, _39951_, _31265_);
  or (_39953_, _39951_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39954_, _39953_, _31351_);
  and (_39955_, _39954_, _39952_);
  nor (_39956_, _39477_, _38672_);
  and (_39957_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39958_, _39957_, _39956_);
  and (_39959_, _39958_, _30651_);
  and (_39960_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39961_, _39960_, rst);
  or (_39962_, _39961_, _39959_);
  or (_40851_, _39962_, _39955_);
  and (_39963_, _39468_, _33344_);
  nand (_39964_, _39963_, _31265_);
  or (_39965_, _39963_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_39966_, _39965_, _31351_);
  and (_39967_, _39966_, _39964_);
  nor (_39968_, _39477_, _38665_);
  and (_39969_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39970_, _39969_, _39968_);
  and (_39971_, _39970_, _30651_);
  and (_39972_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39973_, _39972_, rst);
  or (_39974_, _39973_, _39971_);
  or (_40852_, _39974_, _39967_);
  and (_39975_, _39468_, _34052_);
  nand (_39976_, _39975_, _31265_);
  or (_39977_, _39975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_39978_, _39977_, _31351_);
  and (_39979_, _39978_, _39976_);
  nor (_39984_, _39477_, _38658_);
  and (_39986_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39987_, _39986_, _39984_);
  and (_39988_, _39987_, _30651_);
  and (_39989_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39990_, _39989_, rst);
  or (_39991_, _39990_, _39988_);
  or (_40854_, _39991_, _39979_);
  and (_39992_, _39468_, _34791_);
  nand (_39993_, _39992_, _31265_);
  or (_39994_, _39992_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_39995_, _39994_, _31351_);
  and (_39996_, _39995_, _39993_);
  nor (_39997_, _39477_, _38650_);
  and (_39998_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39999_, _39998_, _39997_);
  and (_40000_, _39999_, _30651_);
  and (_40001_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_40002_, _40001_, rst);
  or (_40003_, _40002_, _40000_);
  or (_40856_, _40003_, _39996_);
  and (_40004_, _39468_, _35607_);
  nand (_40005_, _40004_, _31265_);
  or (_40006_, _40004_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_40007_, _40006_, _31351_);
  and (_40008_, _40007_, _40005_);
  nor (_40009_, _39477_, _38642_);
  and (_40010_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_40011_, _40010_, _40009_);
  and (_40012_, _40011_, _30651_);
  and (_40020_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_40031_, _40020_, rst);
  or (_40042_, _40031_, _40012_);
  or (_40858_, _40042_, _40008_);
  and (_40044_, _39468_, _36336_);
  nand (_40045_, _40044_, _31265_);
  or (_40046_, _40044_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_40047_, _40046_, _31351_);
  and (_40048_, _40047_, _40045_);
  nor (_40049_, _39477_, _38635_);
  and (_40050_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_40051_, _40050_, _40049_);
  and (_40052_, _40051_, _30651_);
  and (_40053_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_40054_, _40053_, rst);
  or (_40055_, _40054_, _40052_);
  or (_40860_, _40055_, _40048_);
  and (_41311_, t0_i, _43100_);
  and (_41314_, t1_i, _43100_);
  nor (_40056_, _26740_, _27650_);
  and (_40057_, _40056_, _38621_);
  and (_40058_, _40057_, _30651_);
  not (_40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_40060_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_40061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_40062_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _40061_);
  nor (_40063_, _40062_, _40060_);
  or (_40064_, _40063_, _40058_);
  and (_40065_, _40064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_40066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_40067_, t1_i);
  and (_40068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _40067_);
  nor (_40069_, _40068_, _40066_);
  not (_40071_, _40069_);
  not (_40077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_40078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _40077_);
  nor (_40079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_40080_, _40079_);
  and (_40081_, _40080_, _40078_);
  and (_40082_, _40081_, _40071_);
  not (_40083_, _40082_);
  nand (_40084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_40085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or (_40086_, _40085_, _40084_);
  nor (_40087_, _40086_, _40083_);
  and (_40088_, _40087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_40089_, _40088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_40090_, _40089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_40091_, _40090_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_40092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_40093_, _40086_, _40092_);
  and (_40094_, _40093_, _40082_);
  and (_40095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_40096_, _40095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_40097_, _40096_, _40094_);
  nor (_40098_, _40097_, _40063_);
  and (_40099_, _40098_, _40091_);
  and (_40100_, _40097_, _40060_);
  and (_40101_, _40100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_40102_, _40101_, _40099_);
  nor (_40103_, _40102_, _40058_);
  or (_40104_, _40103_, _40065_);
  and (_40105_, _34052_, _27661_);
  and (_40106_, _40105_, _38620_);
  and (_40107_, _40106_, _30651_);
  not (_40108_, _40107_);
  and (_40109_, _40108_, _40104_);
  nor (_40110_, _40108_, _38704_);
  or (_40111_, _40110_, _40109_);
  and (_41317_, _40111_, _43100_);
  not (_40112_, _30651_);
  nor (_40113_, _40112_, _27650_);
  and (_40114_, _40113_, _38751_);
  and (_40115_, _40114_, _43100_);
  and (_40116_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_40117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40118_, _40117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_40119_, _40096_, _40093_);
  and (_40120_, _40119_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_40121_, _40120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_40122_, _40121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_40123_, _40122_, _40082_);
  and (_40124_, _40123_, _40118_);
  and (_40125_, _40124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40126_, _40125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_40127_, _40125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_40128_, _40127_, _40126_);
  and (_40129_, _40128_, _40062_);
  and (_40130_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_40131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_40132_, _40131_, _40093_);
  and (_40133_, _40132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_40134_, _40133_, _40082_);
  and (_40135_, _40134_, _40118_);
  and (_40136_, _40135_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40137_, _40136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_40138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_40139_, _40136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_40140_, _40139_, _40138_);
  nor (_40141_, _40140_, _40137_);
  or (_40142_, _40141_, _40130_);
  nor (_40143_, _40142_, _40129_);
  nor (_40144_, _40143_, _40058_);
  not (_40145_, _38704_);
  and (_40146_, _40058_, _40145_);
  or (_40147_, _40146_, _40144_);
  nor (_40148_, _40114_, rst);
  and (_40149_, _40148_, _40147_);
  or (_41320_, _40149_, _40116_);
  and (_40150_, _40083_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or (_40151_, _40150_, _40126_);
  and (_40152_, _40151_, _40062_);
  or (_40153_, _40150_, _40137_);
  and (_40154_, _40153_, _40138_);
  nand (_40155_, _40082_, _40059_);
  and (_40160_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_40167_, _40160_, _40155_);
  or (_40168_, _40167_, _40100_);
  or (_40169_, _40168_, _40154_);
  nor (_40170_, _40169_, _40152_);
  nor (_40171_, _40170_, _40058_);
  and (_41323_, _40171_, _40148_);
  and (_40172_, _40113_, _34791_);
  and (_40173_, _40172_, _38620_);
  nor (_40174_, _40173_, rst);
  and (_40175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_40177_, _40176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40178_, _40177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40179_, _40178_, _40175_);
  and (_40180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_40181_, _40180_, _40179_);
  or (_40182_, _40181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_40183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_40184_, _40183_);
  and (_40185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_40186_, _40185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_40187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_40188_, t0_i);
  and (_40189_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _40188_);
  nor (_40190_, _40189_, _40187_);
  not (_40191_, _40190_);
  not (_40192_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_40193_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_40194_, _40193_, _40192_);
  and (_40195_, _40194_, _40191_);
  and (_40196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_40197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_40198_, _40197_, _40196_);
  and (_40199_, _40198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_40200_, _40199_, _40195_);
  and (_40201_, _40200_, _40186_);
  and (_40202_, _40201_, _40184_);
  and (_40203_, _40202_, _40182_);
  not (_40204_, _40195_);
  and (_40205_, _40204_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and (_40206_, _40200_, _40179_);
  and (_40207_, _40206_, _40180_);
  and (_40208_, _40207_, _40183_);
  or (_40209_, _40208_, _40205_);
  nor (_40210_, _40209_, _40203_);
  and (_40211_, _40113_, _33344_);
  and (_40212_, _40211_, _38620_);
  nor (_40213_, _40212_, _40210_);
  and (_41326_, _40213_, _40174_);
  and (_40214_, _40113_, _38848_);
  nand (_40215_, _40214_, _38704_);
  and (_40216_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_40217_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _40217_);
  not (_40219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40220_, _40219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_40221_, _40220_, _40218_);
  not (_40222_, _40201_);
  and (_40223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40224_, _40223_, _40222_);
  or (_40225_, _40224_, _40221_);
  nand (_40226_, _40220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_40227_, _40226_, _40201_);
  and (_40228_, _40227_, _40225_);
  or (_40229_, _40228_, _40216_);
  or (_40230_, _40229_, _40173_);
  and (_40231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand (_40232_, _40231_, _40200_);
  nor (_40233_, _40232_, _40173_);
  or (_40234_, _40233_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_40235_, _40234_, _40230_);
  or (_40236_, _40235_, _40214_);
  and (_40238_, _40236_, _43100_);
  and (_41329_, _40238_, _40215_);
  nand (_40242_, _40173_, _38704_);
  not (_40243_, _40212_);
  not (_40244_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_40245_, _40199_, _40186_);
  and (_40246_, _40195_, _40217_);
  and (_40247_, _40246_, _40245_);
  and (_40248_, _40247_, _40179_);
  and (_40249_, _40248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_40250_, _40249_, _40244_);
  and (_40251_, _40249_, _40244_);
  or (_40252_, _40251_, _40250_);
  and (_40253_, _40252_, _40221_);
  and (_40254_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_40255_, _40254_, _40178_);
  and (_40256_, _40255_, _40175_);
  and (_40257_, _40256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40267_, _40257_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_40268_, _40254_, _40181_);
  and (_40269_, _40268_, _40267_);
  and (_40270_, _40269_, _40223_);
  and (_40271_, _40206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40272_, _40271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_40273_, _40207_, _40184_);
  and (_40274_, _40273_, _40272_);
  or (_40275_, _40274_, _40270_);
  or (_40276_, _40275_, _40253_);
  or (_40277_, _40276_, _40173_);
  and (_40278_, _40277_, _40243_);
  and (_40279_, _40278_, _40242_);
  and (_40280_, _40212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_40281_, _40280_, _40279_);
  and (_41332_, _40281_, _43100_);
  or (_40282_, _40254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_40283_, _40223_, _43100_);
  nand (_40284_, _40283_, _40282_);
  nor (_40285_, _40284_, _40173_);
  not (_40286_, _40254_);
  nor (_40287_, _40286_, _40181_);
  nor (_40288_, _40287_, _40212_);
  and (_41335_, _40288_, _40285_);
  and (_40289_, _40113_, _38622_);
  or (_40290_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_40291_, _40290_, _43100_);
  nand (_40292_, _40289_, _38704_);
  and (_41338_, _40292_, _40291_);
  and (_40293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_40294_, _40293_, _40058_);
  and (_40295_, _40294_, _40082_);
  or (_40296_, _40295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  not (_40297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_40298_, _40060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_40299_, _40298_, _40119_);
  nor (_40300_, _40299_, _40058_);
  nor (_40301_, _40300_, _40297_);
  nand (_40302_, _40301_, _40295_);
  and (_40303_, _40302_, _40148_);
  and (_40304_, _40303_, _40296_);
  and (_40305_, _40115_, _38683_);
  or (_41820_, _40305_, _40304_);
  not (_40306_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_40307_, _40294_, _40306_);
  not (_40308_, _40293_);
  and (_40309_, _40082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_40310_, _40309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_40311_, _40309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_40312_, _40311_, _40310_);
  and (_40313_, _40312_, _40308_);
  and (_40314_, _40090_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_40315_, _40314_, _40060_);
  and (_40316_, _40315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_40317_, _40316_, _40313_);
  nor (_40318_, _40317_, _40058_);
  or (_40319_, _40318_, _40307_);
  and (_40320_, _40319_, _40108_);
  nor (_40321_, _40108_, _38672_);
  or (_40322_, _40321_, _40320_);
  and (_41822_, _40322_, _43100_);
  not (_40323_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_40324_, _40294_, _40323_);
  nor (_40325_, _40310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_40326_, _40310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_40327_, _40326_, _40325_);
  and (_40328_, _40327_, _40308_);
  and (_40329_, _40100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_40330_, _40329_, _40328_);
  nor (_40331_, _40330_, _40058_);
  or (_40332_, _40331_, _40324_);
  and (_40333_, _40332_, _40148_);
  not (_40334_, _38665_);
  and (_40335_, _40115_, _40334_);
  or (_41823_, _40335_, _40333_);
  not (_40336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_40337_, _40294_, _40336_);
  or (_40338_, _40326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_40339_, _40293_, _40087_);
  and (_40340_, _40339_, _40338_);
  and (_40341_, _40100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_40342_, _40341_, _40340_);
  nor (_40343_, _40342_, _40058_);
  or (_40344_, _40343_, _40337_);
  and (_40345_, _40344_, _40148_);
  not (_40346_, _38658_);
  and (_40347_, _40115_, _40346_);
  or (_41825_, _40347_, _40345_);
  nor (_40348_, _40294_, _40092_);
  or (_40349_, _40087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_40350_, _40293_, _40094_);
  and (_40351_, _40350_, _40349_);
  and (_40352_, _40100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_40353_, _40352_, _40351_);
  nor (_40354_, _40353_, _40058_);
  or (_40355_, _40354_, _40348_);
  and (_40356_, _40355_, _40148_);
  not (_40357_, _38650_);
  and (_40358_, _40115_, _40357_);
  or (_41827_, _40358_, _40356_);
  and (_40359_, _40064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_40360_, _40315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_40361_, _40063_);
  and (_40362_, _40094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_40363_, _40094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_40364_, _40363_, _40362_);
  and (_40365_, _40364_, _40361_);
  nor (_40366_, _40365_, _40360_);
  nor (_40367_, _40366_, _40058_);
  or (_40368_, _40367_, _40359_);
  and (_40369_, _40368_, _40148_);
  not (_40370_, _38642_);
  and (_40371_, _40115_, _40370_);
  or (_41829_, _40371_, _40369_);
  and (_40372_, _40064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_40373_, _40060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40374_, _40373_, _40082_);
  and (_40375_, _40374_, _40119_);
  or (_40376_, _40362_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_40377_, _40376_, _40361_);
  nor (_40378_, _40377_, _40090_);
  nor (_40379_, _40378_, _40375_);
  nor (_40380_, _40379_, _40058_);
  or (_40381_, _40380_, _40372_);
  and (_40382_, _40381_, _40148_);
  not (_40383_, _38635_);
  and (_40384_, _40115_, _40383_);
  or (_41831_, _40384_, _40382_);
  not (_40385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_40386_, _40094_, _40061_);
  nor (_40387_, _40096_, _40059_);
  not (_40388_, _40387_);
  and (_40389_, _40388_, _40386_);
  nor (_40390_, _40389_, _40385_);
  and (_40391_, _40389_, _40385_);
  or (_40392_, _40391_, _40390_);
  or (_40393_, _40392_, _40058_);
  nand (_40394_, _40058_, _38682_);
  and (_40395_, _40394_, _40148_);
  and (_40396_, _40395_, _40393_);
  and (_40397_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_41833_, _40397_, _40396_);
  nand (_40398_, _40058_, _38672_);
  not (_40399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not (_40400_, _40062_);
  nor (_40401_, _40097_, _40400_);
  not (_40402_, _40401_);
  nor (_40403_, _40386_, _40062_);
  nor (_40404_, _40403_, _40385_);
  and (_40405_, _40404_, _40402_);
  nor (_40406_, _40405_, _40399_);
  and (_40407_, _40405_, _40399_);
  or (_40408_, _40407_, _40406_);
  or (_40409_, _40408_, _40058_);
  and (_40410_, _40409_, _40148_);
  and (_40411_, _40410_, _40398_);
  and (_40412_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_41835_, _40412_, _40411_);
  and (_40413_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand (_40414_, _40058_, _38665_);
  and (_40415_, _40131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_40416_, _40415_, _40094_);
  nand (_40417_, _40416_, _40061_);
  or (_40418_, _40417_, _40387_);
  and (_40419_, _40418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_40420_, _40387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_40421_, _40420_);
  not (_40422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_40423_, _40131_, _40422_);
  and (_40424_, _40423_, _40094_);
  and (_40425_, _40424_, _40421_);
  or (_40426_, _40425_, _40419_);
  or (_40427_, _40426_, _40058_);
  and (_40428_, _40427_, _40148_);
  and (_40429_, _40428_, _40414_);
  or (_41837_, _40429_, _40413_);
  and (_40430_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_40431_, _40058_, _38658_);
  and (_40432_, _40416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_40433_, _40432_, _40096_);
  or (_40434_, _40123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_40435_, _40434_, _40062_);
  nor (_40436_, _40435_, _40433_);
  and (_40437_, _40417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_40438_, _40417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_40439_, _40438_, _40437_);
  and (_40440_, _40439_, _40400_);
  or (_40441_, _40440_, _40436_);
  or (_40442_, _40441_, _40058_);
  and (_40443_, _40442_, _40148_);
  and (_40444_, _40443_, _40431_);
  or (_41839_, _40444_, _40430_);
  nand (_40445_, _40058_, _38650_);
  or (_40446_, _40433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_40447_, _40446_, _40062_);
  and (_40448_, _40433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_40449_, _40448_, _40447_);
  and (_40450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40451_, _40134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_40452_, _40451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_40453_, _40451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40454_, _40453_, _40452_);
  and (_40455_, _40454_, _40138_);
  or (_40456_, _40455_, _40450_);
  or (_40457_, _40456_, _40449_);
  or (_40458_, _40457_, _40058_);
  and (_40459_, _40458_, _40148_);
  and (_40460_, _40459_, _40445_);
  and (_40461_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_41840_, _40461_, _40460_);
  nand (_40462_, _40058_, _38642_);
  and (_40463_, _40432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40464_, _40463_, _40138_);
  and (_40465_, _40448_, _40062_);
  nor (_40466_, _40465_, _40464_);
  and (_40467_, _40466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_40468_, _40466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_40469_, _40468_, _40467_);
  or (_40470_, _40469_, _40058_);
  and (_40471_, _40470_, _40148_);
  and (_40472_, _40471_, _40462_);
  and (_40473_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_41842_, _40473_, _40472_);
  nand (_40474_, _40058_, _38635_);
  and (_40475_, _40463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_40476_, _40421_, _40475_);
  or (_40477_, _40476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_40478_, _40476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40479_, _40478_, _40477_);
  or (_40480_, _40479_, _40058_);
  and (_40481_, _40480_, _40148_);
  and (_40482_, _40481_, _40474_);
  and (_40483_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_41844_, _40483_, _40482_);
  nor (_40484_, _40204_, _40173_);
  or (_40485_, _40484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_40486_, _40195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_40487_, _40220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40488_, _40487_, _40245_);
  nand (_40489_, _40488_, _40486_);
  or (_40490_, _40489_, _40173_);
  and (_40491_, _40490_, _40485_);
  or (_40492_, _40491_, _40212_);
  nand (_40493_, _40212_, _38682_);
  and (_40494_, _40493_, _43100_);
  and (_41846_, _40494_, _40492_);
  not (_40495_, _40214_);
  nor (_40496_, _40486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_40497_, _40486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_40498_, _40497_, _40496_);
  and (_40499_, _40220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40500_, _40499_, _40201_);
  nor (_40501_, _40500_, _40498_);
  nor (_40502_, _40501_, _40173_);
  and (_40503_, _40173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_40504_, _40503_, _40502_);
  and (_40505_, _40504_, _40495_);
  nor (_40506_, _40243_, _38672_);
  or (_40507_, _40506_, _40505_);
  and (_41848_, _40507_, _43100_);
  nor (_40508_, _40497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_40509_, _40486_, _40196_);
  nor (_40510_, _40509_, _40508_);
  and (_40511_, _40220_, _40201_);
  and (_40512_, _40511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_40513_, _40512_, _40510_);
  nor (_40514_, _40513_, _40173_);
  and (_40515_, _40173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_40516_, _40515_, _40514_);
  and (_40517_, _40516_, _40495_);
  nor (_40518_, _40243_, _38665_);
  or (_40519_, _40518_, _40517_);
  and (_41850_, _40519_, _43100_);
  and (_40520_, _40198_, _40195_);
  nor (_40521_, _40509_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_40522_, _40521_, _40520_);
  and (_40523_, _40511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_40524_, _40523_, _40522_);
  nor (_40525_, _40524_, _40173_);
  and (_40526_, _40173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_40527_, _40526_, _40525_);
  and (_40528_, _40527_, _40495_);
  nor (_40529_, _40243_, _38658_);
  or (_40530_, _40529_, _40528_);
  and (_41852_, _40530_, _43100_);
  nor (_40531_, _40520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_40532_, _40531_, _40200_);
  and (_40533_, _40511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_40534_, _40533_, _40532_);
  or (_40535_, _40534_, _40173_);
  not (_40536_, _40173_);
  or (_40537_, _40536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_40538_, _40537_, _40243_);
  and (_40539_, _40538_, _40535_);
  nor (_40540_, _40243_, _38650_);
  or (_40541_, _40540_, _40539_);
  and (_41854_, _40541_, _43100_);
  nand (_40542_, _40214_, _38642_);
  or (_40543_, _40536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_40544_, _40511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40545_, _40200_, _40184_);
  or (_40546_, _40545_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_40547_, _40545_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_40548_, _40547_);
  or (_40549_, _40548_, _40173_);
  and (_40550_, _40549_, _40546_);
  or (_40551_, _40550_, _40544_);
  and (_40552_, _40551_, _40543_);
  or (_40553_, _40552_, _40214_);
  and (_40554_, _40553_, _43100_);
  and (_41855_, _40554_, _40542_);
  and (_40555_, _40220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_40556_, _40555_, _40195_);
  and (_40557_, _40556_, _40245_);
  nor (_40558_, _40548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_40559_, _40558_, _40557_);
  nor (_40560_, _40559_, _40173_);
  and (_40561_, _40549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_40562_, _40561_, _40560_);
  and (_40563_, _40562_, _40495_);
  nor (_40564_, _40243_, _38635_);
  or (_40565_, _40564_, _40563_);
  and (_41857_, _40565_, _43100_);
  or (_40566_, _40247_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40567_, _40566_, _40221_);
  and (_40568_, _40247_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_40569_, _40568_, _40567_);
  and (_40570_, _40254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_40571_, _40254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40572_, _40571_, _40223_);
  nor (_40573_, _40572_, _40570_);
  and (_40574_, _40200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_40575_, _40200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40576_, _40575_, _40183_);
  nor (_40577_, _40576_, _40574_);
  or (_40578_, _40577_, _40573_);
  or (_40579_, _40578_, _40569_);
  or (_40580_, _40579_, _40173_);
  nand (_40581_, _40173_, _38682_);
  and (_40582_, _40581_, _40580_);
  or (_40583_, _40582_, _40214_);
  or (_40584_, _40495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_40585_, _40584_, _43100_);
  and (_41859_, _40585_, _40583_);
  nand (_40586_, _40173_, _38672_);
  or (_40587_, _40568_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40588_, _40245_, _40195_);
  and (_40589_, _40588_, _40176_);
  not (_40590_, _40589_);
  or (_40591_, _40590_, _40220_);
  and (_40592_, _40591_, _40221_);
  and (_40593_, _40592_, _40587_);
  not (_40594_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_40595_, _40570_, _40594_);
  and (_40596_, _40570_, _40594_);
  or (_40597_, _40596_, _40595_);
  and (_40598_, _40597_, _40223_);
  and (_40599_, _40574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_40600_, _40574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_40601_, _40600_, _40183_);
  nor (_40602_, _40601_, _40599_);
  or (_40603_, _40602_, _40598_);
  or (_40604_, _40603_, _40593_);
  or (_40605_, _40604_, _40173_);
  and (_40606_, _40605_, _40243_);
  and (_40607_, _40606_, _40586_);
  and (_40608_, _40212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_40609_, _40608_, _40607_);
  and (_41861_, _40609_, _43100_);
  nor (_40610_, _40536_, _38665_);
  or (_40611_, _40589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40612_, _40588_, _40177_);
  not (_40613_, _40612_);
  and (_40614_, _40613_, _40218_);
  and (_40615_, _40614_, _40611_);
  or (_40616_, _40599_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40617_, _40200_, _40177_);
  nor (_40618_, _40617_, _40184_);
  and (_40619_, _40618_, _40616_);
  and (_40620_, _40176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40621_, _40620_, _40254_);
  or (_40622_, _40621_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40623_, _40254_, _40177_);
  nand (_40624_, _40623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40625_, _40624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40626_, _40625_, _40622_);
  or (_40627_, _40626_, _40619_);
  nor (_40628_, _40627_, _40615_);
  nor (_40629_, _40628_, _40173_);
  or (_40630_, _40629_, _40214_);
  or (_40631_, _40630_, _40610_);
  or (_40632_, _40495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40633_, _40632_, _43100_);
  and (_41863_, _40633_, _40631_);
  nor (_40634_, _40536_, _38658_);
  not (_40635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40636_, _40612_, _40217_);
  nor (_40637_, _40636_, _40635_);
  and (_40638_, _40636_, _40635_);
  or (_40639_, _40638_, _40637_);
  and (_40640_, _40639_, _40221_);
  or (_40641_, _40623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_40642_, _40255_);
  and (_40643_, _40642_, _40223_);
  and (_40644_, _40643_, _40641_);
  or (_40645_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40646_, _40200_, _40178_);
  nor (_40647_, _40646_, _40184_);
  and (_40648_, _40647_, _40645_);
  or (_40649_, _40648_, _40644_);
  nor (_40650_, _40649_, _40640_);
  nor (_40651_, _40650_, _40173_);
  or (_40652_, _40651_, _40214_);
  or (_40653_, _40652_, _40634_);
  nand (_40654_, _40214_, _40635_);
  and (_40655_, _40654_, _43100_);
  and (_41865_, _40655_, _40653_);
  nand (_40656_, _40173_, _38650_);
  or (_40657_, _40646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40658_, _40599_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40659_, _40658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40660_, _40659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_40661_, _40660_, _40184_);
  and (_40662_, _40661_, _40657_);
  and (_40663_, _40588_, _40178_);
  or (_40664_, _40663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_40665_, _40663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40666_, _40665_, _40218_);
  and (_40667_, _40666_, _40664_);
  and (_40668_, _40255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_40669_, _40668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40670_, _40669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40671_, _40255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_40672_, _40671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40673_, _40672_, _40670_);
  or (_40674_, _40673_, _40667_);
  or (_40675_, _40674_, _40662_);
  or (_40676_, _40675_, _40173_);
  and (_40677_, _40676_, _40243_);
  and (_40678_, _40677_, _40656_);
  and (_40679_, _40212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_40680_, _40679_, _40678_);
  and (_41867_, _40680_, _43100_);
  nor (_40681_, _40536_, _38642_);
  not (_40682_, _40660_);
  nor (_40683_, _40682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40684_, _40682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_40685_, _40684_, _40683_);
  and (_40686_, _40685_, _40183_);
  nor (_40687_, _40665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_40688_, _40687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_40689_, _40687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40690_, _40689_, _40221_);
  and (_40691_, _40690_, _40688_);
  not (_40692_, _40256_);
  and (_40693_, _40692_, _40223_);
  or (_40694_, _40671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40695_, _40694_, _40693_);
  or (_40696_, _40695_, _40691_);
  or (_40697_, _40696_, _40686_);
  and (_40698_, _40697_, _40536_);
  or (_40699_, _40698_, _40214_);
  or (_40700_, _40699_, _40681_);
  or (_40701_, _40495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40702_, _40701_, _43100_);
  and (_41869_, _40702_, _40700_);
  nand (_40703_, _40173_, _38635_);
  or (_40704_, _40248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_40705_, _40704_, _40221_);
  nor (_40706_, _40705_, _40249_);
  or (_40707_, _40256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_40708_, _40257_);
  and (_40709_, _40708_, _40223_);
  and (_40710_, _40709_, _40707_);
  or (_40711_, _40206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_40712_, _40271_, _40184_);
  and (_40713_, _40712_, _40711_);
  or (_40714_, _40713_, _40710_);
  or (_40715_, _40714_, _40706_);
  or (_40716_, _40715_, _40173_);
  and (_40717_, _40716_, _40243_);
  and (_40718_, _40717_, _40703_);
  and (_40719_, _40212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40720_, _40719_, _40718_);
  and (_41870_, _40720_, _43100_);
  nor (_40721_, _40289_, _40219_);
  and (_40722_, _40289_, _38683_);
  or (_40723_, _40722_, _40721_);
  and (_41872_, _40723_, _43100_);
  or (_40724_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40725_, _40724_, _43100_);
  nand (_40726_, _40289_, _38672_);
  and (_41874_, _40726_, _40725_);
  or (_40727_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_40728_, _40727_, _43100_);
  nand (_40729_, _40289_, _38665_);
  and (_41876_, _40729_, _40728_);
  or (_40730_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_40731_, _40730_, _43100_);
  nand (_40732_, _40289_, _38658_);
  and (_41877_, _40732_, _40731_);
  or (_40733_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_40734_, _40733_, _43100_);
  nand (_40735_, _40289_, _38650_);
  and (_41879_, _40735_, _40734_);
  or (_40736_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_40737_, _40736_, _43100_);
  nand (_40738_, _40289_, _38642_);
  and (_41881_, _40738_, _40737_);
  or (_40739_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_40740_, _40739_, _43100_);
  nand (_40741_, _40289_, _38635_);
  and (_41883_, _40741_, _40740_);
  not (_40742_, _27825_);
  nor (_40743_, _39246_, _27650_);
  nand (_40744_, _40743_, _40742_);
  nor (_40745_, _40744_, _27496_);
  and (_40746_, _40745_, _39451_);
  and (_40747_, _40746_, _31308_);
  nand (_40748_, _40747_, _31265_);
  and (_40749_, _38617_, _31308_);
  and (_40750_, _40749_, _39475_);
  nor (_40751_, _40747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nor (_40752_, _40751_, _40750_);
  and (_40753_, _40752_, _40748_);
  and (_40754_, _39469_, _30651_);
  and (_40755_, _40754_, _40145_);
  or (_40756_, _40755_, _40753_);
  and (_43045_, _40756_, _43100_);
  and (_40757_, _40113_, _27003_);
  and (_40758_, _40757_, _39458_);
  not (_40759_, _40758_);
  and (_40760_, _27825_, _27661_);
  and (_40761_, _40760_, _39247_);
  and (_40762_, _40761_, _39451_);
  and (_40763_, _40762_, _31308_);
  or (_40764_, _40763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_40765_, _40764_, _40759_);
  nand (_40766_, _40763_, _31265_);
  and (_40767_, _40766_, _40765_);
  nor (_40768_, _40759_, _38704_);
  or (_40769_, _40768_, _40767_);
  and (_43048_, _40769_, _43100_);
  and (_40770_, _40757_, _38620_);
  and (_40771_, _40743_, _27825_);
  and (_40772_, _40771_, _27507_);
  and (_40773_, _40772_, _39420_);
  nand (_40774_, _40773_, _26981_);
  and (_40775_, _40774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40776_, _40775_, _40770_);
  or (_40777_, _26992_, _33333_);
  and (_40778_, _40777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40779_, _40778_, _39222_);
  and (_40780_, _40779_, _40773_);
  or (_40781_, _40780_, _40776_);
  nand (_40782_, _40770_, _38635_);
  and (_40783_, _40782_, _43100_);
  and (_43050_, _40783_, _40781_);
  not (_40784_, _40770_);
  nor (_40785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_40786_, _40785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not (_40787_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_40788_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40790_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40789_);
  and (_40791_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40792_, _40791_, _40790_);
  nor (_40793_, _40792_, _40788_);
  or (_40794_, _40793_, _40787_);
  and (_40795_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_40796_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_40797_, _40796_, _40795_);
  nor (_40798_, _40797_, _40788_);
  and (_40799_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40789_);
  and (_40800_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40801_, _40800_, _40799_);
  nand (_40802_, _40801_, _40798_);
  or (_40803_, _40802_, _40794_);
  and (_40804_, _40803_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_40805_, _40804_, _40786_);
  and (_40806_, _38620_, _31308_);
  and (_40807_, _40806_, _40743_);
  or (_40809_, _40807_, _40805_);
  and (_40811_, _40809_, _40784_);
  nand (_40813_, _40807_, _31265_);
  and (_40815_, _40813_, _40811_);
  nor (_40817_, _40784_, _38704_);
  or (_40819_, _40817_, _40815_);
  and (_43052_, _40819_, _43100_);
  and (_40822_, _40057_, _31351_);
  nand (_40824_, _40822_, _31265_);
  not (_40826_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_40828_, _40826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_40830_, _40801_, _40788_);
  not (_40832_, _40830_);
  or (_40834_, _40832_, _40798_);
  or (_40836_, _40834_, _40794_);
  and (_40838_, _40836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_40840_, _40838_, _40828_);
  or (_40842_, _40840_, _40822_);
  and (_40844_, _40842_, _40784_);
  and (_40846_, _40844_, _40824_);
  nor (_40848_, _40784_, _38642_);
  or (_40850_, _40848_, _40846_);
  and (_43054_, _40850_, _43100_);
  not (_40853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_40855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _40853_);
  nand (_40857_, _40793_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_40859_, _40830_, _40798_);
  or (_40861_, _40859_, _40857_);
  and (_40862_, _40861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_40863_, _40862_, _40855_);
  and (_40864_, _40743_, _38622_);
  or (_40865_, _40864_, _40863_);
  and (_40866_, _40865_, _40784_);
  nand (_40867_, _40864_, _31265_);
  and (_40868_, _40867_, _40866_);
  nor (_40869_, _40784_, _38672_);
  or (_40870_, _40869_, _40868_);
  and (_43056_, _40870_, _43100_);
  and (_40871_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_40872_, _40857_, _40834_);
  and (_40873_, _40872_, _40871_);
  and (_40874_, _40743_, _38751_);
  or (_40875_, _40874_, _40873_);
  and (_40876_, _40875_, _40784_);
  nand (_40877_, _40874_, _31265_);
  and (_40878_, _40877_, _40876_);
  nor (_40879_, _40784_, _38658_);
  or (_40880_, _40879_, _40878_);
  and (_43058_, _40880_, _43100_);
  and (_40881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40882_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40789_);
  nor (_40883_, _40882_, _40881_);
  and (_40884_, _40883_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_40885_, _40884_, _40788_);
  and (_40886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40887_, _40886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_40888_, _40887_);
  and (_40889_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40890_, _40889_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_40891_, _40890_);
  and (_40892_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40893_, _40892_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40894_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_40895_, _40894_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_40896_, _40895_, _40893_);
  and (_40897_, _40896_, _40891_);
  and (_40898_, _40897_, _40888_);
  not (_40899_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_40900_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_40901_, _40900_, _40899_);
  nand (_40902_, _40901_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_40903_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_40904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_40905_, _40904_, _40903_);
  and (_40906_, _40905_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_40907_, _40906_);
  and (_40908_, _40907_, _40902_);
  and (_40909_, _40908_, _40898_);
  nor (_40910_, _40909_, _40885_);
  and (_40911_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_40912_, _40911_, _40789_);
  and (_40913_, _40912_, _40910_);
  not (_40914_, _40913_);
  not (_40915_, _40912_);
  and (_40916_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _40788_);
  not (_40917_, _40916_);
  not (_40918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40919_, _40889_, _40918_);
  not (_40920_, _40919_);
  not (_40921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40922_, _40892_, _40921_);
  not (_40923_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_40924_, _40894_, _40923_);
  nor (_40925_, _40924_, _40922_);
  and (_40926_, _40925_, _40920_);
  nor (_40927_, _40926_, _40917_);
  not (_40928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40929_, _40901_, _40928_);
  not (_40930_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40931_, _40905_, _40930_);
  nor (_40932_, _40931_, _40929_);
  not (_40933_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40934_, _40886_, _40933_);
  not (_40935_, _40934_);
  and (_40936_, _40935_, _40932_);
  nor (_40937_, _40936_, _40917_);
  nor (_40938_, _40937_, _40927_);
  or (_40939_, _40938_, _40915_);
  and (_40940_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _43100_);
  and (_40941_, _40940_, _40939_);
  and (_43087_, _40941_, _40914_);
  nor (_40942_, _40911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40943_, _40942_);
  not (_40944_, _40910_);
  and (_40945_, _40938_, _40944_);
  nor (_40946_, _40945_, _40943_);
  nand (_40947_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _43100_);
  nor (_43089_, _40947_, _40946_);
  and (_40948_, _40908_, _40888_);
  nand (_40949_, _40948_, _40910_);
  or (_40950_, _40937_, _40910_);
  and (_40951_, _40950_, _40912_);
  and (_40952_, _40951_, _40949_);
  or (_40953_, _40952_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_40954_, _40914_, _40897_);
  nor (_40955_, _40915_, _40910_);
  nand (_40956_, _40955_, _40927_);
  and (_40957_, _40956_, _43100_);
  and (_40958_, _40957_, _40954_);
  and (_43091_, _40958_, _40953_);
  and (_40959_, _40949_, _40942_);
  or (_40960_, _40959_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40961_, _40942_, _40910_);
  not (_40962_, _40961_);
  or (_40963_, _40962_, _40897_);
  or (_40964_, _40937_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand (_40965_, _40942_, _40927_);
  and (_40966_, _40965_, _40964_);
  or (_40967_, _40966_, _40910_);
  and (_40968_, _40967_, _43100_);
  and (_40969_, _40968_, _40963_);
  and (_43093_, _40969_, _40960_);
  nand (_40970_, _40945_, _40788_);
  nor (_40971_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_40972_, _40971_, _40911_);
  and (_40973_, _40972_, _43100_);
  and (_43094_, _40973_, _40970_);
  and (_40974_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_40975_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_40976_, _40975_, _40971_);
  nor (_40977_, _40976_, _40944_);
  or (_40978_, _40977_, _40911_);
  or (_40984_, _40978_, _40974_);
  not (_40990_, _40911_);
  or (_40996_, _40976_, _40990_);
  and (_41002_, _40996_, _43100_);
  and (_43096_, _41002_, _40984_);
  and (_41006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _43100_);
  and (_43098_, _41006_, _40911_);
  nor (_43102_, _40785_, rst);
  and (_43104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _43100_);
  nor (_41007_, _40945_, _40911_);
  and (_41008_, _40911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_41009_, _41008_, _41007_);
  and (_00131_, _41009_, _43100_);
  and (_41010_, _40911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_41011_, _41010_, _41007_);
  and (_00133_, _41011_, _43100_);
  and (_41012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _43100_);
  and (_00135_, _41012_, _40911_);
  not (_41015_, _40924_);
  nor (_41019_, _40931_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_41023_, _41019_, _40929_);
  or (_41024_, _41023_, _40934_);
  and (_41025_, _41024_, _41015_);
  or (_41026_, _41025_, _40922_);
  nor (_41032_, _40938_, _40910_);
  and (_41036_, _41032_, _40920_);
  and (_41037_, _41036_, _41026_);
  not (_41039_, _40895_);
  or (_41040_, _40906_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_41046_, _41040_, _40902_);
  or (_41049_, _41046_, _40887_);
  and (_41050_, _41049_, _41039_);
  or (_41051_, _41050_, _40893_);
  and (_41057_, _40910_, _40891_);
  and (_41061_, _41057_, _41051_);
  or (_41062_, _41061_, _40911_);
  or (_41064_, _41062_, _41037_);
  or (_41065_, _40990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_41073_, _41065_, _43100_);
  and (_00137_, _41073_, _41064_);
  not (_41074_, _40893_);
  or (_41076_, _40895_, _40887_);
  and (_41082_, _40908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_41085_, _41082_, _41076_);
  and (_41086_, _41085_, _41074_);
  and (_41087_, _41086_, _41057_);
  nor (_41093_, _40922_, _40919_);
  or (_41097_, _40934_, _40924_);
  and (_41098_, _40932_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_41099_, _41098_, _41097_);
  and (_41105_, _41099_, _41093_);
  and (_41109_, _41105_, _41032_);
  or (_41110_, _41109_, _40911_);
  or (_41111_, _41110_, _41087_);
  or (_41113_, _40990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_41119_, _41113_, _43100_);
  and (_00139_, _41119_, _41111_);
  and (_41122_, _40935_, _40916_);
  nand (_41129_, _41122_, _40926_);
  nor (_41130_, _41129_, _40932_);
  nor (_41133_, _40908_, _40885_);
  or (_41134_, _41133_, _41130_);
  or (_41135_, _40898_, _40885_);
  and (_41141_, _41135_, _41134_);
  or (_41145_, _41141_, _40911_);
  or (_41146_, _40990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_41147_, _41146_, _43100_);
  and (_00140_, _41147_, _41145_);
  and (_41156_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _43100_);
  and (_00142_, _41156_, _40911_);
  and (_41157_, _40911_, _40789_);
  or (_41161_, _41157_, _40946_);
  or (_41167_, _41161_, _40955_);
  and (_00144_, _41167_, _43100_);
  not (_41168_, _41007_);
  and (_41172_, _41168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_41178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_41179_, _40906_, _40789_);
  or (_41180_, _41179_, _41178_);
  nor (_41183_, _40902_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_41189_, _41183_, _40887_);
  nand (_41191_, _41189_, _41180_);
  or (_41192_, _40888_, _40791_);
  and (_41195_, _41192_, _41191_);
  or (_41201_, _41195_, _40895_);
  or (_41202_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40789_);
  or (_41203_, _41202_, _41039_);
  and (_41204_, _41203_, _41074_);
  and (_41205_, _41204_, _41201_);
  and (_41206_, _40893_, _40791_);
  or (_41207_, _41206_, _40890_);
  or (_41208_, _41207_, _41205_);
  or (_41209_, _41202_, _40891_);
  and (_41210_, _41209_, _40910_);
  and (_41211_, _41210_, _41208_);
  and (_41212_, _40931_, _40789_);
  or (_41213_, _41212_, _41178_);
  and (_41214_, _40929_, _40789_);
  nor (_41215_, _41214_, _40934_);
  nand (_41216_, _41215_, _41213_);
  or (_41217_, _40935_, _40791_);
  and (_41218_, _41217_, _41216_);
  or (_41219_, _41218_, _40924_);
  not (_41220_, _40922_);
  or (_41221_, _41202_, _41015_);
  and (_41222_, _41221_, _41220_);
  and (_41223_, _41222_, _41219_);
  and (_41224_, _40922_, _40791_);
  or (_41225_, _41224_, _40919_);
  or (_41226_, _41225_, _41223_);
  and (_41227_, _41202_, _41032_);
  or (_41228_, _41227_, _41036_);
  and (_41229_, _41228_, _41226_);
  or (_41230_, _41229_, _41211_);
  and (_41231_, _41230_, _40990_);
  or (_41232_, _41231_, _41172_);
  and (_00146_, _41232_, _43100_);
  and (_41233_, _41168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_41234_, _41179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_41235_, _41234_, _41189_);
  and (_41236_, _40887_, _40800_);
  or (_41237_, _41236_, _41235_);
  and (_41238_, _41237_, _40896_);
  not (_41239_, _40896_);
  or (_41240_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40789_);
  and (_41241_, _41240_, _41239_);
  or (_41242_, _41241_, _40890_);
  or (_41243_, _41242_, _41238_);
  or (_41244_, _40891_, _40800_);
  and (_41245_, _41244_, _40910_);
  and (_41246_, _41245_, _41243_);
  and (_41247_, _40919_, _40800_);
  and (_41248_, _41240_, _40920_);
  or (_41249_, _41248_, _40926_);
  and (_41250_, _40934_, _40800_);
  not (_41251_, _40925_);
  or (_41252_, _41212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_41253_, _41252_, _41215_);
  or (_41254_, _41253_, _41251_);
  or (_41255_, _41254_, _41250_);
  and (_41256_, _41255_, _41249_);
  or (_41257_, _41256_, _41247_);
  and (_41258_, _41257_, _41032_);
  or (_41259_, _41258_, _41246_);
  and (_41260_, _41259_, _40990_);
  or (_41261_, _41260_, _41233_);
  and (_00148_, _41261_, _43100_);
  and (_41262_, _41168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_41263_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_41264_, _41263_, _40891_);
  and (_41265_, _41264_, _40910_);
  not (_41266_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_41267_, _40906_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_41268_, _41267_, _41266_);
  nor (_41269_, _40902_, _40789_);
  nor (_41270_, _41269_, _40887_);
  nand (_41271_, _41270_, _41268_);
  or (_41272_, _40888_, _40790_);
  and (_41273_, _41272_, _41271_);
  or (_41274_, _41273_, _40895_);
  or (_41275_, _41263_, _41039_);
  and (_41276_, _41275_, _41074_);
  and (_41277_, _41276_, _41274_);
  and (_41278_, _40893_, _40790_);
  or (_41279_, _41278_, _40890_);
  or (_41280_, _41279_, _41277_);
  and (_41281_, _41280_, _41265_);
  or (_41282_, _41263_, _40920_);
  and (_41283_, _40931_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_41284_, _41283_, _41266_);
  and (_41285_, _40929_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_41286_, _41285_, _40934_);
  nand (_41287_, _41286_, _41284_);
  or (_41288_, _40935_, _40790_);
  and (_41289_, _41288_, _41287_);
  or (_41290_, _41289_, _40924_);
  or (_41291_, _41263_, _41015_);
  and (_41292_, _41291_, _41220_);
  and (_41293_, _41292_, _41290_);
  and (_41294_, _40922_, _40790_);
  or (_41295_, _41294_, _40919_);
  or (_41296_, _41295_, _41293_);
  and (_41297_, _41296_, _41032_);
  and (_41298_, _41297_, _41282_);
  or (_41299_, _41298_, _41281_);
  and (_41300_, _41299_, _40990_);
  or (_41301_, _41300_, _41262_);
  and (_00150_, _41301_, _43100_);
  and (_41302_, _41168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_41303_, _41267_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_41304_, _41303_, _41270_);
  and (_41305_, _40887_, _40799_);
  or (_41306_, _41305_, _41304_);
  and (_41307_, _41306_, _40896_);
  or (_41308_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_41309_, _41308_, _41239_);
  or (_41310_, _41309_, _40890_);
  or (_41312_, _41310_, _41307_);
  or (_41313_, _40891_, _40799_);
  and (_41315_, _41313_, _40910_);
  and (_41316_, _41315_, _41312_);
  and (_41318_, _40919_, _40799_);
  and (_41319_, _41308_, _40920_);
  or (_41321_, _41319_, _40926_);
  and (_41322_, _40934_, _40799_);
  or (_41324_, _41283_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_41325_, _41324_, _41286_);
  or (_41327_, _41325_, _41251_);
  or (_41328_, _41327_, _41322_);
  and (_41330_, _41328_, _41321_);
  or (_41331_, _41330_, _41318_);
  and (_41333_, _41331_, _41032_);
  or (_41334_, _41333_, _41316_);
  and (_41336_, _41334_, _40990_);
  or (_41337_, _41336_, _41302_);
  and (_00151_, _41337_, _43100_);
  or (_41339_, _40943_, _40938_);
  and (_41340_, _41339_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_41341_, _41340_, _40961_);
  and (_00153_, _41341_, _43100_);
  and (_41342_, _40939_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_41343_, _41342_, _40913_);
  and (_00155_, _41343_, _43100_);
  and (_41344_, _40773_, _27003_);
  or (_41345_, _41344_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_41346_, _41345_, _40784_);
  nand (_41347_, _41344_, _31265_);
  and (_41348_, _41347_, _41346_);
  and (_41349_, _40770_, _38683_);
  or (_41350_, _41349_, _41348_);
  and (_00157_, _41350_, _43100_);
  and (_41351_, _40773_, _33344_);
  or (_41352_, _41351_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_41353_, _41352_, _40784_);
  nand (_41354_, _41351_, _31265_);
  and (_41355_, _41354_, _41353_);
  nor (_41356_, _40784_, _38665_);
  or (_41357_, _41356_, _41355_);
  and (_00159_, _41357_, _43100_);
  and (_41358_, _40773_, _34791_);
  or (_41359_, _41358_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_41360_, _41359_, _40784_);
  nand (_41361_, _41358_, _31265_);
  and (_41362_, _41361_, _41360_);
  nor (_41363_, _40784_, _38650_);
  or (_41364_, _41363_, _41362_);
  and (_00161_, _41364_, _43100_);
  and (_41365_, _40762_, _27003_);
  or (_41366_, _41365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_41367_, _41366_, _40759_);
  nand (_41368_, _41365_, _31265_);
  and (_41369_, _41368_, _41367_);
  and (_41370_, _40758_, _38683_);
  or (_41371_, _41370_, _41369_);
  and (_00162_, _41371_, _43100_);
  and (_41372_, _40762_, _32604_);
  or (_41373_, _41372_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_41374_, _41373_, _40759_);
  nand (_41375_, _41372_, _31265_);
  and (_41376_, _41375_, _41374_);
  nor (_41377_, _40759_, _38672_);
  or (_41378_, _41377_, _41376_);
  and (_00164_, _41378_, _43100_);
  nand (_41379_, _40762_, _39511_);
  and (_41380_, _41379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_41381_, _41380_, _40758_);
  and (_41382_, _33377_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_41383_, _41382_, _33366_);
  and (_41384_, _41383_, _40762_);
  or (_41385_, _41384_, _41381_);
  nand (_41386_, _40758_, _38665_);
  and (_41387_, _41386_, _43100_);
  and (_00166_, _41387_, _41385_);
  and (_41388_, _40762_, _34052_);
  or (_41389_, _41388_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_41390_, _41389_, _40759_);
  nand (_41391_, _41388_, _31265_);
  and (_41392_, _41391_, _41390_);
  nor (_41393_, _40759_, _38658_);
  or (_41394_, _41393_, _41392_);
  and (_00168_, _41394_, _43100_);
  and (_41395_, _40762_, _34791_);
  or (_41396_, _41395_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_41397_, _41396_, _40759_);
  nand (_41398_, _41395_, _31265_);
  and (_41399_, _41398_, _41397_);
  nor (_41400_, _40759_, _38650_);
  or (_41401_, _41400_, _41399_);
  and (_00170_, _41401_, _43100_);
  and (_41402_, _40762_, _35607_);
  or (_41403_, _41402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_41404_, _41403_, _40759_);
  nand (_41405_, _41402_, _31265_);
  and (_41406_, _41405_, _41404_);
  nor (_41407_, _40759_, _38642_);
  or (_41408_, _41407_, _41406_);
  and (_00172_, _41408_, _43100_);
  and (_41409_, _40762_, _36336_);
  or (_41410_, _41409_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_41411_, _41410_, _40759_);
  nand (_41412_, _41409_, _31265_);
  and (_41413_, _41412_, _41411_);
  nor (_41414_, _40759_, _38635_);
  or (_41415_, _41414_, _41413_);
  and (_00173_, _41415_, _43100_);
  and (_41416_, _40746_, _27003_);
  nand (_41417_, _41416_, _31265_);
  nor (_41418_, _41416_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_41419_, _41418_, _40750_);
  and (_41420_, _41419_, _41417_);
  and (_41421_, _40754_, _38683_);
  or (_41422_, _41421_, _41420_);
  and (_00175_, _41422_, _43100_);
  and (_41423_, _40746_, _32604_);
  nand (_41424_, _41423_, _31265_);
  nor (_41425_, _41423_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_41426_, _41425_, _40750_);
  and (_41427_, _41426_, _41424_);
  not (_41428_, _38672_);
  and (_41429_, _40754_, _41428_);
  or (_41430_, _41429_, _41427_);
  and (_00177_, _41430_, _43100_);
  and (_41431_, _33377_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_41432_, _41431_, _33366_);
  and (_41433_, _41432_, _40746_);
  nand (_41434_, _40746_, _39511_);
  and (_41435_, _41434_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_41436_, _41435_, _40750_);
  or (_41437_, _41436_, _41433_);
  nand (_41438_, _40750_, _38665_);
  and (_41439_, _41438_, _43100_);
  and (_00179_, _41439_, _41437_);
  and (_41440_, _40746_, _34052_);
  nand (_41441_, _41440_, _31265_);
  nor (_41442_, _41440_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor (_41443_, _41442_, _40750_);
  and (_41444_, _41443_, _41441_);
  and (_41445_, _40754_, _40346_);
  or (_41446_, _41445_, _41444_);
  and (_00181_, _41446_, _43100_);
  and (_41447_, _40746_, _34791_);
  nand (_41448_, _41447_, _31265_);
  nor (_41449_, _41447_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nor (_41450_, _41449_, _40750_);
  and (_41451_, _41450_, _41448_);
  and (_41452_, _40754_, _40357_);
  or (_41453_, _41452_, _41451_);
  and (_00183_, _41453_, _43100_);
  not (_41454_, _40750_);
  and (_41455_, _40746_, _35607_);
  and (_41456_, _41455_, _31265_);
  nor (_41457_, _41455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_41458_, _41457_, _41456_);
  nand (_41459_, _41458_, _41454_);
  nand (_41460_, _40750_, _38642_);
  and (_41461_, _41460_, _43100_);
  and (_00184_, _41461_, _41459_);
  and (_41462_, _40746_, _36336_);
  nand (_41463_, _41462_, _31265_);
  nor (_41464_, _41462_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nor (_41465_, _41464_, _40750_);
  and (_41466_, _41465_, _41463_);
  and (_41467_, _40754_, _40383_);
  or (_41468_, _41467_, _41466_);
  and (_00186_, _41468_, _43100_);
  and (_41469_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_41470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_41471_, _40785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_41472_, _41471_, _41470_);
  not (_41473_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_41474_, _41473_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_41475_, _41474_, _41472_);
  nor (_41476_, _41475_, _41469_);
  or (_41477_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_41478_, _41477_, _43100_);
  nor (_00546_, _41478_, _41476_);
  nor (_41479_, _41476_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_41480_, _41479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_41481_, _41479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_41482_, _41481_, _43100_);
  and (_00549_, _41482_, _41480_);
  not (_41483_, rxd_i);
  and (_41484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _41483_);
  nor (_41485_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_41486_, _41485_);
  and (_41487_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_41488_, _41487_, _41486_);
  and (_41489_, _41488_, _41484_);
  not (_41490_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_41491_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _41490_);
  and (_41492_, _41491_, _41485_);
  or (_41493_, _41492_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or (_41494_, _41493_, _41489_);
  and (_41495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _43100_);
  and (_00552_, _41495_, _41494_);
  and (_41496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_41497_, _41496_, _41486_);
  not (_41498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_41499_, _41485_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41500_, _41499_, _41498_);
  nor (_41501_, _41500_, _41497_);
  not (_41502_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_41503_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _41502_);
  not (_41504_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_41505_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _41504_);
  and (_41506_, _41505_, _41503_);
  not (_41507_, _41506_);
  or (_41508_, _41507_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and (_41509_, _41506_, _41497_);
  and (_41510_, _41497_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41511_, _41510_, _41509_);
  and (_41512_, _41511_, _41508_);
  or (_41513_, _41512_, _41501_);
  not (_41514_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand (_41515_, _41485_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_41516_, _41515_, _41514_);
  not (_41517_, _41516_);
  or (_41518_, _41517_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_41519_, _41518_, _41513_);
  nand (_00554_, _41519_, _41495_);
  not (_41520_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_41521_, _41497_);
  nor (_41522_, _41498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_41523_, _41522_);
  not (_41524_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41525_, _41485_, _41524_);
  and (_41526_, _41525_, _41523_);
  and (_41527_, _41526_, _41521_);
  nor (_41528_, _41527_, _41520_);
  and (_41529_, _41527_, rxd_i);
  or (_41530_, _41529_, rst);
  or (_00557_, _41530_, _41528_);
  nor (_41531_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41532_, _41531_, _41503_);
  and (_41533_, _41532_, _41510_);
  nand (_41534_, _41533_, _41483_);
  or (_41535_, _41533_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_41536_, _41535_, _43100_);
  and (_00560_, _41536_, _41534_);
  and (_41537_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41538_, _41537_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41539_, _41538_, _41502_);
  and (_41540_, _41539_, _41510_);
  and (_41541_, _41488_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41542_, _41541_, _41510_);
  nor (_41543_, _41538_, _41521_);
  or (_41544_, _41543_, _41542_);
  and (_41545_, _41544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_41546_, _41545_, _41540_);
  and (_00562_, _41546_, _43100_);
  and (_41547_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _43100_);
  nand (_41548_, _41547_, _41524_);
  nand (_41549_, _41495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand (_00565_, _41549_, _41548_);
  and (_41550_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41524_);
  not (_41551_, _41488_);
  nand (_41552_, _41492_, _41514_);
  and (_41553_, _41552_, _41551_);
  nand (_41554_, _41553_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand (_41555_, _41554_, _41521_);
  or (_41556_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_41557_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_41558_, _41557_, _41509_);
  and (_41559_, _41558_, _41556_);
  and (_41560_, _41559_, _41555_);
  or (_41561_, _41560_, _41516_);
  nand (_41562_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_41563_, _41562_, _41497_);
  or (_41564_, _41563_, _41507_);
  and (_41565_, _41564_, _41517_);
  or (_41566_, _41565_, rxd_i);
  and (_41567_, _41566_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41568_, _41567_, _41561_);
  or (_41569_, _41568_, _41550_);
  and (_00568_, _41569_, _43100_);
  and (_41570_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_41571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_41572_, _41471_, _41571_);
  or (_41573_, _41572_, _41474_);
  nor (_41574_, _41573_, _41570_);
  or (_41575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_41576_, _41575_, _43100_);
  nor (_00571_, _41576_, _41574_);
  nor (_41577_, _41574_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_41578_, _41577_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_41579_, _41577_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_41580_, _41579_, _43100_);
  and (_00573_, _41580_, _41578_);
  not (_41581_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_41582_, _32604_, _27661_);
  and (_41583_, _41582_, _30651_);
  and (_41584_, _41583_, _39442_);
  and (_41585_, _41584_, _43100_);
  nand (_41586_, _41585_, _41581_);
  not (_41587_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_41588_, _41515_, _41587_);
  nor (_41589_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not (_41590_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_41591_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_41592_, _41591_, _41590_);
  and (_41593_, _41592_, _41589_);
  not (_41594_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_41595_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_41596_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41597_, _41596_, _41595_);
  and (_41598_, _41597_, _41594_);
  and (_41599_, _41598_, _41593_);
  or (_41600_, _41599_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand (_41601_, _41599_, _41581_);
  nand (_41602_, _41601_, _41600_);
  nand (_41603_, _41602_, _41588_);
  nor (_41604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41605_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_41606_, _41605_, _41604_);
  and (_41607_, _41486_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_41608_, _41607_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_41609_, _41608_, _41606_);
  not (_41610_, _41609_);
  or (_41611_, _41610_, _41600_);
  and (_41612_, _41606_, _41607_);
  or (_41613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _41587_);
  or (_41614_, _41613_, _41612_);
  or (_41615_, _41614_, _41588_);
  and (_41616_, _41615_, _41611_);
  nand (_41617_, _41616_, _41603_);
  nor (_41618_, _41584_, rst);
  nand (_41619_, _41618_, _41617_);
  and (_00576_, _41619_, _41586_);
  not (_41620_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and (_41621_, _41599_, _41620_);
  nand (_41622_, _41612_, _41621_);
  and (_41623_, _41599_, _41588_);
  or (_41624_, _41587_, rst);
  nor (_41625_, _41624_, _41623_);
  and (_41626_, _41625_, _41622_);
  or (_00579_, _41626_, _41585_);
  or (_41627_, _41610_, _41621_);
  or (_41628_, _41612_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_41629_, _41515_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_41630_, _41629_, _41628_);
  and (_41631_, _41630_, _41627_);
  or (_41632_, _41631_, _41623_);
  and (_00581_, _41632_, _41618_);
  and (_41633_, _41608_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_41634_, _41633_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_41635_, _41634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or (_41636_, _41635_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_41637_, _41635_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_41638_, _41637_, _41636_);
  and (_00584_, _41638_, _41618_);
  nor (_41639_, _41609_, _41588_);
  and (_41640_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_41641_, _41640_, _41618_);
  and (_41642_, _41585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_00587_, _41642_, _41641_);
  and (_41643_, _40749_, _38620_);
  or (_41644_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_41645_, _41644_, _43100_);
  nand (_41646_, _41643_, _38704_);
  and (_00589_, _41646_, _41645_);
  and (_41647_, _40745_, _39420_);
  and (_41648_, _41647_, _31308_);
  nand (_41649_, _41648_, _31265_);
  and (_41650_, _40757_, _39442_);
  nor (_41651_, _41648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_41652_, _41651_, _41650_);
  and (_41653_, _41652_, _41649_);
  not (_41654_, _41650_);
  nor (_41655_, _41654_, _38704_);
  or (_41656_, _41655_, _41653_);
  and (_00592_, _41656_, _43100_);
  nor (_41657_, _41516_, _41509_);
  not (_41658_, _41657_);
  nor (_41659_, _41553_, _41497_);
  nor (_41660_, _41659_, _41658_);
  nor (_41661_, _41660_, _41524_);
  or (_41662_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_41663_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _41524_);
  or (_41664_, _41663_, _41657_);
  and (_41665_, _41664_, _43100_);
  and (_01211_, _41665_, _41662_);
  or (_41666_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_41667_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _41524_);
  or (_41668_, _41667_, _41657_);
  and (_41669_, _41668_, _43100_);
  and (_01213_, _41669_, _41666_);
  or (_41670_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_41671_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41524_);
  or (_41672_, _41671_, _41657_);
  and (_41673_, _41672_, _43100_);
  and (_01215_, _41673_, _41670_);
  or (_41674_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_41675_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41524_);
  or (_41676_, _41675_, _41657_);
  and (_41677_, _41676_, _43100_);
  and (_01217_, _41677_, _41674_);
  or (_41678_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_41679_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41524_);
  or (_41680_, _41679_, _41657_);
  and (_41681_, _41680_, _43100_);
  and (_01219_, _41681_, _41678_);
  or (_41682_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_41683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41524_);
  or (_41684_, _41683_, _41657_);
  and (_41685_, _41684_, _43100_);
  and (_01221_, _41685_, _41682_);
  or (_41686_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_41687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41524_);
  or (_41688_, _41687_, _41657_);
  and (_41689_, _41688_, _43100_);
  and (_01223_, _41689_, _41686_);
  or (_41690_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_41691_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _41524_);
  or (_41692_, _41691_, _41657_);
  and (_41693_, _41692_, _43100_);
  and (_01224_, _41693_, _41690_);
  nor (_41694_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_41695_, _41694_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_41696_, _41507_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or (_41697_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_41698_, _41697_, _41497_);
  and (_41699_, _41698_, _41696_);
  or (_41700_, _41488_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_41701_, _41700_, _41552_);
  and (_41702_, _41701_, _41521_);
  or (_41703_, _41702_, _41699_);
  or (_41704_, _41703_, _41516_);
  or (_41705_, _41517_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_41706_, _41705_, _41495_);
  and (_41707_, _41706_, _41704_);
  or (_01226_, _41707_, _41695_);
  and (_41708_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_41709_, _41708_, _41553_);
  or (_41710_, _41709_, _41660_);
  and (_41711_, _41710_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_41712_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _41524_);
  nand (_41713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41714_, _41713_, _41657_);
  or (_41715_, _41714_, _41712_);
  or (_41716_, _41715_, _41711_);
  and (_01228_, _41716_, _43100_);
  not (_41717_, _41661_);
  and (_41718_, _41717_, _41547_);
  or (_41719_, _41709_, _41658_);
  and (_41720_, _41495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_41721_, _41720_, _41719_);
  or (_01230_, _41721_, _41718_);
  or (_41722_, _41540_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_41723_, _41540_, _41483_);
  and (_41724_, _41723_, _43100_);
  and (_01232_, _41724_, _41722_);
  or (_41725_, _41542_, _41504_);
  or (_41726_, _41510_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41727_, _41726_, _43100_);
  and (_01234_, _41727_, _41725_);
  and (_41728_, _41542_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_41729_, _41531_, _41537_);
  and (_41730_, _41729_, _41510_);
  or (_41731_, _41730_, _41728_);
  and (_01236_, _41731_, _43100_);
  and (_41732_, _41544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41733_, _41537_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41734_, _41733_, _41543_);
  or (_41735_, _41734_, _41732_);
  and (_01238_, _41735_, _43100_);
  and (_41736_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41524_);
  and (_41737_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41738_, _41737_, _41736_);
  and (_01240_, _41738_, _43100_);
  and (_41739_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41524_);
  and (_41740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41741_, _41740_, _41739_);
  and (_01242_, _41741_, _43100_);
  and (_41742_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41524_);
  and (_41743_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41744_, _41743_, _41742_);
  and (_01244_, _41744_, _43100_);
  and (_41745_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41524_);
  and (_41746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41747_, _41746_, _41745_);
  and (_01246_, _41747_, _43100_);
  and (_41748_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41524_);
  and (_41749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41750_, _41749_, _41748_);
  and (_01248_, _41750_, _43100_);
  and (_41751_, _41495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_01250_, _41751_, _41695_);
  and (_41752_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41753_, _41752_, _41712_);
  and (_01252_, _41753_, _43100_);
  nor (_41754_, _41608_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41755_, _41754_, _41633_);
  and (_01254_, _41755_, _41618_);
  nor (_41756_, _41633_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_41757_, _41756_, _41634_);
  and (_01256_, _41757_, _41618_);
  nor (_41758_, _41634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_41759_, _41758_, _41635_);
  and (_01258_, _41759_, _41618_);
  and (_41760_, _41609_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_41761_, _41588_, _41620_);
  nor (_41762_, _41761_, _41609_);
  or (_41763_, _41762_, _41760_);
  and (_41764_, _41599_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41765_, _41764_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41766_, _41765_, _41588_);
  nor (_41767_, _41766_, _41763_);
  nor (_41768_, _41767_, _41584_);
  nor (_41769_, _41486_, _38682_);
  and (_41770_, _41769_, _41584_);
  or (_41771_, _41770_, _41768_);
  and (_01259_, _41771_, _43100_);
  not (_41772_, _41639_);
  and (_41773_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_41774_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_41775_, _41774_, _41773_);
  and (_41776_, _41775_, _41618_);
  nand (_41777_, _41485_, _38672_);
  nand (_41778_, _41486_, _38682_);
  and (_41779_, _41778_, _41585_);
  and (_41780_, _41779_, _41777_);
  or (_01261_, _41780_, _41776_);
  nor (_41781_, _41639_, _41594_);
  and (_41782_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or (_41783_, _41782_, _41781_);
  and (_41784_, _41783_, _41618_);
  nand (_41785_, _41485_, _38665_);
  nand (_41786_, _41486_, _38672_);
  and (_41787_, _41786_, _41585_);
  and (_41788_, _41787_, _41785_);
  or (_01263_, _41788_, _41784_);
  nor (_41789_, _41639_, _41590_);
  and (_41790_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or (_41791_, _41790_, _41789_);
  and (_41792_, _41791_, _41618_);
  nand (_41793_, _41486_, _38665_);
  nand (_41794_, _41485_, _38658_);
  and (_41795_, _41794_, _41585_);
  and (_41796_, _41795_, _41793_);
  or (_01265_, _41796_, _41792_);
  and (_41797_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41798_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or (_41799_, _41798_, _41797_);
  and (_41800_, _41799_, _41618_);
  nand (_41801_, _41485_, _38650_);
  nand (_41802_, _41486_, _38658_);
  and (_41803_, _41802_, _41585_);
  and (_41804_, _41803_, _41801_);
  or (_01267_, _41804_, _41800_);
  and (_41805_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_41806_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or (_41807_, _41806_, _41805_);
  and (_41808_, _41807_, _41618_);
  nand (_41809_, _41486_, _38650_);
  nand (_41810_, _41485_, _38642_);
  and (_41811_, _41810_, _41585_);
  and (_41812_, _41811_, _41809_);
  or (_01269_, _41812_, _41808_);
  and (_41813_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_41814_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or (_41815_, _41814_, _41813_);
  and (_41816_, _41815_, _41618_);
  nand (_41817_, _41485_, _38635_);
  nand (_41818_, _41486_, _38642_);
  and (_41819_, _41818_, _41585_);
  and (_41821_, _41819_, _41817_);
  or (_01271_, _41821_, _41816_);
  and (_41824_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_41826_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_41828_, _41826_, _41824_);
  and (_41830_, _41828_, _41618_);
  nand (_41832_, _41485_, _38704_);
  nand (_41834_, _41486_, _38635_);
  and (_41836_, _41834_, _41585_);
  and (_41838_, _41836_, _41832_);
  or (_01273_, _41838_, _41830_);
  and (_41841_, _41584_, _41486_);
  nand (_41843_, _41841_, _38704_);
  or (_41845_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_41847_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_41849_, _41847_, _41845_);
  or (_41851_, _41849_, _41584_);
  and (_41853_, _41851_, _43100_);
  and (_01275_, _41853_, _41843_);
  and (_41856_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_41858_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_41860_, _41858_, _41856_);
  and (_41862_, _41860_, _41618_);
  or (_41864_, _41473_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_41866_, _41864_, _41486_);
  and (_41868_, _41866_, _41585_);
  or (_01277_, _41868_, _41862_);
  nand (_41871_, _41643_, _38682_);
  or (_41873_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_41875_, _41873_, _43100_);
  and (_01279_, _41875_, _41871_);
  or (_41878_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_41880_, _41878_, _43100_);
  nand (_41882_, _41643_, _38672_);
  and (_01281_, _41882_, _41880_);
  or (_41884_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_41885_, _41884_, _43100_);
  nand (_41886_, _41643_, _38665_);
  and (_01283_, _41886_, _41885_);
  or (_41887_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_41888_, _41887_, _43100_);
  nand (_41889_, _41643_, _38658_);
  and (_01285_, _41889_, _41888_);
  or (_41890_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_41891_, _41890_, _43100_);
  nand (_41892_, _41643_, _38650_);
  and (_01287_, _41892_, _41891_);
  or (_41893_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_41894_, _41893_, _43100_);
  nand (_41895_, _41643_, _38642_);
  and (_01289_, _41895_, _41894_);
  or (_41896_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_41897_, _41896_, _43100_);
  nand (_41898_, _41643_, _38635_);
  and (_01291_, _41898_, _41897_);
  not (_41899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_41900_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41899_);
  or (_41901_, _41900_, _41485_);
  nor (_41902_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41903_, _41902_, _41901_);
  or (_41904_, _41903_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_41905_, _41904_, _41647_);
  or (_41906_, _27003_, _41490_);
  nand (_41907_, _41906_, _41647_);
  or (_41908_, _41907_, _39268_);
  and (_41909_, _41908_, _41905_);
  or (_41910_, _41909_, _41650_);
  nand (_41911_, _41650_, _38682_);
  and (_41912_, _41911_, _43100_);
  and (_01293_, _41912_, _41910_);
  or (_41913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_41914_, _41913_, _41647_);
  not (_41915_, _32604_);
  nor (_41916_, _41915_, _31265_);
  nand (_41917_, _41915_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_41918_, _41917_, _41647_);
  or (_41919_, _41918_, _41916_);
  and (_41920_, _41919_, _41914_);
  or (_41921_, _41920_, _41650_);
  nand (_41922_, _41650_, _38672_);
  and (_41923_, _41922_, _43100_);
  and (_01294_, _41923_, _41921_);
  not (_41924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not (_41925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_41926_, _41499_, _41925_);
  nor (_41927_, _41926_, _41924_);
  and (_41928_, _41926_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_41929_, _41928_, _41927_);
  or (_41930_, _41929_, _41647_);
  or (_41931_, _33344_, _41924_);
  nand (_41932_, _41931_, _41647_);
  or (_41933_, _41932_, _33366_);
  and (_41934_, _41933_, _41930_);
  or (_41935_, _41934_, _41650_);
  nand (_41936_, _41650_, _38665_);
  and (_41937_, _41936_, _43100_);
  and (_01296_, _41937_, _41935_);
  and (_41938_, _41647_, _34052_);
  nand (_41939_, _41938_, _31265_);
  nor (_41940_, _41938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor (_41941_, _41940_, _41650_);
  and (_41942_, _41941_, _41939_);
  nor (_41943_, _41654_, _38658_);
  or (_41944_, _41943_, _41942_);
  and (_01298_, _41944_, _43100_);
  and (_41945_, _41647_, _34791_);
  nand (_41946_, _41945_, _31265_);
  nor (_41947_, _41945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_41948_, _41947_, _41650_);
  and (_41949_, _41948_, _41946_);
  nor (_41950_, _41654_, _38650_);
  or (_41951_, _41950_, _41949_);
  and (_01300_, _41951_, _43100_);
  and (_41952_, _41647_, _35607_);
  nand (_41953_, _41952_, _31265_);
  nor (_41954_, _41952_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  nor (_41955_, _41954_, _41650_);
  and (_41956_, _41955_, _41953_);
  nor (_41957_, _41654_, _38642_);
  or (_41958_, _41957_, _41956_);
  and (_01302_, _41958_, _43100_);
  and (_41959_, _41647_, _36336_);
  nand (_41960_, _41959_, _31265_);
  nor (_41961_, _41959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nor (_41962_, _41961_, _41650_);
  and (_41963_, _41962_, _41960_);
  nor (_41964_, _41654_, _38635_);
  or (_41965_, _41964_, _41963_);
  and (_01304_, _41965_, _43100_);
  and (_01630_, t2_i, _43100_);
  nor (_41966_, t2_i, rst);
  and (_01633_, _41966_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand (_41967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _43100_);
  nor (_01636_, _41967_, t2ex_i);
  and (_01639_, t2ex_i, _43100_);
  and (_41968_, _38618_, _39112_);
  and (_41969_, _41968_, _40211_);
  nand (_41970_, _41969_, _38704_);
  and (_41971_, _40113_, _34052_);
  and (_41972_, _41968_, _41971_);
  not (_41973_, _41972_);
  and (_41974_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_41975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_41976_, _41975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41977_, _41976_, _41974_);
  not (_41978_, _41977_);
  and (_41979_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_41980_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_41981_, _41980_, _41979_);
  or (_41982_, _41969_, _41981_);
  and (_41983_, _41982_, _41973_);
  and (_41984_, _41983_, _41970_);
  and (_41985_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_41986_, _41985_, _41984_);
  and (_01642_, _41986_, _43100_);
  nand (_41987_, _41972_, _38704_);
  nor (_41988_, _41969_, _41978_);
  or (_41989_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_41990_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_41991_, _41988_, _41990_);
  and (_41992_, _41991_, _41989_);
  or (_41993_, _41992_, _41972_);
  and (_41994_, _41993_, _43100_);
  and (_01645_, _41994_, _41987_);
  and (_41995_, _41968_, _35607_);
  and (_41996_, _41995_, _40113_);
  and (_41997_, _41968_, _40172_);
  nor (_41998_, _41997_, _41996_);
  not (_41999_, _41975_);
  or (_42000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_42001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_42002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _42001_);
  and (_42003_, _42002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_42004_, _42003_, _42000_);
  and (_42005_, _42004_, _41999_);
  and (_42006_, _42005_, _41998_);
  and (_42007_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_42008_, _42007_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_42009_, _42008_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_42010_, _42009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_42011_, _42010_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_42012_, _42011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_42013_, _42012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_42014_, _42013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_42015_, _42014_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_42016_, _42015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_42017_, _42016_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_42018_, _42017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_42019_, _42018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_42020_, _42019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_42021_, _42020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_42022_, _42021_);
  nand (_42023_, _42022_, _42006_);
  or (_42024_, _42006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_42025_, _42024_, _43100_);
  and (_01648_, _42025_, _42023_);
  nand (_42026_, _41997_, _38704_);
  not (_42027_, _41996_);
  not (_42028_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_42029_, _41974_, _42028_);
  and (_42030_, _42029_, _41975_);
  and (_42031_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not (_42032_, _42030_);
  not (_42033_, _41976_);
  and (_42034_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_42035_, _42021_, _42004_);
  and (_42036_, _42035_, _42034_);
  and (_42037_, _42012_, _42004_);
  or (_42038_, _42037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_42039_, _42037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_42040_, _42039_, _42038_);
  or (_42041_, _42040_, _42036_);
  and (_42042_, _42041_, _42032_);
  or (_42043_, _42042_, _42031_);
  or (_42044_, _42043_, _41997_);
  and (_42045_, _42044_, _42027_);
  and (_42046_, _42045_, _42026_);
  and (_42047_, _41996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_42048_, _42047_, _42046_);
  and (_01651_, _42048_, _43100_);
  nand (_42049_, _41996_, _38704_);
  nor (_42050_, _42030_, _41990_);
  and (_42051_, _42032_, _42004_);
  and (_42052_, _42051_, _42020_);
  or (_42053_, _42052_, _42050_);
  nand (_42054_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand (_42055_, _42054_, _42035_);
  and (_42056_, _42055_, _42053_);
  nand (_42057_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand (_42058_, _42057_, _41998_);
  or (_42059_, _42058_, _42056_);
  nand (_42060_, _41997_, _41990_);
  and (_42061_, _42060_, _43100_);
  and (_42062_, _42061_, _42059_);
  and (_01654_, _42062_, _42049_);
  and (_42063_, _41975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_42064_, _42063_, _42052_);
  nand (_42065_, _42064_, _41998_);
  or (_42066_, _41998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_42067_, _42066_, _43100_);
  and (_01657_, _42067_, _42065_);
  or (_42068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_42069_, _40761_, _39096_);
  or (_42070_, _42069_, _42068_);
  nand (_42071_, _39099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_42072_, _42071_, _42069_);
  or (_42073_, _42072_, _39100_);
  and (_42074_, _42073_, _42070_);
  and (_42075_, _41968_, _40757_);
  or (_42076_, _42075_, _42074_);
  nand (_42077_, _42075_, _38704_);
  and (_42078_, _42077_, _43100_);
  and (_01660_, _42078_, _42076_);
  not (_42079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor (_42080_, _41977_, _42079_);
  and (_42081_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_42082_, _42081_, _42080_);
  or (_42083_, _42082_, _41969_);
  nand (_42084_, _41969_, _38682_);
  and (_42085_, _42084_, _42083_);
  or (_42086_, _42085_, _41972_);
  nand (_42087_, _41972_, _42079_);
  and (_42088_, _42087_, _43100_);
  and (_02112_, _42088_, _42086_);
  nand (_42089_, _41969_, _38672_);
  and (_42090_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_42091_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_42092_, _42091_, _42090_);
  or (_42093_, _42092_, _41969_);
  and (_42094_, _42093_, _41973_);
  and (_42095_, _42094_, _42089_);
  and (_42096_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_42097_, _42096_, _42095_);
  and (_02114_, _42097_, _43100_);
  nand (_42098_, _41969_, _38665_);
  and (_42099_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_42100_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_42101_, _42100_, _42099_);
  or (_42102_, _42101_, _41969_);
  and (_42103_, _42102_, _41973_);
  and (_42104_, _42103_, _42098_);
  and (_42105_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_42106_, _42105_, _42104_);
  and (_02116_, _42106_, _43100_);
  not (_42107_, _41969_);
  nor (_42108_, _42107_, _38658_);
  and (_42109_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_42110_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_42111_, _42110_, _42109_);
  nor (_42112_, _42111_, _41969_);
  or (_42113_, _42112_, _41972_);
  or (_42114_, _42113_, _42108_);
  or (_42115_, _41973_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_42116_, _42115_, _43100_);
  and (_02117_, _42116_, _42114_);
  nand (_42117_, _41969_, _38650_);
  and (_42118_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_42119_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_42120_, _42119_, _42118_);
  or (_42121_, _42120_, _41969_);
  and (_42122_, _42121_, _41973_);
  and (_42123_, _42122_, _42117_);
  and (_42124_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_42125_, _42124_, _42123_);
  and (_02119_, _42125_, _43100_);
  nand (_42126_, _41969_, _38642_);
  and (_42127_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_42128_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_42129_, _42128_, _42127_);
  or (_42130_, _42129_, _41969_);
  and (_42131_, _42130_, _41973_);
  and (_42132_, _42131_, _42126_);
  and (_42133_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_42134_, _42133_, _42132_);
  and (_02121_, _42134_, _43100_);
  nand (_42135_, _41969_, _38635_);
  and (_42136_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_42137_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_42138_, _42137_, _42136_);
  or (_42139_, _42138_, _41969_);
  and (_42140_, _42139_, _41973_);
  and (_42141_, _42140_, _42135_);
  and (_42142_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_42143_, _42142_, _42141_);
  and (_02123_, _42143_, _43100_);
  or (_42144_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_42145_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_42146_, _41988_, _42145_);
  and (_42147_, _42146_, _42144_);
  or (_42148_, _42147_, _41972_);
  nand (_42149_, _41972_, _38682_);
  and (_42150_, _42149_, _43100_);
  and (_02124_, _42150_, _42148_);
  not (_42151_, _41988_);
  and (_42152_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_42153_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_42154_, _42153_, _42152_);
  or (_42155_, _42154_, _41972_);
  nand (_42156_, _41972_, _38672_);
  and (_42157_, _42156_, _43100_);
  and (_02126_, _42157_, _42155_);
  nand (_42158_, _41972_, _38665_);
  and (_42159_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_42160_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_42161_, _42160_, _42159_);
  or (_42162_, _42161_, _41972_);
  and (_42163_, _42162_, _43100_);
  and (_02128_, _42163_, _42158_);
  nand (_42164_, _41972_, _38658_);
  and (_42165_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_42166_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_42167_, _42166_, _42165_);
  or (_42168_, _42167_, _41972_);
  and (_42169_, _42168_, _43100_);
  and (_02130_, _42169_, _42164_);
  nand (_42170_, _41972_, _38650_);
  and (_42171_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_42172_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_42173_, _42172_, _42171_);
  or (_42174_, _42173_, _41972_);
  and (_42175_, _42174_, _43100_);
  and (_02131_, _42175_, _42170_);
  nand (_42176_, _41972_, _38642_);
  and (_42177_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_42178_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_42179_, _42178_, _42177_);
  or (_42180_, _42179_, _41972_);
  and (_42181_, _42180_, _43100_);
  and (_02133_, _42181_, _42176_);
  nand (_42182_, _41972_, _38635_);
  and (_42183_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_42184_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_42185_, _42184_, _42183_);
  or (_42186_, _42185_, _41972_);
  and (_42187_, _42186_, _43100_);
  and (_02135_, _42187_, _42182_);
  and (_42188_, _42004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_42189_, _41976_, _42079_);
  nand (_42190_, _42189_, _42021_);
  nand (_42191_, _42190_, _42188_);
  or (_42192_, _42004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_42193_, _42192_, _42032_);
  and (_42194_, _42193_, _42191_);
  and (_42195_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_42196_, _42195_, _41997_);
  or (_42197_, _42196_, _42194_);
  and (_42198_, _41997_, _38682_);
  nor (_42199_, _42198_, _41996_);
  and (_42200_, _42199_, _42197_);
  and (_42201_, _41996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_42202_, _42201_, _42200_);
  and (_02137_, _42202_, _43100_);
  and (_42203_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_42204_, _42203_, _42051_);
  and (_42205_, _42204_, _42021_);
  and (_42206_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_42207_, _42188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_42208_, _42007_, _42004_);
  nor (_42209_, _42208_, _42030_);
  and (_42210_, _42209_, _42207_);
  nor (_42211_, _42210_, _42206_);
  nand (_42212_, _42211_, _41998_);
  or (_42213_, _42212_, _42205_);
  nand (_42214_, _41997_, _38672_);
  or (_42215_, _42027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_42216_, _42215_, _43100_);
  and (_42217_, _42216_, _42214_);
  and (_02138_, _42217_, _42213_);
  and (_42218_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_42219_, _42218_, _42035_);
  not (_42220_, _42208_);
  nor (_42221_, _42220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_42222_, _42220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_42223_, _42222_, _42221_);
  or (_42224_, _42223_, _42219_);
  and (_42225_, _42224_, _42032_);
  nand (_42226_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand (_42227_, _42226_, _41998_);
  or (_42228_, _42227_, _42225_);
  nand (_42229_, _41997_, _38665_);
  or (_42230_, _42027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_42231_, _42230_, _43100_);
  and (_42232_, _42231_, _42229_);
  and (_02140_, _42232_, _42228_);
  not (_42233_, _41997_);
  and (_42234_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_42235_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_42236_, _42235_, _42035_);
  nand (_42237_, _42008_, _42004_);
  nor (_42238_, _42237_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_42239_, _42237_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_42240_, _42239_, _42238_);
  or (_42241_, _42240_, _42236_);
  and (_42242_, _42241_, _42032_);
  or (_42243_, _42242_, _42234_);
  and (_42244_, _42243_, _42233_);
  nor (_42245_, _42233_, _38658_);
  or (_42246_, _42245_, _42244_);
  and (_42247_, _42246_, _42027_);
  and (_42248_, _41996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_42249_, _42248_, _42247_);
  and (_02142_, _42249_, _43100_);
  and (_42250_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_42251_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_42252_, _42251_, _42035_);
  nand (_42253_, _42009_, _42004_);
  nor (_42254_, _42253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_42255_, _42253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_42256_, _42255_, _42254_);
  or (_42257_, _42256_, _42252_);
  and (_42258_, _42257_, _42032_);
  or (_42259_, _42258_, _42250_);
  and (_42260_, _42259_, _42233_);
  nor (_42261_, _42233_, _38650_);
  or (_42262_, _42261_, _41996_);
  or (_42263_, _42262_, _42260_);
  or (_42264_, _42027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_42265_, _42264_, _43100_);
  and (_02144_, _42265_, _42263_);
  and (_42266_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_42267_, _42266_, _42035_);
  nand (_42268_, _42010_, _42004_);
  nor (_42269_, _42268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_42270_, _42268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_42271_, _42270_, _42269_);
  or (_42272_, _42271_, _42267_);
  and (_42273_, _42272_, _42032_);
  nand (_42274_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nand (_42275_, _42274_, _41998_);
  or (_42276_, _42275_, _42273_);
  nand (_42277_, _41997_, _38642_);
  or (_42278_, _42027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_42279_, _42278_, _43100_);
  and (_42280_, _42279_, _42277_);
  and (_02145_, _42280_, _42276_);
  nor (_42281_, _42233_, _38635_);
  and (_42282_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_42283_, _42282_, _42035_);
  and (_42284_, _42011_, _42004_);
  nor (_42285_, _42284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_42286_, _42285_, _42037_);
  or (_42287_, _42286_, _42030_);
  or (_42288_, _42287_, _42283_);
  or (_42289_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_42290_, _42289_, _41998_);
  and (_42291_, _42290_, _42288_);
  and (_42292_, _41996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_42293_, _42292_, _42291_);
  or (_42294_, _42293_, _42281_);
  and (_02147_, _42294_, _43100_);
  not (_42295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_42296_, _41976_, _42295_);
  and (_42297_, _42296_, _42035_);
  and (_42298_, _42013_, _42004_);
  or (_42299_, _42298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_42300_, _42298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_42301_, _42300_, _42299_);
  or (_42302_, _42301_, _42030_);
  or (_42303_, _42302_, _42297_);
  nand (_42304_, _42030_, _42295_);
  and (_42305_, _42304_, _41998_);
  and (_42306_, _42305_, _42303_);
  and (_42307_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_42308_, _41996_, _38683_);
  or (_42309_, _42308_, _42307_);
  or (_42310_, _42309_, _42306_);
  and (_02149_, _42310_, _43100_);
  and (_42311_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_42312_, _42311_, _42035_);
  and (_42313_, _42014_, _42004_);
  or (_42314_, _42313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_42315_, _42313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_42316_, _42315_, _42314_);
  or (_42317_, _42316_, _42030_);
  or (_42318_, _42317_, _42312_);
  not (_42319_, _41998_);
  nor (_42320_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_42321_, _42320_, _42319_);
  and (_42322_, _42321_, _42318_);
  and (_42323_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_42324_, _42027_, _38672_);
  or (_42325_, _42324_, _42323_);
  or (_42326_, _42325_, _42322_);
  and (_02151_, _42326_, _43100_);
  and (_42327_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_42328_, _42327_, _42035_);
  and (_42329_, _42015_, _42004_);
  or (_42330_, _42329_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand (_42331_, _42329_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_42332_, _42331_, _42330_);
  or (_42333_, _42332_, _42030_);
  or (_42334_, _42333_, _42328_);
  nor (_42335_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_42336_, _42335_, _42319_);
  and (_42337_, _42336_, _42334_);
  nor (_42338_, _42027_, _38665_);
  and (_42339_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_42340_, _42339_, _42338_);
  or (_42341_, _42340_, _42337_);
  and (_02152_, _42341_, _43100_);
  and (_42342_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_42343_, _42342_, _42035_);
  nand (_42344_, _42016_, _42004_);
  nor (_42345_, _42344_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_42346_, _42344_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_42347_, _42346_, _42030_);
  or (_42348_, _42347_, _42345_);
  or (_42349_, _42348_, _42343_);
  or (_42350_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_42351_, _42350_, _41998_);
  and (_42352_, _42351_, _42349_);
  and (_42353_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_42354_, _42353_, _42352_);
  nor (_42355_, _42027_, _38658_);
  or (_42356_, _42355_, _42354_);
  and (_02154_, _42356_, _43100_);
  and (_42357_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_42358_, _42357_, _42035_);
  nand (_42359_, _42017_, _42004_);
  nor (_42360_, _42359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_42361_, _42359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_42362_, _42361_, _42030_);
  or (_42363_, _42362_, _42360_);
  or (_42364_, _42363_, _42358_);
  or (_42365_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_42366_, _42365_, _41998_);
  and (_42367_, _42366_, _42364_);
  and (_42368_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_42369_, _42368_, _42367_);
  nor (_42370_, _42027_, _38650_);
  or (_42371_, _42370_, _42369_);
  and (_02156_, _42371_, _43100_);
  and (_42372_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_42373_, _42372_, _42035_);
  nand (_42374_, _42018_, _42004_);
  and (_42375_, _42374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_42376_, _42374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_42377_, _42376_, _42030_);
  or (_42378_, _42377_, _42375_);
  or (_42379_, _42378_, _42373_);
  or (_42380_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_42381_, _42380_, _41998_);
  and (_42382_, _42381_, _42379_);
  and (_42383_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_42384_, _42027_, _38642_);
  or (_42385_, _42384_, _42383_);
  or (_42386_, _42385_, _42382_);
  and (_02158_, _42386_, _43100_);
  and (_42387_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_42388_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_42389_, _42388_, _42035_);
  nand (_42390_, _42019_, _42004_);
  and (_42391_, _42390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_42392_, _42390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_42393_, _42392_, _42030_);
  or (_42394_, _42393_, _42391_);
  or (_42395_, _42394_, _42389_);
  or (_42396_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_42397_, _42396_, _41998_);
  and (_42398_, _42397_, _42395_);
  or (_42399_, _42398_, _42387_);
  nor (_42400_, _42027_, _38635_);
  or (_42401_, _42400_, _42399_);
  and (_02159_, _42401_, _43100_);
  not (_42402_, _42075_);
  and (_42403_, _42069_, _27003_);
  or (_42404_, _42403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_42405_, _42404_, _42402_);
  nand (_42406_, _42403_, _31265_);
  and (_42407_, _42406_, _42405_);
  and (_42408_, _42075_, _38683_);
  or (_42409_, _42408_, _42407_);
  and (_02161_, _42409_, _43100_);
  and (_42410_, _42069_, _32604_);
  or (_42411_, _42410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_42412_, _42411_, _42402_);
  nand (_42413_, _42410_, _31265_);
  and (_42414_, _42413_, _42412_);
  nor (_42415_, _42402_, _38672_);
  or (_42416_, _42415_, _42414_);
  and (_02163_, _42416_, _43100_);
  nand (_42417_, _42069_, _39511_);
  and (_42418_, _42417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_42419_, _42418_, _42075_);
  and (_42420_, _33377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_42421_, _42420_, _33366_);
  and (_42422_, _42421_, _42069_);
  or (_42423_, _42422_, _42419_);
  nand (_42424_, _42075_, _38665_);
  and (_42425_, _42424_, _43100_);
  and (_02165_, _42425_, _42423_);
  and (_42426_, _42069_, _34052_);
  or (_42427_, _42426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_42428_, _42427_, _42402_);
  nand (_42429_, _42426_, _31265_);
  and (_42430_, _42429_, _42428_);
  nor (_42431_, _42402_, _38658_);
  or (_42432_, _42431_, _42430_);
  and (_02166_, _42432_, _43100_);
  and (_42433_, _42069_, _34791_);
  or (_42434_, _42433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_42435_, _42434_, _42402_);
  nand (_42436_, _42433_, _31265_);
  and (_42437_, _42436_, _42435_);
  nor (_42438_, _42402_, _38650_);
  or (_42439_, _42438_, _42437_);
  and (_02167_, _42439_, _43100_);
  and (_42440_, _42069_, _35607_);
  or (_42441_, _42440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_42442_, _42441_, _42402_);
  nand (_42443_, _42440_, _31265_);
  and (_42444_, _42443_, _42442_);
  nor (_42445_, _42402_, _38642_);
  or (_42446_, _42445_, _42444_);
  and (_02168_, _42446_, _43100_);
  not (_42447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_42448_, _41974_, _42447_);
  or (_42449_, _42448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_42450_, _42449_, _42069_);
  nand (_42451_, _39221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_42452_, _42451_, _42069_);
  or (_42453_, _42452_, _39222_);
  and (_42454_, _42453_, _42450_);
  or (_42455_, _42454_, _42075_);
  nand (_42456_, _42075_, _38635_);
  and (_42457_, _42456_, _43100_);
  and (_02169_, _42457_, _42455_);
  nor (_42458_, _27496_, _26476_);
  nor (_42459_, _42458_, _30629_);
  and (_42460_, _38706_, _38615_);
  not (_42461_, _42460_);
  not (_42462_, _38614_);
  and (_42463_, _42462_, _38577_);
  nand (_42464_, _38006_, _26981_);
  or (_42465_, _38006_, _26981_);
  not (_42466_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_42467_, _30618_, _42466_);
  and (_42468_, _42467_, _33377_);
  and (_42469_, _42468_, _27496_);
  and (_42470_, _42469_, _42465_);
  and (_42471_, _42470_, _42464_);
  and (_42472_, _39111_, _39112_);
  and (_42473_, _42472_, _39113_);
  not (_42474_, _42473_);
  and (_42475_, _42474_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_42476_, _42475_, _39168_);
  and (_42477_, _42476_, _27661_);
  nor (_42478_, _42476_, _27661_);
  nor (_42479_, _42478_, _42477_);
  and (_42480_, _42479_, _42471_);
  not (_42481_, _42480_);
  and (_42482_, _42476_, _38479_);
  and (_42483_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_42484_, _42476_, _38006_);
  and (_42485_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_42486_, _42485_, _42483_);
  nor (_42487_, _42476_, _38479_);
  and (_42488_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_42489_, _42476_, _38006_);
  and (_42490_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_42491_, _42490_, _42488_);
  and (_42492_, _42491_, _42486_);
  and (_42493_, _42492_, _42481_);
  and (_42494_, _42480_, _38704_);
  nor (_42495_, _42494_, _42493_);
  and (_42496_, _42495_, _42463_);
  not (_42497_, _42496_);
  not (_42498_, _38477_);
  nor (_42499_, _42462_, _38577_);
  not (_42500_, _36509_);
  and (_42501_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_42502_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_42503_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_42504_, _42503_, _42502_);
  and (_42505_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_42506_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_42507_, _42506_, _42505_);
  and (_42508_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_42509_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_42510_, _42509_, _42508_);
  and (_42511_, _42510_, _42507_);
  and (_42512_, _42511_, _42504_);
  and (_42513_, _38017_, _36509_);
  not (_42514_, _42513_);
  nor (_42515_, _42514_, _42512_);
  nor (_42516_, _42515_, _42501_);
  not (_42517_, _42516_);
  and (_42518_, _42517_, _42499_);
  nor (_42519_, _42518_, _42498_);
  and (_42520_, _42519_, _42497_);
  and (_42521_, _42520_, _42461_);
  not (_42522_, _38550_);
  and (_42523_, _42522_, _38544_);
  nor (_42524_, _38539_, _38535_);
  nor (_42525_, _38547_, _38532_);
  and (_42526_, _42525_, _42524_);
  and (_42527_, _38561_, _38523_);
  and (_42528_, _42527_, _42526_);
  and (_42529_, _42528_, _42523_);
  nor (_42530_, _42529_, _36466_);
  nor (_42531_, _38559_, _38555_);
  not (_42532_, _38466_);
  nor (_42533_, _42532_, _42531_);
  nor (_42534_, _42533_, _42530_);
  not (_42535_, _42534_);
  and (_42536_, _42535_, _42521_);
  and (_42537_, _42499_, _38477_);
  and (_42538_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_42539_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_42540_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_42541_, _42540_, _42539_);
  and (_42542_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_42543_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_42544_, _42543_, _42542_);
  and (_42545_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_42546_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_42547_, _42546_, _42545_);
  and (_42548_, _42547_, _42544_);
  and (_42549_, _42548_, _42541_);
  nor (_42550_, _42549_, _42514_);
  nor (_42551_, _42550_, _42538_);
  not (_42552_, _42551_);
  and (_42553_, _42552_, _42537_);
  not (_42554_, _42553_);
  and (_42555_, _42498_, _38614_);
  and (_42556_, _38614_, _38577_);
  and (_42557_, _42556_, _38477_);
  and (_42558_, _42474_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_42559_, _42558_, _39181_);
  and (_42560_, _42559_, _42557_);
  nor (_42561_, _42560_, _42555_);
  and (_42562_, _42561_, _42554_);
  not (_42563_, _38738_);
  and (_42564_, _42563_, _38616_);
  and (_42565_, _42463_, _38477_);
  and (_42566_, _42480_, _40357_);
  and (_42567_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_42568_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_42569_, _42568_, _42567_);
  and (_42570_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_42571_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_42572_, _42571_, _42570_);
  and (_42573_, _42572_, _42569_);
  nor (_42574_, _42573_, _42480_);
  nor (_42575_, _42574_, _42566_);
  not (_42576_, _42575_);
  and (_42577_, _42576_, _42565_);
  nor (_42578_, _42577_, _42564_);
  and (_42579_, _42578_, _42562_);
  not (_42580_, _42579_);
  and (_42581_, _42580_, _42536_);
  and (_42582_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_42583_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_42584_, _42583_, _42582_);
  and (_42585_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_42586_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_42587_, _42586_, _42585_);
  and (_42588_, _42587_, _42584_);
  nor (_42589_, _42588_, _42480_);
  and (_42590_, _42480_, _41428_);
  nor (_42591_, _42590_, _42589_);
  not (_42592_, _42591_);
  and (_42593_, _42592_, _42565_);
  and (_42594_, _42463_, _42498_);
  not (_42595_, _38720_);
  and (_42596_, _42595_, _38616_);
  or (_42597_, _42596_, _42594_);
  and (_42598_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_42599_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_42600_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_42601_, _42600_, _42599_);
  and (_42602_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_42603_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_42604_, _42603_, _42602_);
  and (_42605_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_42606_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_42607_, _42606_, _42605_);
  and (_42608_, _42607_, _42604_);
  and (_42609_, _42608_, _42601_);
  nor (_42610_, _42609_, _42514_);
  nor (_42611_, _42610_, _42598_);
  not (_42612_, _42611_);
  and (_42613_, _42612_, _42537_);
  and (_42614_, _42557_, _38270_);
  or (_42615_, _42614_, _42613_);
  or (_42616_, _42615_, _42597_);
  nor (_42617_, _42616_, _42593_);
  nor (_42618_, _42617_, _42535_);
  nor (_42619_, _42618_, _42581_);
  and (_42620_, _27496_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42621_, _42620_, _40742_);
  nor (_42622_, _26860_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42623_, _42622_, _42621_);
  nand (_42624_, _42623_, _42619_);
  or (_42625_, _42623_, _42619_);
  and (_42626_, _42625_, _42624_);
  and (_42627_, _42620_, _27661_);
  nor (_42628_, _26981_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42629_, _42628_, _42627_);
  not (_42630_, _42629_);
  not (_42631_, _42476_);
  and (_42632_, _42557_, _42631_);
  and (_42633_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_42634_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_42635_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_42636_, _42635_, _42634_);
  and (_42637_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_42638_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_42639_, _42638_, _42637_);
  and (_42640_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_42641_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_42642_, _42641_, _42640_);
  and (_42643_, _42642_, _42639_);
  and (_42644_, _42643_, _42636_);
  nor (_42645_, _42644_, _42514_);
  nor (_42646_, _42645_, _42633_);
  not (_42647_, _42646_);
  and (_42648_, _42647_, _42537_);
  nor (_42649_, _42648_, _42632_);
  not (_42650_, _38732_);
  and (_42651_, _42650_, _38616_);
  and (_42652_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_42653_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_42654_, _42653_, _42652_);
  and (_42655_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_42656_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_42657_, _42656_, _42655_);
  and (_42658_, _42657_, _42654_);
  nor (_42659_, _42658_, _42480_);
  and (_42660_, _42480_, _40346_);
  nor (_42661_, _42660_, _42659_);
  not (_42662_, _42661_);
  and (_42663_, _42662_, _42565_);
  nor (_42664_, _42663_, _42651_);
  and (_42665_, _42664_, _42649_);
  not (_42666_, _42665_);
  and (_42667_, _42666_, _42536_);
  and (_42668_, _42557_, _38006_);
  and (_42669_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_42670_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_42671_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_42672_, _42671_, _42670_);
  and (_42673_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_42674_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_42675_, _42674_, _42673_);
  and (_42676_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_42677_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_42678_, _42677_, _42676_);
  and (_42679_, _42678_, _42675_);
  and (_42680_, _42679_, _42672_);
  nor (_42681_, _42680_, _42514_);
  nor (_42682_, _42681_, _42669_);
  not (_42683_, _42682_);
  and (_42684_, _42683_, _42537_);
  nor (_42685_, _42684_, _42668_);
  not (_42686_, _38714_);
  and (_42687_, _42686_, _38616_);
  and (_42688_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_42689_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_42690_, _42689_, _42688_);
  and (_42691_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_42692_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_42693_, _42692_, _42691_);
  and (_42694_, _42693_, _42690_);
  nor (_42695_, _42694_, _42480_);
  and (_42696_, _42480_, _38683_);
  nor (_42697_, _42696_, _42695_);
  not (_42698_, _42697_);
  and (_42699_, _42698_, _42565_);
  nor (_42700_, _42699_, _42687_);
  and (_42701_, _42700_, _42685_);
  nor (_42702_, _42701_, _42535_);
  nor (_42703_, _42702_, _42667_);
  and (_42704_, _42703_, _42630_);
  nor (_42705_, _42703_, _42630_);
  nor (_42706_, _42705_, _42704_);
  not (_42707_, _42706_);
  nor (_42708_, _42707_, _42626_);
  nor (_42709_, _42666_, _42536_);
  nor (_42710_, _42463_, _38477_);
  and (_42711_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_42712_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_42713_, _42712_, _42711_);
  and (_42714_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_42715_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_42716_, _42715_, _42714_);
  and (_42717_, _42716_, _42713_);
  nor (_42718_, _42717_, _42480_);
  and (_42719_, _42480_, _40383_);
  nor (_42720_, _42719_, _42718_);
  not (_42721_, _42720_);
  and (_42722_, _42721_, _42565_);
  nor (_42723_, _42722_, _42710_);
  not (_42724_, _38750_);
  and (_42725_, _42724_, _38616_);
  and (_42726_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_42727_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_42728_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_42729_, _42728_, _42727_);
  and (_42730_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_42731_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_42732_, _42731_, _42730_);
  and (_42733_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_42734_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_42735_, _42734_, _42733_);
  and (_42736_, _42735_, _42732_);
  and (_42737_, _42736_, _42729_);
  nor (_42738_, _42737_, _42514_);
  nor (_42739_, _42738_, _42726_);
  not (_42740_, _42739_);
  and (_42741_, _42740_, _42537_);
  nor (_42742_, _42741_, _42725_);
  and (_42743_, _42742_, _42723_);
  and (_42744_, _42743_, _42536_);
  nor (_42745_, _42744_, _42709_);
  nor (_42746_, _42620_, _27661_);
  and (_42747_, _42620_, _27211_);
  nor (_42748_, _42747_, _42746_);
  not (_42749_, _42748_);
  and (_42750_, _42749_, _42745_);
  nor (_42751_, _42749_, _42745_);
  nor (_42752_, _42751_, _42750_);
  and (_42753_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_42754_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_42755_, _42754_, _42753_);
  and (_42756_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_42757_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_42758_, _42757_, _42756_);
  and (_42759_, _42758_, _42755_);
  and (_42760_, _42759_, _42481_);
  and (_42761_, _42480_, _38642_);
  nor (_42762_, _42761_, _42760_);
  and (_42763_, _42762_, _42565_);
  and (_42764_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_42765_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_42766_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_42767_, _42766_, _42765_);
  and (_42768_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_42769_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_42770_, _42769_, _42768_);
  and (_42771_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_42772_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_42773_, _42772_, _42771_);
  and (_42774_, _42773_, _42770_);
  and (_42775_, _42774_, _42767_);
  nor (_42776_, _42775_, _42514_);
  nor (_42777_, _42776_, _42764_);
  not (_42778_, _42777_);
  and (_42779_, _42778_, _42537_);
  nor (_42780_, _42779_, _42763_);
  nor (_42781_, _38744_, _38614_);
  nor (_42782_, _42781_, _42498_);
  or (_42783_, _42556_, _38615_);
  not (_42784_, _42783_);
  nor (_42785_, _42784_, _42782_);
  not (_42786_, _42785_);
  and (_42787_, _42786_, _42780_);
  not (_42788_, _42787_);
  and (_42789_, _42788_, _42536_);
  and (_42790_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_42791_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_42792_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_42793_, _42792_, _42791_);
  and (_42794_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_42795_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_42796_, _42795_, _42794_);
  and (_42797_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_42798_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_42799_, _42798_, _42797_);
  and (_42800_, _42799_, _42796_);
  and (_42801_, _42800_, _42793_);
  nor (_42802_, _42801_, _42514_);
  nor (_42803_, _42802_, _42790_);
  not (_42804_, _42803_);
  and (_42805_, _42804_, _42537_);
  and (_42806_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_42807_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_42808_, _42807_, _42806_);
  and (_42809_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_42810_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_42811_, _42810_, _42809_);
  and (_42812_, _42811_, _42808_);
  nor (_42813_, _42812_, _42480_);
  and (_42814_, _42480_, _40334_);
  nor (_42815_, _42814_, _42813_);
  not (_42816_, _42815_);
  and (_42817_, _42816_, _42565_);
  nor (_42818_, _42817_, _42805_);
  not (_42819_, _38726_);
  and (_42820_, _42819_, _38616_);
  and (_42821_, _42557_, _38414_);
  nor (_42822_, _42821_, _42820_);
  and (_42823_, _42822_, _42818_);
  nor (_42824_, _42823_, _42535_);
  nor (_42825_, _42824_, _42789_);
  and (_42826_, _42620_, _39095_);
  nor (_42827_, _26740_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42828_, _42827_, _42826_);
  not (_42829_, _42828_);
  nor (_42830_, _42829_, _42825_);
  and (_42831_, _42829_, _42825_);
  nor (_42832_, _42831_, _42830_);
  and (_42833_, _42832_, _42752_);
  and (_42834_, _42833_, _42708_);
  and (_42835_, _42834_, _42459_);
  nor (_42836_, _42788_, _42536_);
  nor (_42837_, _42620_, _39095_);
  not (_42838_, _42837_);
  nor (_42839_, _42838_, _42836_);
  and (_42840_, _42838_, _42836_);
  nor (_42841_, _42840_, _42839_);
  nor (_42842_, _42579_, _42536_);
  nor (_42843_, _42620_, _27825_);
  not (_42844_, _42843_);
  nor (_42845_, _42844_, _42842_);
  and (_42846_, _42844_, _42842_);
  nor (_42847_, _42846_, _42845_);
  and (_42848_, _42847_, _42841_);
  nor (_42849_, _42743_, _42536_);
  nor (_42850_, _42620_, _27211_);
  not (_42851_, _42850_);
  nor (_42852_, _42851_, _42849_);
  and (_42853_, _42851_, _42849_);
  nor (_42854_, _42853_, _42852_);
  nor (_42855_, _42521_, _27496_);
  and (_42856_, _42521_, _27496_);
  nor (_42857_, _42856_, _42855_);
  not (_42858_, _42857_);
  and (_42859_, _42858_, _42854_);
  and (_42860_, _42859_, _42848_);
  and (_42861_, _42860_, _42835_);
  not (_42862_, _42825_);
  not (_42863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_42864_, _42703_, _42863_);
  and (_42865_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_42866_, _42865_, _42619_);
  or (_42867_, _42866_, _42864_);
  and (_42868_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_42869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_42870_, _42703_, _42869_);
  nand (_42871_, _42870_, _42619_);
  or (_42872_, _42871_, _42868_);
  and (_42873_, _42872_, _42867_);
  or (_42874_, _42873_, _42862_);
  not (_42875_, _42745_);
  not (_42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_42877_, _42703_, _42876_);
  and (_42878_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_42879_, _42878_, _42619_);
  or (_42880_, _42879_, _42877_);
  and (_42881_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not (_42882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_42883_, _42703_, _42882_);
  nand (_42884_, _42883_, _42619_);
  or (_42885_, _42884_, _42881_);
  and (_42886_, _42885_, _42880_);
  or (_42887_, _42886_, _42825_);
  and (_42888_, _42887_, _42875_);
  and (_42889_, _42888_, _42874_);
  not (_42890_, _42619_);
  not (_42891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_42892_, _42703_, _42891_);
  or (_42893_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_42894_, _42893_, _42892_);
  or (_42895_, _42894_, _42890_);
  or (_42896_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_42897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_42898_, _42703_, _42897_);
  and (_42899_, _42898_, _42896_);
  or (_42900_, _42899_, _42619_);
  and (_42901_, _42900_, _42895_);
  or (_42902_, _42901_, _42862_);
  not (_42903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_42904_, _42703_, _42903_);
  or (_42905_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_42906_, _42905_, _42904_);
  or (_42907_, _42906_, _42890_);
  or (_42908_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_42909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_42910_, _42703_, _42909_);
  and (_42911_, _42910_, _42908_);
  or (_42912_, _42911_, _42619_);
  and (_42913_, _42912_, _42907_);
  or (_42914_, _42913_, _42825_);
  and (_42915_, _42914_, _42745_);
  and (_42916_, _42915_, _42902_);
  or (_42917_, _42916_, _42889_);
  or (_42918_, _42917_, _42861_);
  not (_42919_, _42861_);
  or (_42920_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_42921_, _42835_);
  nor (_42922_, _42861_, _42921_);
  nor (_42923_, _42922_, rst);
  and (_42924_, _42923_, _42920_);
  and (_42925_, _42924_, _42918_);
  and (_42926_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_42927_, _42926_, _28659_);
  nor (_42928_, _42927_, _31265_);
  nand (_42929_, _28659_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42930_, _20043_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42931_, _42930_, _42929_);
  nor (_42932_, _38704_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_42933_, _42932_, _42931_);
  or (_42934_, _42933_, _42928_);
  and (_40239_, _42934_, _43100_);
  and (_42935_, _40239_, _42922_);
  or (_02567_, _42935_, _42925_);
  not (_42936_, _42459_);
  nor (_42937_, _42629_, _42936_);
  nor (_42938_, _42936_, _42623_);
  and (_42939_, _42938_, _42937_);
  and (_42940_, _42748_, _42459_);
  nor (_42941_, _42936_, _42828_);
  and (_42942_, _42941_, _42940_);
  and (_42943_, _42942_, _42939_);
  and (_42944_, _42934_, _42459_);
  and (_42945_, _42944_, _42943_);
  not (_42946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_42947_, _42943_, _42946_);
  or (_02578_, _42947_, _42945_);
  nor (_42948_, _42941_, _42940_);
  nor (_42949_, _42938_, _42937_);
  and (_42950_, _42949_, _42459_);
  and (_42951_, _42950_, _42948_);
  and (_42952_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _28648_);
  and (_42953_, _42952_, _28692_);
  nand (_42954_, _42953_, _31265_);
  not (_42955_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42956_, _38682_, _42955_);
  or (_42957_, _18880_, _42955_);
  and (_42958_, _42957_, _42956_);
  or (_42959_, _42958_, _42953_);
  and (_42960_, _42959_, _42954_);
  and (_42961_, _42960_, _42951_);
  not (_42962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_42963_, _42951_, _42962_);
  or (_02802_, _42963_, _42961_);
  not (_42964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_42965_, _42951_, _42964_);
  nand (_42966_, _42952_, _28736_);
  nor (_42967_, _42966_, _31265_);
  nor (_42968_, _38672_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42969_, _42952_, _28757_);
  and (_42970_, _42952_, _28659_);
  or (_42971_, _42970_, _42926_);
  or (_42972_, _42971_, _42969_);
  and (_42973_, _42972_, _19874_);
  or (_42974_, _42973_, _42968_);
  or (_42975_, _42974_, _42967_);
  and (_42976_, _42975_, _42951_);
  or (_02807_, _42976_, _42965_);
  not (_42977_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_42978_, _42951_, _42977_);
  nand (_42979_, _42952_, _28768_);
  nor (_42980_, _42979_, _31265_);
  nor (_42981_, _38665_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42982_, _42952_, _28725_);
  or (_42983_, _42982_, _42971_);
  and (_42984_, _42983_, _18518_);
  or (_42985_, _42984_, _42981_);
  or (_42986_, _42985_, _42980_);
  and (_42987_, _42986_, _42951_);
  or (_02812_, _42987_, _42978_);
  and (_42988_, _42970_, _31885_);
  nor (_42989_, _38658_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_42990_, _42969_, _42926_);
  or (_42991_, _42990_, _42982_);
  and (_42992_, _42991_, _19547_);
  or (_42993_, _42992_, _42989_);
  or (_42994_, _42993_, _42988_);
  and (_42995_, _42994_, _42951_);
  not (_42996_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_42997_, _42951_, _42996_);
  or (_02817_, _42997_, _42995_);
  nand (_42998_, _42926_, _28692_);
  nor (_42999_, _42998_, _31265_);
  nor (_43000_, _38650_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_43001_, _28692_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_43002_, _18716_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_43003_, _43002_, _43001_);
  or (_43004_, _43003_, _43000_);
  or (_43005_, _43004_, _42999_);
  and (_43006_, _43005_, _42951_);
  not (_43007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_43008_, _42951_, _43007_);
  or (_02822_, _43008_, _43006_);
  nand (_43009_, _42926_, _28736_);
  nor (_43010_, _43009_, _31265_);
  nor (_43011_, _38642_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_43012_, _28736_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_43013_, _19699_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_43014_, _43013_, _43012_);
  or (_43015_, _43014_, _43011_);
  or (_43016_, _43015_, _43010_);
  and (_43017_, _43016_, _42951_);
  not (_43018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_43019_, _42951_, _43018_);
  or (_02827_, _43019_, _43017_);
  nand (_43020_, _42926_, _28768_);
  nor (_43021_, _43020_, _31265_);
  nor (_43022_, _38635_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_43023_, _28768_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_43024_, _19056_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_43025_, _43024_, _43023_);
  or (_43026_, _43025_, _43022_);
  or (_43027_, _43026_, _43021_);
  and (_43028_, _43027_, _42951_);
  not (_43029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_43030_, _42951_, _43029_);
  or (_02832_, _43030_, _43028_);
  not (_43031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_43032_, _42951_, _43031_);
  and (_43033_, _42951_, _42934_);
  or (_02834_, _43033_, _43032_);
  and (_43034_, _42960_, _42459_);
  and (_43035_, _42937_, _42623_);
  and (_43036_, _43035_, _42948_);
  and (_43037_, _43036_, _43034_);
  not (_43038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_43039_, _43036_, _43038_);
  or (_02842_, _43039_, _43037_);
  and (_43040_, _42975_, _42459_);
  and (_43041_, _43036_, _43040_);
  not (_43042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_43043_, _43036_, _43042_);
  or (_02845_, _43043_, _43041_);
  and (_43044_, _42986_, _42459_);
  and (_43046_, _43036_, _43044_);
  not (_43047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_43049_, _43036_, _43047_);
  or (_02848_, _43049_, _43046_);
  and (_43051_, _42994_, _42459_);
  and (_43053_, _43036_, _43051_);
  not (_43055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_43057_, _43036_, _43055_);
  or (_02853_, _43057_, _43053_);
  and (_43059_, _43005_, _42459_);
  and (_43060_, _43036_, _43059_);
  not (_43061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_43062_, _43036_, _43061_);
  or (_02856_, _43062_, _43060_);
  and (_43063_, _43016_, _42459_);
  and (_43064_, _43036_, _43063_);
  not (_43065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_43066_, _43036_, _43065_);
  or (_02859_, _43066_, _43064_);
  and (_43067_, _43027_, _42459_);
  and (_43068_, _43036_, _43067_);
  not (_43069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_43070_, _43036_, _43069_);
  or (_02862_, _43070_, _43068_);
  and (_43071_, _43036_, _42944_);
  nor (_43072_, _43036_, _42869_);
  or (_02865_, _43072_, _43071_);
  and (_43073_, _42938_, _42629_);
  and (_43074_, _43073_, _42948_);
  and (_43075_, _43074_, _43034_);
  not (_43076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_43077_, _43074_, _43076_);
  or (_02871_, _43077_, _43075_);
  and (_43078_, _43074_, _43040_);
  not (_43079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_43080_, _43074_, _43079_);
  or (_02875_, _43080_, _43078_);
  and (_43081_, _43074_, _43044_);
  not (_43082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_43083_, _43074_, _43082_);
  or (_02879_, _43083_, _43081_);
  and (_43084_, _43074_, _43051_);
  not (_43085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_43086_, _43074_, _43085_);
  or (_02882_, _43086_, _43084_);
  and (_43088_, _43074_, _43059_);
  not (_43090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_43092_, _43074_, _43090_);
  or (_02886_, _43092_, _43088_);
  and (_43095_, _43074_, _43063_);
  not (_43097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_43099_, _43074_, _43097_);
  or (_02889_, _43099_, _43095_);
  and (_43101_, _43074_, _43067_);
  not (_43103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_43105_, _43074_, _43103_);
  or (_02893_, _43105_, _43101_);
  and (_43106_, _43074_, _42944_);
  not (_43107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_43108_, _43074_, _43107_);
  or (_02895_, _43108_, _43106_);
  and (_43109_, _42948_, _42939_);
  and (_43110_, _43109_, _43034_);
  not (_43111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_43112_, _43109_, _43111_);
  or (_02901_, _43112_, _43110_);
  and (_43113_, _43109_, _43040_);
  not (_43114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_43115_, _43109_, _43114_);
  or (_02904_, _43115_, _43113_);
  and (_43116_, _43109_, _43044_);
  not (_43117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_43118_, _43109_, _43117_);
  or (_02907_, _43118_, _43116_);
  and (_43119_, _43109_, _43051_);
  not (_43120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_43121_, _43109_, _43120_);
  or (_02910_, _43121_, _43119_);
  and (_43122_, _43109_, _43059_);
  not (_43123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_43124_, _43109_, _43123_);
  or (_02914_, _43124_, _43122_);
  and (_43125_, _43109_, _43063_);
  not (_43126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_43127_, _43109_, _43126_);
  or (_02917_, _43127_, _43125_);
  and (_43128_, _43109_, _43067_);
  not (_43129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_43130_, _43109_, _43129_);
  or (_02922_, _43130_, _43128_);
  and (_43131_, _43109_, _42944_);
  nor (_43132_, _43109_, _42863_);
  or (_02925_, _43132_, _43131_);
  and (_43133_, _42941_, _42749_);
  and (_43134_, _43133_, _42949_);
  and (_43135_, _43134_, _43034_);
  not (_43136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_43137_, _43134_, _43136_);
  or (_02933_, _43137_, _43135_);
  and (_43138_, _43134_, _43040_);
  not (_43139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_43140_, _43134_, _43139_);
  or (_02937_, _43140_, _43138_);
  and (_43141_, _43134_, _43044_);
  not (_43142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_43143_, _43134_, _43142_);
  or (_02940_, _43143_, _43141_);
  and (_43144_, _43134_, _43051_);
  not (_43145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_43146_, _43134_, _43145_);
  or (_02945_, _43146_, _43144_);
  and (_43147_, _43134_, _43059_);
  not (_43148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_43149_, _43134_, _43148_);
  or (_02949_, _43149_, _43147_);
  and (_43150_, _43134_, _43063_);
  not (_43151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_43152_, _43134_, _43151_);
  or (_02952_, _43152_, _43150_);
  and (_43153_, _43134_, _43067_);
  not (_43154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_43155_, _43134_, _43154_);
  or (_02956_, _43155_, _43153_);
  and (_43156_, _43134_, _42944_);
  not (_43157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_43158_, _43134_, _43157_);
  or (_02959_, _43158_, _43156_);
  and (_43159_, _43133_, _43035_);
  and (_43160_, _43159_, _43034_);
  not (_43161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_43162_, _43159_, _43161_);
  or (_02963_, _43162_, _43160_);
  and (_43163_, _43159_, _43040_);
  not (_43164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_43165_, _43159_, _43164_);
  or (_02966_, _43165_, _43163_);
  and (_43166_, _43159_, _43044_);
  not (_43167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_43168_, _43159_, _43167_);
  or (_02971_, _43168_, _43166_);
  and (_43169_, _43159_, _43051_);
  not (_43170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_43171_, _43159_, _43170_);
  or (_02974_, _43171_, _43169_);
  and (_43172_, _43159_, _43059_);
  not (_43173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_43174_, _43159_, _43173_);
  or (_02977_, _43174_, _43172_);
  and (_43175_, _43159_, _43063_);
  not (_43176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_43177_, _43159_, _43176_);
  or (_02981_, _43177_, _43175_);
  and (_43178_, _43159_, _43067_);
  not (_43179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_43180_, _43159_, _43179_);
  or (_02985_, _43180_, _43178_);
  and (_43181_, _43159_, _42944_);
  nor (_43182_, _43159_, _42882_);
  or (_02987_, _43182_, _43181_);
  and (_43183_, _43133_, _43073_);
  and (_43184_, _43183_, _43034_);
  not (_43185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_43186_, _43183_, _43185_);
  or (_02992_, _43186_, _43184_);
  and (_43187_, _43183_, _43040_);
  not (_43188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_43189_, _43183_, _43188_);
  or (_02996_, _43189_, _43187_);
  and (_43190_, _43183_, _43044_);
  not (_43191_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_43192_, _43183_, _43191_);
  or (_03000_, _43192_, _43190_);
  and (_43193_, _43183_, _43051_);
  not (_43194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_43195_, _43183_, _43194_);
  or (_03003_, _43195_, _43193_);
  and (_43196_, _43183_, _43059_);
  not (_43197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_43198_, _43183_, _43197_);
  or (_03008_, _43198_, _43196_);
  and (_43199_, _43183_, _43063_);
  not (_43200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_43201_, _43183_, _43200_);
  or (_03012_, _43201_, _43199_);
  and (_43202_, _43183_, _43067_);
  not (_43203_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_43204_, _43183_, _43203_);
  or (_03015_, _43204_, _43202_);
  and (_43205_, _43183_, _42944_);
  not (_43206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_43207_, _43183_, _43206_);
  or (_03018_, _43207_, _43205_);
  and (_43208_, _43133_, _42939_);
  and (_43209_, _43208_, _43034_);
  not (_43210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_43211_, _43208_, _43210_);
  or (_03023_, _43211_, _43209_);
  and (_43212_, _43208_, _43040_);
  not (_43213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_43214_, _43208_, _43213_);
  or (_03027_, _43214_, _43212_);
  and (_43215_, _43208_, _43044_);
  not (_43216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_43217_, _43208_, _43216_);
  or (_03030_, _43217_, _43215_);
  and (_43218_, _43208_, _43051_);
  not (_43219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_43220_, _43208_, _43219_);
  or (_03034_, _43220_, _43218_);
  and (_43221_, _43208_, _43059_);
  not (_43222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_43223_, _43208_, _43222_);
  or (_03038_, _43223_, _43221_);
  and (_43224_, _43208_, _43063_);
  not (_43225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_43226_, _43208_, _43225_);
  or (_03041_, _43226_, _43224_);
  and (_43227_, _43208_, _43067_);
  not (_43228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_43229_, _43208_, _43228_);
  or (_03045_, _43229_, _43227_);
  and (_43230_, _43208_, _42944_);
  nor (_43231_, _43208_, _42876_);
  or (_03047_, _43231_, _43230_);
  and (_43232_, _42940_, _42828_);
  and (_43233_, _43232_, _42949_);
  and (_43234_, _43233_, _43034_);
  not (_43235_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_43236_, _43233_, _43235_);
  or (_03054_, _43236_, _43234_);
  and (_43237_, _43233_, _43040_);
  not (_43238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_43239_, _43233_, _43238_);
  or (_03058_, _43239_, _43237_);
  and (_43240_, _43233_, _43044_);
  not (_43241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_43242_, _43233_, _43241_);
  or (_03062_, _43242_, _43240_);
  and (_43243_, _43233_, _43051_);
  not (_43244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_43245_, _43233_, _43244_);
  or (_03065_, _43245_, _43243_);
  and (_43246_, _43233_, _43059_);
  not (_43247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_43248_, _43233_, _43247_);
  or (_03069_, _43248_, _43246_);
  and (_43249_, _43233_, _43063_);
  not (_43250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_43251_, _43233_, _43250_);
  or (_03072_, _43251_, _43249_);
  and (_43252_, _43233_, _43067_);
  not (_43253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_43254_, _43233_, _43253_);
  or (_03076_, _43254_, _43252_);
  and (_43255_, _43233_, _42944_);
  nor (_43256_, _43233_, _42891_);
  or (_03078_, _43256_, _43255_);
  and (_43257_, _43232_, _43035_);
  and (_43258_, _43257_, _43034_);
  not (_43259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_43260_, _43257_, _43259_);
  or (_03083_, _43260_, _43258_);
  and (_43261_, _43257_, _43040_);
  not (_43262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_43263_, _43257_, _43262_);
  or (_03086_, _43263_, _43261_);
  and (_43264_, _43257_, _43044_);
  not (_43265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_43266_, _43257_, _43265_);
  or (_03090_, _43266_, _43264_);
  and (_43267_, _43257_, _43051_);
  not (_43268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_43269_, _43257_, _43268_);
  or (_03094_, _43269_, _43267_);
  and (_43270_, _43257_, _43059_);
  not (_43271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_43272_, _43257_, _43271_);
  or (_03097_, _43272_, _43270_);
  and (_43273_, _43257_, _43063_);
  not (_43274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_43275_, _43257_, _43274_);
  or (_03101_, _43275_, _43273_);
  and (_43276_, _43257_, _43067_);
  not (_43277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_43278_, _43257_, _43277_);
  or (_03104_, _43278_, _43276_);
  and (_43279_, _43257_, _42944_);
  not (_43280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_43281_, _43257_, _43280_);
  or (_03107_, _43281_, _43279_);
  and (_43282_, _43232_, _43073_);
  and (_43283_, _43282_, _43034_);
  not (_43284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_43285_, _43282_, _43284_);
  or (_03111_, _43285_, _43283_);
  and (_43286_, _43282_, _43040_);
  not (_43287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_43288_, _43282_, _43287_);
  or (_03115_, _43288_, _43286_);
  and (_43289_, _43282_, _43044_);
  not (_43290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_43291_, _43282_, _43290_);
  or (_03119_, _43291_, _43289_);
  and (_43292_, _43282_, _43051_);
  not (_43293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_43294_, _43282_, _43293_);
  or (_03122_, _43294_, _43292_);
  and (_43295_, _43282_, _43059_);
  not (_43296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_43297_, _43282_, _43296_);
  or (_03127_, _43297_, _43295_);
  and (_43298_, _43282_, _43063_);
  not (_43299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_43300_, _43282_, _43299_);
  or (_03130_, _43300_, _43298_);
  and (_43301_, _43282_, _43067_);
  not (_43302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_43303_, _43282_, _43302_);
  or (_03134_, _43303_, _43301_);
  and (_43304_, _43282_, _42944_);
  nor (_43305_, _43282_, _42897_);
  or (_03137_, _43305_, _43304_);
  and (_43306_, _43232_, _42939_);
  and (_43307_, _43306_, _43034_);
  not (_43308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_43309_, _43306_, _43308_);
  or (_03141_, _43309_, _43307_);
  and (_43310_, _43306_, _43040_);
  not (_43311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_43312_, _43306_, _43311_);
  or (_03145_, _43312_, _43310_);
  and (_43313_, _43306_, _43044_);
  not (_43314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_43315_, _43306_, _43314_);
  or (_03148_, _43315_, _43313_);
  and (_43316_, _43306_, _43051_);
  not (_43317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_43318_, _43306_, _43317_);
  or (_03152_, _43318_, _43316_);
  and (_43319_, _43306_, _43059_);
  not (_43320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_43321_, _43306_, _43320_);
  or (_03155_, _43321_, _43319_);
  and (_43322_, _43306_, _43063_);
  not (_43323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_43324_, _43306_, _43323_);
  or (_03159_, _43324_, _43322_);
  and (_43325_, _43306_, _43067_);
  not (_43326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_43327_, _43306_, _43326_);
  or (_03162_, _43327_, _43325_);
  and (_43328_, _43306_, _42944_);
  not (_43329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_43330_, _43306_, _43329_);
  or (_03165_, _43330_, _43328_);
  and (_43331_, _42949_, _42942_);
  and (_43332_, _43331_, _43034_);
  not (_43333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_43334_, _43331_, _43333_);
  or (_03170_, _43334_, _43332_);
  and (_43335_, _43331_, _43040_);
  not (_43336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_43337_, _43331_, _43336_);
  or (_03173_, _43337_, _43335_);
  and (_43338_, _43331_, _43044_);
  not (_43339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_43340_, _43331_, _43339_);
  or (_03177_, _43340_, _43338_);
  and (_43341_, _43331_, _43051_);
  not (_43342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_43343_, _43331_, _43342_);
  or (_03181_, _43343_, _43341_);
  and (_43344_, _43331_, _43059_);
  not (_43345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_43346_, _43331_, _43345_);
  or (_03185_, _43346_, _43344_);
  and (_43347_, _43331_, _43063_);
  not (_43348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_43349_, _43331_, _43348_);
  or (_03189_, _43349_, _43347_);
  and (_43350_, _43331_, _43067_);
  not (_43351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_43352_, _43331_, _43351_);
  or (_03193_, _43352_, _43350_);
  and (_43353_, _43331_, _42944_);
  nor (_43354_, _43331_, _42903_);
  or (_03196_, _43354_, _43353_);
  and (_43355_, _43035_, _42942_);
  and (_43356_, _43355_, _43034_);
  not (_43357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_43358_, _43355_, _43357_);
  or (_03201_, _43358_, _43356_);
  and (_43359_, _43355_, _43040_);
  not (_43360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_43361_, _43355_, _43360_);
  or (_03205_, _43361_, _43359_);
  and (_43362_, _43355_, _43044_);
  not (_43363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_43364_, _43355_, _43363_);
  or (_03209_, _43364_, _43362_);
  and (_43365_, _43355_, _43051_);
  not (_43366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_43367_, _43355_, _43366_);
  or (_03213_, _43367_, _43365_);
  and (_43368_, _43355_, _43059_);
  not (_43369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_43370_, _43355_, _43369_);
  or (_03217_, _43370_, _43368_);
  and (_43371_, _43355_, _43063_);
  not (_43372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_43373_, _43355_, _43372_);
  or (_03221_, _43373_, _43371_);
  and (_43374_, _43355_, _43067_);
  not (_43375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_43376_, _43355_, _43375_);
  or (_03225_, _43376_, _43374_);
  and (_43377_, _43355_, _42944_);
  not (_43378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_43379_, _43355_, _43378_);
  or (_03228_, _43379_, _43377_);
  and (_43380_, _43073_, _42942_);
  and (_43381_, _43380_, _43034_);
  not (_43382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_43383_, _43380_, _43382_);
  or (_03233_, _43383_, _43381_);
  and (_43384_, _43380_, _43040_);
  not (_43385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_43386_, _43380_, _43385_);
  or (_03237_, _43386_, _43384_);
  and (_43387_, _43380_, _43044_);
  not (_43388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_43389_, _43380_, _43388_);
  or (_03241_, _43389_, _43387_);
  and (_43390_, _43380_, _43051_);
  not (_43391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_43392_, _43380_, _43391_);
  or (_03245_, _43392_, _43390_);
  and (_43393_, _43380_, _43059_);
  not (_43394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_43395_, _43380_, _43394_);
  or (_03249_, _43395_, _43393_);
  and (_43396_, _43380_, _43063_);
  not (_43397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_43398_, _43380_, _43397_);
  or (_03253_, _43398_, _43396_);
  and (_43399_, _43380_, _43067_);
  not (_43400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_43401_, _43380_, _43400_);
  or (_03257_, _43401_, _43399_);
  and (_43402_, _43380_, _42944_);
  nor (_43403_, _43380_, _42909_);
  or (_03260_, _43403_, _43402_);
  and (_43404_, _43034_, _42943_);
  not (_43405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_43406_, _42943_, _43405_);
  or (_03265_, _43406_, _43404_);
  and (_43407_, _43040_, _42943_);
  not (_43408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_43409_, _42943_, _43408_);
  or (_03269_, _43409_, _43407_);
  and (_43410_, _43044_, _42943_);
  not (_43411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_43412_, _42943_, _43411_);
  or (_03273_, _43412_, _43410_);
  and (_43413_, _43051_, _42943_);
  not (_43414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_43415_, _42943_, _43414_);
  or (_03277_, _43415_, _43413_);
  and (_43416_, _43059_, _42943_);
  not (_43417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_43418_, _42943_, _43417_);
  or (_03281_, _43418_, _43416_);
  and (_43419_, _43063_, _42943_);
  not (_43420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_43421_, _42943_, _43420_);
  or (_03285_, _43421_, _43419_);
  and (_43422_, _43067_, _42943_);
  not (_43423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_43424_, _42943_, _43423_);
  or (_03289_, _43424_, _43422_);
  nor (_43425_, _42703_, _43111_);
  and (_43426_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_43427_, _43426_, _42619_);
  or (_43428_, _43427_, _43425_);
  and (_43429_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_43430_, _42703_, _43038_);
  nand (_43431_, _43430_, _42619_);
  or (_43432_, _43431_, _43429_);
  and (_43433_, _43432_, _43428_);
  or (_43434_, _43433_, _42862_);
  nor (_43435_, _42703_, _43210_);
  and (_43436_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_43437_, _43436_, _42619_);
  or (_43438_, _43437_, _43435_);
  and (_43439_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_43440_, _42703_, _43161_);
  nand (_43441_, _43440_, _42619_);
  or (_43442_, _43441_, _43439_);
  and (_43443_, _43442_, _43438_);
  or (_43444_, _43443_, _42825_);
  and (_43445_, _43444_, _42875_);
  and (_43446_, _43445_, _43434_);
  nand (_43447_, _42703_, _43235_);
  or (_43448_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_43449_, _43448_, _43447_);
  or (_43450_, _43449_, _42890_);
  or (_43451_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand (_43452_, _42703_, _43284_);
  and (_43453_, _43452_, _43451_);
  or (_43454_, _43453_, _42619_);
  and (_43455_, _43454_, _43450_);
  or (_43456_, _43455_, _42862_);
  nand (_43457_, _42703_, _43333_);
  or (_43458_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_43459_, _43458_, _43457_);
  or (_43460_, _43459_, _42890_);
  or (_43461_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand (_43462_, _42703_, _43382_);
  and (_43463_, _43462_, _43461_);
  or (_43464_, _43463_, _42619_);
  and (_43465_, _43464_, _43460_);
  or (_43466_, _43465_, _42825_);
  and (_43467_, _43466_, _42745_);
  and (_43468_, _43467_, _43456_);
  or (_43469_, _43468_, _43446_);
  or (_43470_, _43469_, _42861_);
  or (_43471_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_43472_, _43471_, _42923_);
  and (_43473_, _43472_, _43470_);
  and (_40258_, _42960_, _43100_);
  and (_43474_, _40258_, _42922_);
  or (_05085_, _43474_, _43473_);
  nor (_43475_, _42703_, _43114_);
  and (_43476_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_43477_, _43476_, _42619_);
  or (_43478_, _43477_, _43475_);
  and (_43479_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_43480_, _42703_, _43042_);
  nand (_43481_, _43480_, _42619_);
  or (_43482_, _43481_, _43479_);
  and (_43483_, _43482_, _43478_);
  or (_43484_, _43483_, _42862_);
  nor (_43485_, _42703_, _43213_);
  and (_43486_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_43487_, _43486_, _42619_);
  or (_43488_, _43487_, _43485_);
  and (_43489_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_43490_, _42703_, _43164_);
  nand (_43491_, _43490_, _42619_);
  or (_43492_, _43491_, _43489_);
  and (_43493_, _43492_, _43488_);
  or (_43494_, _43493_, _42825_);
  and (_43495_, _43494_, _42875_);
  and (_43496_, _43495_, _43484_);
  nand (_43497_, _42703_, _43238_);
  or (_43498_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_43499_, _43498_, _43497_);
  or (_43500_, _43499_, _42890_);
  or (_43501_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand (_43502_, _42703_, _43287_);
  and (_43503_, _43502_, _43501_);
  or (_43504_, _43503_, _42619_);
  and (_43505_, _43504_, _43500_);
  or (_43506_, _43505_, _42862_);
  nand (_43507_, _42703_, _43336_);
  or (_43508_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_43509_, _43508_, _43507_);
  or (_43510_, _43509_, _42890_);
  or (_43511_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand (_43512_, _42703_, _43385_);
  and (_43513_, _43512_, _43511_);
  or (_43514_, _43513_, _42619_);
  and (_43515_, _43514_, _43510_);
  or (_43516_, _43515_, _42825_);
  and (_43517_, _43516_, _42745_);
  and (_43518_, _43517_, _43506_);
  or (_43519_, _43518_, _43496_);
  or (_43520_, _43519_, _42861_);
  or (_43521_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_43522_, _43521_, _42923_);
  and (_43523_, _43522_, _43520_);
  and (_40259_, _42975_, _43100_);
  and (_43524_, _40259_, _42922_);
  or (_05087_, _43524_, _43523_);
  nor (_43525_, _42703_, _43117_);
  and (_43526_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_43527_, _43526_, _42619_);
  or (_43528_, _43527_, _43525_);
  and (_43529_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_43530_, _42703_, _43047_);
  nand (_43531_, _43530_, _42619_);
  or (_43532_, _43531_, _43529_);
  and (_43533_, _43532_, _43528_);
  or (_43534_, _43533_, _42862_);
  nor (_43535_, _42703_, _43216_);
  and (_43536_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_43537_, _43536_, _42619_);
  or (_43538_, _43537_, _43535_);
  and (_43539_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_43540_, _42703_, _43167_);
  nand (_43541_, _43540_, _42619_);
  or (_43542_, _43541_, _43539_);
  and (_43543_, _43542_, _43538_);
  or (_43544_, _43543_, _42825_);
  and (_43545_, _43544_, _42875_);
  and (_43546_, _43545_, _43534_);
  nand (_43547_, _42703_, _43241_);
  or (_43548_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_43549_, _43548_, _43547_);
  or (_43550_, _43549_, _42890_);
  or (_43551_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_43552_, _42703_, _43290_);
  and (_43553_, _43552_, _43551_);
  or (_43554_, _43553_, _42619_);
  and (_43555_, _43554_, _43550_);
  or (_43556_, _43555_, _42862_);
  nand (_43557_, _42703_, _43339_);
  or (_43558_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_43559_, _43558_, _43557_);
  or (_43560_, _43559_, _42890_);
  or (_43561_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_43562_, _42703_, _43388_);
  and (_43563_, _43562_, _43561_);
  or (_43564_, _43563_, _42619_);
  and (_43565_, _43564_, _43560_);
  or (_43566_, _43565_, _42825_);
  and (_43567_, _43566_, _42745_);
  and (_43568_, _43567_, _43556_);
  or (_43569_, _43568_, _43546_);
  or (_43570_, _43569_, _42861_);
  or (_43571_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_43572_, _43571_, _42923_);
  and (_43573_, _43572_, _43570_);
  and (_40260_, _42986_, _43100_);
  and (_43574_, _40260_, _42922_);
  or (_05089_, _43574_, _43573_);
  nor (_43575_, _42703_, _43120_);
  and (_43576_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_43577_, _43576_, _42619_);
  or (_43578_, _43577_, _43575_);
  and (_43579_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_43580_, _42703_, _43055_);
  nand (_43581_, _43580_, _42619_);
  or (_43582_, _43581_, _43579_);
  and (_43583_, _43582_, _43578_);
  or (_43584_, _43583_, _42862_);
  nor (_43585_, _42703_, _43219_);
  and (_43586_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_43587_, _43586_, _42619_);
  or (_43588_, _43587_, _43585_);
  and (_43589_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_43590_, _42703_, _43170_);
  nand (_43591_, _43590_, _42619_);
  or (_43592_, _43591_, _43589_);
  and (_43593_, _43592_, _43588_);
  or (_43597_, _43593_, _42825_);
  and (_43602_, _43597_, _42875_);
  and (_43610_, _43602_, _43584_);
  nand (_43616_, _42703_, _43244_);
  or (_43620_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_43627_, _43620_, _43616_);
  or (_43635_, _43627_, _42890_);
  or (_43639_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_43644_, _42703_, _43293_);
  and (_43652_, _43644_, _43639_);
  or (_43658_, _43652_, _42619_);
  and (_43662_, _43658_, _43635_);
  or (_43669_, _43662_, _42862_);
  nand (_43677_, _42703_, _43342_);
  or (_43681_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_43686_, _43681_, _43677_);
  or (_43688_, _43686_, _42890_);
  or (_43699_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_43704_, _42703_, _43391_);
  and (_43712_, _43704_, _43699_);
  or (_43718_, _43712_, _42619_);
  and (_43722_, _43718_, _43688_);
  or (_43729_, _43722_, _42825_);
  and (_43737_, _43729_, _42745_);
  and (_43741_, _43737_, _43669_);
  or (_43746_, _43741_, _43610_);
  or (_43754_, _43746_, _42861_);
  or (_43760_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_43764_, _43760_, _42923_);
  and (_43771_, _43764_, _43754_);
  and (_40261_, _42994_, _43100_);
  and (_43782_, _40261_, _42922_);
  or (_05091_, _43782_, _43771_);
  and (_43787_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_43788_, _42703_, _43061_);
  nand (_43789_, _43788_, _42619_);
  or (_43790_, _43789_, _43787_);
  nor (_43791_, _42703_, _43123_);
  and (_43792_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_43793_, _43792_, _42619_);
  or (_43794_, _43793_, _43791_);
  and (_43795_, _43794_, _43790_);
  or (_43796_, _43795_, _42862_);
  nor (_43797_, _42703_, _43222_);
  and (_43798_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_43799_, _43798_, _42619_);
  or (_43800_, _43799_, _43797_);
  and (_43801_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_43802_, _42703_, _43173_);
  nand (_43803_, _43802_, _42619_);
  or (_43804_, _43803_, _43801_);
  and (_43805_, _43804_, _43800_);
  or (_43806_, _43805_, _42825_);
  and (_43807_, _43806_, _42875_);
  and (_43808_, _43807_, _43796_);
  nor (_43809_, _42703_, _43320_);
  and (_43810_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_43811_, _43810_, _42619_);
  or (_43812_, _43811_, _43809_);
  and (_43813_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_43814_, _42703_, _43271_);
  nand (_43815_, _43814_, _42619_);
  or (_43816_, _43815_, _43813_);
  and (_43817_, _43816_, _43812_);
  or (_43818_, _43817_, _42862_);
  nor (_43819_, _42703_, _43417_);
  and (_43820_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_43821_, _43820_, _42619_);
  or (_43822_, _43821_, _43819_);
  and (_43823_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_43824_, _42703_, _43369_);
  nand (_43825_, _43824_, _42619_);
  or (_43826_, _43825_, _43823_);
  and (_43827_, _43826_, _43822_);
  or (_43828_, _43827_, _42825_);
  and (_43829_, _43828_, _42745_);
  and (_43830_, _43829_, _43818_);
  or (_43831_, _43830_, _43808_);
  and (_43832_, _43831_, _42921_);
  and (_43833_, _43005_, _42922_);
  and (_43834_, _42861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or (_43835_, _43834_, _43833_);
  or (_43836_, _43835_, _43832_);
  and (_05093_, _43836_, _43100_);
  or (_43837_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_43838_, _42703_, _43397_);
  and (_43839_, _43838_, _43837_);
  or (_43840_, _43839_, _42619_);
  nand (_43841_, _42703_, _43348_);
  or (_43842_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_43843_, _43842_, _43841_);
  or (_43844_, _43843_, _42890_);
  and (_43845_, _43844_, _42745_);
  and (_43846_, _43845_, _43840_);
  and (_43847_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_43848_, _42703_, _43176_);
  nand (_43849_, _43848_, _42619_);
  or (_43850_, _43849_, _43847_);
  nor (_43851_, _42703_, _43225_);
  and (_43852_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_43853_, _43852_, _42619_);
  or (_43854_, _43853_, _43851_);
  and (_43855_, _43854_, _42875_);
  and (_43856_, _43855_, _43850_);
  or (_43857_, _43856_, _43846_);
  and (_43858_, _43857_, _42862_);
  or (_43859_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_43860_, _42703_, _43299_);
  and (_43861_, _43860_, _43859_);
  or (_43862_, _43861_, _42619_);
  nand (_43863_, _42703_, _43250_);
  or (_43864_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_43865_, _43864_, _43863_);
  or (_43866_, _43865_, _42890_);
  and (_43867_, _43866_, _42745_);
  and (_43868_, _43867_, _43862_);
  and (_43869_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_43870_, _42703_, _43065_);
  nand (_43871_, _43870_, _42619_);
  or (_43872_, _43871_, _43869_);
  nor (_43873_, _42703_, _43126_);
  and (_43874_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_43875_, _43874_, _42619_);
  or (_43876_, _43875_, _43873_);
  and (_43877_, _43876_, _42875_);
  and (_43878_, _43877_, _43872_);
  or (_43879_, _43878_, _43868_);
  and (_43880_, _43879_, _42825_);
  or (_43881_, _43880_, _42835_);
  or (_43882_, _43881_, _43858_);
  or (_43883_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_40263_, _43016_, _43100_);
  or (_43884_, _40263_, _42923_);
  and (_43885_, _43884_, _43883_);
  and (_05095_, _43885_, _43882_);
  nor (_43886_, _42703_, _43129_);
  and (_43887_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_43888_, _43887_, _42619_);
  or (_43889_, _43888_, _43886_);
  and (_43890_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_43891_, _42703_, _43069_);
  nand (_43892_, _43891_, _42619_);
  or (_43893_, _43892_, _43890_);
  and (_43894_, _43893_, _43889_);
  or (_43895_, _43894_, _42862_);
  nor (_43896_, _42703_, _43228_);
  and (_43897_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_43898_, _43897_, _42619_);
  or (_43899_, _43898_, _43896_);
  and (_43900_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_43901_, _42703_, _43179_);
  nand (_43902_, _43901_, _42619_);
  or (_43903_, _43902_, _43900_);
  and (_43904_, _43903_, _43899_);
  or (_43905_, _43904_, _42825_);
  and (_43906_, _43905_, _42875_);
  and (_43907_, _43906_, _43895_);
  nand (_43908_, _42703_, _43253_);
  or (_43909_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_43910_, _43909_, _43908_);
  or (_43911_, _43910_, _42890_);
  or (_43912_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_43913_, _42703_, _43302_);
  and (_43914_, _43913_, _43912_);
  or (_43915_, _43914_, _42619_);
  and (_43916_, _43915_, _43911_);
  or (_43917_, _43916_, _42862_);
  nand (_43918_, _42703_, _43351_);
  or (_43919_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_43920_, _43919_, _43918_);
  or (_43921_, _43920_, _42890_);
  or (_43922_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_43923_, _42703_, _43400_);
  and (_43924_, _43923_, _43922_);
  or (_43925_, _43924_, _42619_);
  and (_43926_, _43925_, _43921_);
  or (_43927_, _43926_, _42825_);
  and (_43928_, _43927_, _42745_);
  and (_43929_, _43928_, _43917_);
  or (_43930_, _43929_, _43907_);
  or (_43931_, _43930_, _42861_);
  or (_43932_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_43933_, _43932_, _42923_);
  and (_43934_, _43933_, _43931_);
  and (_40264_, _43027_, _43100_);
  and (_43935_, _40264_, _42922_);
  or (_05097_, _43935_, _43934_);
  or (_43936_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_43937_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_43938_, _43937_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_43939_, _43938_, _43936_);
  nand (_43940_, _43939_, _43100_);
  or (_43941_, \oc8051_gm_cxrom_1.cell0.data [7], _43100_);
  and (_05105_, _43941_, _43940_);
  or (_43942_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43943_, \oc8051_gm_cxrom_1.cell0.data [0], _43937_);
  nand (_43944_, _43943_, _43942_);
  nand (_43945_, _43944_, _43100_);
  or (_43946_, \oc8051_gm_cxrom_1.cell0.data [0], _43100_);
  and (_05111_, _43946_, _43945_);
  or (_43947_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43948_, \oc8051_gm_cxrom_1.cell0.data [1], _43937_);
  nand (_43949_, _43948_, _43947_);
  nand (_43950_, _43949_, _43100_);
  or (_43951_, \oc8051_gm_cxrom_1.cell0.data [1], _43100_);
  and (_05115_, _43951_, _43950_);
  or (_43952_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43953_, \oc8051_gm_cxrom_1.cell0.data [2], _43937_);
  nand (_43954_, _43953_, _43952_);
  nand (_43955_, _43954_, _43100_);
  or (_43956_, \oc8051_gm_cxrom_1.cell0.data [2], _43100_);
  and (_05119_, _43956_, _43955_);
  or (_43957_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43958_, \oc8051_gm_cxrom_1.cell0.data [3], _43937_);
  nand (_43959_, _43958_, _43957_);
  nand (_43960_, _43959_, _43100_);
  or (_43961_, \oc8051_gm_cxrom_1.cell0.data [3], _43100_);
  and (_05123_, _43961_, _43960_);
  or (_43962_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43963_, \oc8051_gm_cxrom_1.cell0.data [4], _43937_);
  nand (_43964_, _43963_, _43962_);
  nand (_43965_, _43964_, _43100_);
  or (_43966_, \oc8051_gm_cxrom_1.cell0.data [4], _43100_);
  and (_05127_, _43966_, _43965_);
  or (_43967_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43968_, \oc8051_gm_cxrom_1.cell0.data [5], _43937_);
  nand (_43969_, _43968_, _43967_);
  nand (_43970_, _43969_, _43100_);
  or (_43971_, \oc8051_gm_cxrom_1.cell0.data [5], _43100_);
  and (_05131_, _43971_, _43970_);
  or (_43972_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43973_, \oc8051_gm_cxrom_1.cell0.data [6], _43937_);
  nand (_43974_, _43973_, _43972_);
  nand (_43975_, _43974_, _43100_);
  or (_43976_, \oc8051_gm_cxrom_1.cell0.data [6], _43100_);
  and (_05135_, _43976_, _43975_);
  or (_43977_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_43978_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_43979_, _43978_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_43980_, _43979_, _43977_);
  nand (_43981_, _43980_, _43100_);
  or (_43982_, \oc8051_gm_cxrom_1.cell1.data [7], _43100_);
  and (_05156_, _43982_, _43981_);
  or (_43983_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43984_, \oc8051_gm_cxrom_1.cell1.data [0], _43978_);
  nand (_43985_, _43984_, _43983_);
  nand (_43986_, _43985_, _43100_);
  or (_43987_, \oc8051_gm_cxrom_1.cell1.data [0], _43100_);
  and (_05163_, _43987_, _43986_);
  or (_43988_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43989_, \oc8051_gm_cxrom_1.cell1.data [1], _43978_);
  nand (_43990_, _43989_, _43988_);
  nand (_43991_, _43990_, _43100_);
  or (_43992_, \oc8051_gm_cxrom_1.cell1.data [1], _43100_);
  and (_05167_, _43992_, _43991_);
  or (_43993_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43994_, \oc8051_gm_cxrom_1.cell1.data [2], _43978_);
  nand (_43995_, _43994_, _43993_);
  nand (_43996_, _43995_, _43100_);
  or (_43997_, \oc8051_gm_cxrom_1.cell1.data [2], _43100_);
  and (_05171_, _43997_, _43996_);
  or (_43998_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43999_, \oc8051_gm_cxrom_1.cell1.data [3], _43978_);
  nand (_44000_, _43999_, _43998_);
  nand (_44001_, _44000_, _43100_);
  or (_44002_, \oc8051_gm_cxrom_1.cell1.data [3], _43100_);
  and (_05175_, _44002_, _44001_);
  or (_44003_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_44004_, \oc8051_gm_cxrom_1.cell1.data [4], _43978_);
  nand (_44005_, _44004_, _44003_);
  nand (_44006_, _44005_, _43100_);
  or (_44007_, \oc8051_gm_cxrom_1.cell1.data [4], _43100_);
  and (_05179_, _44007_, _44006_);
  or (_44008_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_44009_, \oc8051_gm_cxrom_1.cell1.data [5], _43978_);
  nand (_44010_, _44009_, _44008_);
  nand (_44011_, _44010_, _43100_);
  or (_44012_, \oc8051_gm_cxrom_1.cell1.data [5], _43100_);
  and (_05183_, _44012_, _44011_);
  or (_44013_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_44014_, \oc8051_gm_cxrom_1.cell1.data [6], _43978_);
  nand (_44015_, _44014_, _44013_);
  nand (_44016_, _44015_, _43100_);
  or (_44017_, \oc8051_gm_cxrom_1.cell1.data [6], _43100_);
  and (_05186_, _44017_, _44016_);
  or (_44018_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_44019_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_44020_, _44019_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_44021_, _44020_, _44018_);
  nand (_44022_, _44021_, _43100_);
  or (_44023_, \oc8051_gm_cxrom_1.cell2.data [7], _43100_);
  and (_05208_, _44023_, _44022_);
  or (_44024_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_44025_, \oc8051_gm_cxrom_1.cell2.data [0], _44019_);
  nand (_44026_, _44025_, _44024_);
  nand (_44027_, _44026_, _43100_);
  or (_44028_, \oc8051_gm_cxrom_1.cell2.data [0], _43100_);
  and (_05215_, _44028_, _44027_);
  or (_00002_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00003_, \oc8051_gm_cxrom_1.cell2.data [1], _44019_);
  nand (_00004_, _00003_, _00002_);
  nand (_00005_, _00004_, _43100_);
  or (_00006_, \oc8051_gm_cxrom_1.cell2.data [1], _43100_);
  and (_05219_, _00006_, _00005_);
  or (_00007_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00008_, \oc8051_gm_cxrom_1.cell2.data [2], _44019_);
  nand (_00009_, _00008_, _00007_);
  nand (_00010_, _00009_, _43100_);
  or (_00011_, \oc8051_gm_cxrom_1.cell2.data [2], _43100_);
  and (_05222_, _00011_, _00010_);
  or (_00012_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00013_, \oc8051_gm_cxrom_1.cell2.data [3], _44019_);
  nand (_00014_, _00013_, _00012_);
  nand (_00015_, _00014_, _43100_);
  or (_00016_, \oc8051_gm_cxrom_1.cell2.data [3], _43100_);
  and (_05226_, _00016_, _00015_);
  or (_00017_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00018_, \oc8051_gm_cxrom_1.cell2.data [4], _44019_);
  nand (_00019_, _00018_, _00017_);
  nand (_00020_, _00019_, _43100_);
  or (_00021_, \oc8051_gm_cxrom_1.cell2.data [4], _43100_);
  and (_05230_, _00021_, _00020_);
  or (_00022_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00023_, \oc8051_gm_cxrom_1.cell2.data [5], _44019_);
  nand (_00024_, _00023_, _00022_);
  nand (_00025_, _00024_, _43100_);
  or (_00026_, \oc8051_gm_cxrom_1.cell2.data [5], _43100_);
  and (_05234_, _00026_, _00025_);
  or (_00027_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00028_, \oc8051_gm_cxrom_1.cell2.data [6], _44019_);
  nand (_00029_, _00028_, _00027_);
  nand (_00030_, _00029_, _43100_);
  or (_00031_, \oc8051_gm_cxrom_1.cell2.data [6], _43100_);
  and (_05238_, _00031_, _00030_);
  or (_00032_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_00033_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_00034_, _00033_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_00035_, _00034_, _00032_);
  nand (_00036_, _00035_, _43100_);
  or (_00037_, \oc8051_gm_cxrom_1.cell3.data [7], _43100_);
  and (_05259_, _00037_, _00036_);
  or (_00038_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00039_, \oc8051_gm_cxrom_1.cell3.data [0], _00033_);
  nand (_00040_, _00039_, _00038_);
  nand (_00041_, _00040_, _43100_);
  or (_00042_, \oc8051_gm_cxrom_1.cell3.data [0], _43100_);
  and (_05266_, _00042_, _00041_);
  or (_00043_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00044_, \oc8051_gm_cxrom_1.cell3.data [1], _00033_);
  nand (_00045_, _00044_, _00043_);
  nand (_00046_, _00045_, _43100_);
  or (_00047_, \oc8051_gm_cxrom_1.cell3.data [1], _43100_);
  and (_05270_, _00047_, _00046_);
  or (_00048_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00049_, \oc8051_gm_cxrom_1.cell3.data [2], _00033_);
  nand (_00050_, _00049_, _00048_);
  nand (_00051_, _00050_, _43100_);
  or (_00052_, \oc8051_gm_cxrom_1.cell3.data [2], _43100_);
  and (_05274_, _00052_, _00051_);
  or (_00053_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00054_, \oc8051_gm_cxrom_1.cell3.data [3], _00033_);
  nand (_00055_, _00054_, _00053_);
  nand (_00056_, _00055_, _43100_);
  or (_00057_, \oc8051_gm_cxrom_1.cell3.data [3], _43100_);
  and (_05278_, _00057_, _00056_);
  or (_00058_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00059_, \oc8051_gm_cxrom_1.cell3.data [4], _00033_);
  nand (_00060_, _00059_, _00058_);
  nand (_00061_, _00060_, _43100_);
  or (_00062_, \oc8051_gm_cxrom_1.cell3.data [4], _43100_);
  and (_05282_, _00062_, _00061_);
  or (_00063_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00064_, \oc8051_gm_cxrom_1.cell3.data [5], _00033_);
  nand (_00065_, _00064_, _00063_);
  nand (_00066_, _00065_, _43100_);
  or (_00067_, \oc8051_gm_cxrom_1.cell3.data [5], _43100_);
  and (_05286_, _00067_, _00066_);
  or (_00068_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00069_, \oc8051_gm_cxrom_1.cell3.data [6], _00033_);
  nand (_00070_, _00069_, _00068_);
  nand (_00071_, _00070_, _43100_);
  or (_00072_, \oc8051_gm_cxrom_1.cell3.data [6], _43100_);
  and (_05290_, _00072_, _00071_);
  or (_00073_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_00074_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_00075_, _00074_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_00076_, _00075_, _00073_);
  nand (_00077_, _00076_, _43100_);
  or (_00078_, \oc8051_gm_cxrom_1.cell4.data [7], _43100_);
  and (_05311_, _00078_, _00077_);
  or (_00079_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00080_, \oc8051_gm_cxrom_1.cell4.data [0], _00074_);
  nand (_00081_, _00080_, _00079_);
  nand (_00082_, _00081_, _43100_);
  or (_00083_, \oc8051_gm_cxrom_1.cell4.data [0], _43100_);
  and (_05318_, _00083_, _00082_);
  or (_00084_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00085_, \oc8051_gm_cxrom_1.cell4.data [1], _00074_);
  nand (_00086_, _00085_, _00084_);
  nand (_00087_, _00086_, _43100_);
  or (_00088_, \oc8051_gm_cxrom_1.cell4.data [1], _43100_);
  and (_05322_, _00088_, _00087_);
  or (_00089_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00090_, \oc8051_gm_cxrom_1.cell4.data [2], _00074_);
  nand (_00091_, _00090_, _00089_);
  nand (_00092_, _00091_, _43100_);
  or (_00093_, \oc8051_gm_cxrom_1.cell4.data [2], _43100_);
  and (_05326_, _00093_, _00092_);
  or (_00094_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00095_, \oc8051_gm_cxrom_1.cell4.data [3], _00074_);
  nand (_00096_, _00095_, _00094_);
  nand (_00097_, _00096_, _43100_);
  or (_00098_, \oc8051_gm_cxrom_1.cell4.data [3], _43100_);
  and (_05329_, _00098_, _00097_);
  or (_00099_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00100_, \oc8051_gm_cxrom_1.cell4.data [4], _00074_);
  nand (_00101_, _00100_, _00099_);
  nand (_00102_, _00101_, _43100_);
  or (_00103_, \oc8051_gm_cxrom_1.cell4.data [4], _43100_);
  and (_05333_, _00103_, _00102_);
  or (_00104_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00105_, \oc8051_gm_cxrom_1.cell4.data [5], _00074_);
  nand (_00106_, _00105_, _00104_);
  nand (_00107_, _00106_, _43100_);
  or (_00108_, \oc8051_gm_cxrom_1.cell4.data [5], _43100_);
  and (_05337_, _00108_, _00107_);
  or (_00109_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00110_, \oc8051_gm_cxrom_1.cell4.data [6], _00074_);
  nand (_00111_, _00110_, _00109_);
  nand (_00112_, _00111_, _43100_);
  or (_00113_, \oc8051_gm_cxrom_1.cell4.data [6], _43100_);
  and (_05341_, _00113_, _00112_);
  or (_00114_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_00115_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_00116_, _00115_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_00117_, _00116_, _00114_);
  nand (_00118_, _00117_, _43100_);
  or (_00119_, \oc8051_gm_cxrom_1.cell5.data [7], _43100_);
  and (_05363_, _00119_, _00118_);
  or (_00120_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00121_, \oc8051_gm_cxrom_1.cell5.data [0], _00115_);
  nand (_00122_, _00121_, _00120_);
  nand (_00123_, _00122_, _43100_);
  or (_00124_, \oc8051_gm_cxrom_1.cell5.data [0], _43100_);
  and (_05369_, _00124_, _00123_);
  or (_00125_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00126_, \oc8051_gm_cxrom_1.cell5.data [1], _00115_);
  nand (_00127_, _00126_, _00125_);
  nand (_00128_, _00127_, _43100_);
  or (_00129_, \oc8051_gm_cxrom_1.cell5.data [1], _43100_);
  and (_05373_, _00129_, _00128_);
  or (_00130_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00132_, \oc8051_gm_cxrom_1.cell5.data [2], _00115_);
  nand (_00134_, _00132_, _00130_);
  nand (_00136_, _00134_, _43100_);
  or (_00138_, \oc8051_gm_cxrom_1.cell5.data [2], _43100_);
  and (_05377_, _00138_, _00136_);
  or (_00141_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00143_, \oc8051_gm_cxrom_1.cell5.data [3], _00115_);
  nand (_00145_, _00143_, _00141_);
  nand (_00147_, _00145_, _43100_);
  or (_00149_, \oc8051_gm_cxrom_1.cell5.data [3], _43100_);
  and (_05381_, _00149_, _00147_);
  or (_00152_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00154_, \oc8051_gm_cxrom_1.cell5.data [4], _00115_);
  nand (_00156_, _00154_, _00152_);
  nand (_00158_, _00156_, _43100_);
  or (_00160_, \oc8051_gm_cxrom_1.cell5.data [4], _43100_);
  and (_05385_, _00160_, _00158_);
  or (_00163_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00165_, \oc8051_gm_cxrom_1.cell5.data [5], _00115_);
  nand (_00167_, _00165_, _00163_);
  nand (_00169_, _00167_, _43100_);
  or (_00171_, \oc8051_gm_cxrom_1.cell5.data [5], _43100_);
  and (_05389_, _00171_, _00169_);
  or (_00174_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00176_, \oc8051_gm_cxrom_1.cell5.data [6], _00115_);
  nand (_00178_, _00176_, _00174_);
  nand (_00180_, _00178_, _43100_);
  or (_00182_, \oc8051_gm_cxrom_1.cell5.data [6], _43100_);
  and (_05393_, _00182_, _00180_);
  or (_00185_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_00187_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_00188_, _00187_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_00189_, _00188_, _00185_);
  nand (_00190_, _00189_, _43100_);
  or (_00191_, \oc8051_gm_cxrom_1.cell6.data [7], _43100_);
  and (_05414_, _00191_, _00190_);
  or (_00192_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00193_, \oc8051_gm_cxrom_1.cell6.data [0], _00187_);
  nand (_00194_, _00193_, _00192_);
  nand (_00195_, _00194_, _43100_);
  or (_00196_, \oc8051_gm_cxrom_1.cell6.data [0], _43100_);
  and (_05421_, _00196_, _00195_);
  or (_00197_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00198_, \oc8051_gm_cxrom_1.cell6.data [1], _00187_);
  nand (_00199_, _00198_, _00197_);
  nand (_00200_, _00199_, _43100_);
  or (_00201_, \oc8051_gm_cxrom_1.cell6.data [1], _43100_);
  and (_05425_, _00201_, _00200_);
  or (_00202_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00203_, \oc8051_gm_cxrom_1.cell6.data [2], _00187_);
  nand (_00204_, _00203_, _00202_);
  nand (_00205_, _00204_, _43100_);
  or (_00206_, \oc8051_gm_cxrom_1.cell6.data [2], _43100_);
  and (_05429_, _00206_, _00205_);
  or (_00207_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00208_, \oc8051_gm_cxrom_1.cell6.data [3], _00187_);
  nand (_00209_, _00208_, _00207_);
  nand (_00210_, _00209_, _43100_);
  or (_00211_, \oc8051_gm_cxrom_1.cell6.data [3], _43100_);
  and (_05433_, _00211_, _00210_);
  or (_00212_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00213_, \oc8051_gm_cxrom_1.cell6.data [4], _00187_);
  nand (_00214_, _00213_, _00212_);
  nand (_00215_, _00214_, _43100_);
  or (_00216_, \oc8051_gm_cxrom_1.cell6.data [4], _43100_);
  and (_05437_, _00216_, _00215_);
  or (_00217_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00218_, \oc8051_gm_cxrom_1.cell6.data [5], _00187_);
  nand (_00219_, _00218_, _00217_);
  nand (_00220_, _00219_, _43100_);
  or (_00221_, \oc8051_gm_cxrom_1.cell6.data [5], _43100_);
  and (_05441_, _00221_, _00220_);
  or (_00222_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00223_, \oc8051_gm_cxrom_1.cell6.data [6], _00187_);
  nand (_00224_, _00223_, _00222_);
  nand (_00225_, _00224_, _43100_);
  or (_00226_, \oc8051_gm_cxrom_1.cell6.data [6], _43100_);
  and (_05445_, _00226_, _00225_);
  or (_00227_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_00228_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_00229_, _00228_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_00230_, _00229_, _00227_);
  nand (_00231_, _00230_, _43100_);
  or (_00232_, \oc8051_gm_cxrom_1.cell7.data [7], _43100_);
  and (_05467_, _00232_, _00231_);
  or (_00233_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00234_, \oc8051_gm_cxrom_1.cell7.data [0], _00228_);
  nand (_00235_, _00234_, _00233_);
  nand (_00236_, _00235_, _43100_);
  or (_00237_, \oc8051_gm_cxrom_1.cell7.data [0], _43100_);
  and (_05474_, _00237_, _00236_);
  or (_00238_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00239_, \oc8051_gm_cxrom_1.cell7.data [1], _00228_);
  nand (_00240_, _00239_, _00238_);
  nand (_00241_, _00240_, _43100_);
  or (_00242_, \oc8051_gm_cxrom_1.cell7.data [1], _43100_);
  and (_05478_, _00242_, _00241_);
  or (_00243_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00244_, \oc8051_gm_cxrom_1.cell7.data [2], _00228_);
  nand (_00245_, _00244_, _00243_);
  nand (_00246_, _00245_, _43100_);
  or (_00247_, \oc8051_gm_cxrom_1.cell7.data [2], _43100_);
  and (_05482_, _00247_, _00246_);
  or (_00248_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00249_, \oc8051_gm_cxrom_1.cell7.data [3], _00228_);
  nand (_00250_, _00249_, _00248_);
  nand (_00251_, _00250_, _43100_);
  or (_00252_, \oc8051_gm_cxrom_1.cell7.data [3], _43100_);
  and (_05486_, _00252_, _00251_);
  or (_00253_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00254_, \oc8051_gm_cxrom_1.cell7.data [4], _00228_);
  nand (_00255_, _00254_, _00253_);
  nand (_00256_, _00255_, _43100_);
  or (_00257_, \oc8051_gm_cxrom_1.cell7.data [4], _43100_);
  and (_05490_, _00257_, _00256_);
  or (_00258_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00259_, \oc8051_gm_cxrom_1.cell7.data [5], _00228_);
  nand (_00260_, _00259_, _00258_);
  nand (_00261_, _00260_, _43100_);
  or (_00262_, \oc8051_gm_cxrom_1.cell7.data [5], _43100_);
  and (_05494_, _00262_, _00261_);
  or (_00263_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00264_, \oc8051_gm_cxrom_1.cell7.data [6], _00228_);
  nand (_00265_, _00264_, _00263_);
  nand (_00266_, _00265_, _43100_);
  or (_00267_, \oc8051_gm_cxrom_1.cell7.data [6], _43100_);
  and (_05498_, _00267_, _00266_);
  or (_00268_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_00269_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_00270_, _00269_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_00271_, _00270_, _00268_);
  nand (_00272_, _00271_, _43100_);
  or (_00273_, \oc8051_gm_cxrom_1.cell8.data [7], _43100_);
  and (_05520_, _00273_, _00272_);
  or (_00274_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00275_, \oc8051_gm_cxrom_1.cell8.data [0], _00269_);
  nand (_00276_, _00275_, _00274_);
  nand (_00277_, _00276_, _43100_);
  or (_00278_, \oc8051_gm_cxrom_1.cell8.data [0], _43100_);
  and (_05527_, _00278_, _00277_);
  or (_00279_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00280_, \oc8051_gm_cxrom_1.cell8.data [1], _00269_);
  nand (_00281_, _00280_, _00279_);
  nand (_00282_, _00281_, _43100_);
  or (_00283_, \oc8051_gm_cxrom_1.cell8.data [1], _43100_);
  and (_05531_, _00283_, _00282_);
  or (_00284_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00285_, \oc8051_gm_cxrom_1.cell8.data [2], _00269_);
  nand (_00286_, _00285_, _00284_);
  nand (_00287_, _00286_, _43100_);
  or (_00288_, \oc8051_gm_cxrom_1.cell8.data [2], _43100_);
  and (_05535_, _00288_, _00287_);
  or (_00289_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00290_, \oc8051_gm_cxrom_1.cell8.data [3], _00269_);
  nand (_00291_, _00290_, _00289_);
  nand (_00292_, _00291_, _43100_);
  or (_00293_, \oc8051_gm_cxrom_1.cell8.data [3], _43100_);
  and (_05539_, _00293_, _00292_);
  or (_00294_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00295_, \oc8051_gm_cxrom_1.cell8.data [4], _00269_);
  nand (_00296_, _00295_, _00294_);
  nand (_00297_, _00296_, _43100_);
  or (_00298_, \oc8051_gm_cxrom_1.cell8.data [4], _43100_);
  and (_05543_, _00298_, _00297_);
  or (_00299_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00300_, \oc8051_gm_cxrom_1.cell8.data [5], _00269_);
  nand (_00301_, _00300_, _00299_);
  nand (_00302_, _00301_, _43100_);
  or (_00303_, \oc8051_gm_cxrom_1.cell8.data [5], _43100_);
  and (_05547_, _00303_, _00302_);
  or (_00304_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00305_, \oc8051_gm_cxrom_1.cell8.data [6], _00269_);
  nand (_00306_, _00305_, _00304_);
  nand (_00307_, _00306_, _43100_);
  or (_00308_, \oc8051_gm_cxrom_1.cell8.data [6], _43100_);
  and (_05551_, _00308_, _00307_);
  or (_00309_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_00310_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_00311_, _00310_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_00312_, _00311_, _00309_);
  nand (_00313_, _00312_, _43100_);
  or (_00314_, \oc8051_gm_cxrom_1.cell9.data [7], _43100_);
  and (_05573_, _00314_, _00313_);
  or (_00315_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00316_, \oc8051_gm_cxrom_1.cell9.data [0], _00310_);
  nand (_00317_, _00316_, _00315_);
  nand (_00318_, _00317_, _43100_);
  or (_00319_, \oc8051_gm_cxrom_1.cell9.data [0], _43100_);
  and (_05580_, _00319_, _00318_);
  or (_00320_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00321_, \oc8051_gm_cxrom_1.cell9.data [1], _00310_);
  nand (_00322_, _00321_, _00320_);
  nand (_00323_, _00322_, _43100_);
  or (_00324_, \oc8051_gm_cxrom_1.cell9.data [1], _43100_);
  and (_05584_, _00324_, _00323_);
  or (_00325_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00326_, \oc8051_gm_cxrom_1.cell9.data [2], _00310_);
  nand (_00327_, _00326_, _00325_);
  nand (_00328_, _00327_, _43100_);
  or (_00329_, \oc8051_gm_cxrom_1.cell9.data [2], _43100_);
  and (_05588_, _00329_, _00328_);
  or (_00330_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00331_, \oc8051_gm_cxrom_1.cell9.data [3], _00310_);
  nand (_00332_, _00331_, _00330_);
  nand (_00333_, _00332_, _43100_);
  or (_00334_, \oc8051_gm_cxrom_1.cell9.data [3], _43100_);
  and (_05592_, _00334_, _00333_);
  or (_00335_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00336_, \oc8051_gm_cxrom_1.cell9.data [4], _00310_);
  nand (_00337_, _00336_, _00335_);
  nand (_00338_, _00337_, _43100_);
  or (_00339_, \oc8051_gm_cxrom_1.cell9.data [4], _43100_);
  and (_05596_, _00339_, _00338_);
  or (_00340_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00341_, \oc8051_gm_cxrom_1.cell9.data [5], _00310_);
  nand (_00342_, _00341_, _00340_);
  nand (_00343_, _00342_, _43100_);
  or (_00344_, \oc8051_gm_cxrom_1.cell9.data [5], _43100_);
  and (_05600_, _00344_, _00343_);
  or (_00345_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00346_, \oc8051_gm_cxrom_1.cell9.data [6], _00310_);
  nand (_00347_, _00346_, _00345_);
  nand (_00348_, _00347_, _43100_);
  or (_00349_, \oc8051_gm_cxrom_1.cell9.data [6], _43100_);
  and (_05604_, _00349_, _00348_);
  or (_00350_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_00351_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_00352_, _00351_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_00353_, _00352_, _00350_);
  nand (_00354_, _00353_, _43100_);
  or (_00355_, \oc8051_gm_cxrom_1.cell10.data [7], _43100_);
  and (_05626_, _00355_, _00354_);
  or (_00356_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00357_, \oc8051_gm_cxrom_1.cell10.data [0], _00351_);
  nand (_00358_, _00357_, _00356_);
  nand (_00359_, _00358_, _43100_);
  or (_00360_, \oc8051_gm_cxrom_1.cell10.data [0], _43100_);
  and (_05633_, _00360_, _00359_);
  or (_00361_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00362_, \oc8051_gm_cxrom_1.cell10.data [1], _00351_);
  nand (_00363_, _00362_, _00361_);
  nand (_00364_, _00363_, _43100_);
  or (_00365_, \oc8051_gm_cxrom_1.cell10.data [1], _43100_);
  and (_05637_, _00365_, _00364_);
  or (_00366_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00367_, \oc8051_gm_cxrom_1.cell10.data [2], _00351_);
  nand (_00368_, _00367_, _00366_);
  nand (_00369_, _00368_, _43100_);
  or (_00370_, \oc8051_gm_cxrom_1.cell10.data [2], _43100_);
  and (_05641_, _00370_, _00369_);
  or (_00371_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00372_, \oc8051_gm_cxrom_1.cell10.data [3], _00351_);
  nand (_00373_, _00372_, _00371_);
  nand (_00374_, _00373_, _43100_);
  or (_00375_, \oc8051_gm_cxrom_1.cell10.data [3], _43100_);
  and (_05645_, _00375_, _00374_);
  or (_00376_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00377_, \oc8051_gm_cxrom_1.cell10.data [4], _00351_);
  nand (_00378_, _00377_, _00376_);
  nand (_00379_, _00378_, _43100_);
  or (_00380_, \oc8051_gm_cxrom_1.cell10.data [4], _43100_);
  and (_05649_, _00380_, _00379_);
  or (_00381_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00382_, \oc8051_gm_cxrom_1.cell10.data [5], _00351_);
  nand (_00383_, _00382_, _00381_);
  nand (_00384_, _00383_, _43100_);
  or (_00385_, \oc8051_gm_cxrom_1.cell10.data [5], _43100_);
  and (_05653_, _00385_, _00384_);
  or (_00386_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00387_, \oc8051_gm_cxrom_1.cell10.data [6], _00351_);
  nand (_00388_, _00387_, _00386_);
  nand (_00389_, _00388_, _43100_);
  or (_00390_, \oc8051_gm_cxrom_1.cell10.data [6], _43100_);
  and (_05657_, _00390_, _00389_);
  or (_00391_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_00392_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_00393_, _00392_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_00394_, _00393_, _00391_);
  nand (_00395_, _00394_, _43100_);
  or (_00396_, \oc8051_gm_cxrom_1.cell11.data [7], _43100_);
  and (_05679_, _00396_, _00395_);
  or (_00397_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00398_, \oc8051_gm_cxrom_1.cell11.data [0], _00392_);
  nand (_00399_, _00398_, _00397_);
  nand (_00400_, _00399_, _43100_);
  or (_00401_, \oc8051_gm_cxrom_1.cell11.data [0], _43100_);
  and (_05686_, _00401_, _00400_);
  or (_00402_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00403_, \oc8051_gm_cxrom_1.cell11.data [1], _00392_);
  nand (_00404_, _00403_, _00402_);
  nand (_00405_, _00404_, _43100_);
  or (_00406_, \oc8051_gm_cxrom_1.cell11.data [1], _43100_);
  and (_05690_, _00406_, _00405_);
  or (_00407_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00408_, \oc8051_gm_cxrom_1.cell11.data [2], _00392_);
  nand (_00409_, _00408_, _00407_);
  nand (_00410_, _00409_, _43100_);
  or (_00411_, \oc8051_gm_cxrom_1.cell11.data [2], _43100_);
  and (_05694_, _00411_, _00410_);
  or (_00412_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00413_, \oc8051_gm_cxrom_1.cell11.data [3], _00392_);
  nand (_00414_, _00413_, _00412_);
  nand (_00415_, _00414_, _43100_);
  or (_00416_, \oc8051_gm_cxrom_1.cell11.data [3], _43100_);
  and (_05698_, _00416_, _00415_);
  or (_00417_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00418_, \oc8051_gm_cxrom_1.cell11.data [4], _00392_);
  nand (_00419_, _00418_, _00417_);
  nand (_00420_, _00419_, _43100_);
  or (_00421_, \oc8051_gm_cxrom_1.cell11.data [4], _43100_);
  and (_05702_, _00421_, _00420_);
  or (_00422_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00423_, \oc8051_gm_cxrom_1.cell11.data [5], _00392_);
  nand (_00424_, _00423_, _00422_);
  nand (_00425_, _00424_, _43100_);
  or (_00426_, \oc8051_gm_cxrom_1.cell11.data [5], _43100_);
  and (_05706_, _00426_, _00425_);
  or (_00427_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00428_, \oc8051_gm_cxrom_1.cell11.data [6], _00392_);
  nand (_00429_, _00428_, _00427_);
  nand (_00430_, _00429_, _43100_);
  or (_00431_, \oc8051_gm_cxrom_1.cell11.data [6], _43100_);
  and (_05710_, _00431_, _00430_);
  or (_00432_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_00433_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_00434_, _00433_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_00435_, _00434_, _00432_);
  nand (_00436_, _00435_, _43100_);
  or (_00437_, \oc8051_gm_cxrom_1.cell12.data [7], _43100_);
  and (_05732_, _00437_, _00436_);
  or (_00438_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00439_, \oc8051_gm_cxrom_1.cell12.data [0], _00433_);
  nand (_00440_, _00439_, _00438_);
  nand (_00441_, _00440_, _43100_);
  or (_00442_, \oc8051_gm_cxrom_1.cell12.data [0], _43100_);
  and (_05739_, _00442_, _00441_);
  or (_00443_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00444_, \oc8051_gm_cxrom_1.cell12.data [1], _00433_);
  nand (_00445_, _00444_, _00443_);
  nand (_00446_, _00445_, _43100_);
  or (_00447_, \oc8051_gm_cxrom_1.cell12.data [1], _43100_);
  and (_05743_, _00447_, _00446_);
  or (_00448_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00449_, \oc8051_gm_cxrom_1.cell12.data [2], _00433_);
  nand (_00450_, _00449_, _00448_);
  nand (_00451_, _00450_, _43100_);
  or (_00452_, \oc8051_gm_cxrom_1.cell12.data [2], _43100_);
  and (_05747_, _00452_, _00451_);
  or (_00453_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00454_, \oc8051_gm_cxrom_1.cell12.data [3], _00433_);
  nand (_00455_, _00454_, _00453_);
  nand (_00456_, _00455_, _43100_);
  or (_00457_, \oc8051_gm_cxrom_1.cell12.data [3], _43100_);
  and (_05751_, _00457_, _00456_);
  or (_00458_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00459_, \oc8051_gm_cxrom_1.cell12.data [4], _00433_);
  nand (_00460_, _00459_, _00458_);
  nand (_00461_, _00460_, _43100_);
  or (_00462_, \oc8051_gm_cxrom_1.cell12.data [4], _43100_);
  and (_05755_, _00462_, _00461_);
  or (_00463_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00464_, \oc8051_gm_cxrom_1.cell12.data [5], _00433_);
  nand (_00465_, _00464_, _00463_);
  nand (_00466_, _00465_, _43100_);
  or (_00467_, \oc8051_gm_cxrom_1.cell12.data [5], _43100_);
  and (_05759_, _00467_, _00466_);
  or (_00468_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00469_, \oc8051_gm_cxrom_1.cell12.data [6], _00433_);
  nand (_00470_, _00469_, _00468_);
  nand (_00471_, _00470_, _43100_);
  or (_00472_, \oc8051_gm_cxrom_1.cell12.data [6], _43100_);
  and (_05763_, _00472_, _00471_);
  or (_00473_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_00474_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_00475_, _00474_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_00476_, _00475_, _00473_);
  nand (_00477_, _00476_, _43100_);
  or (_00478_, \oc8051_gm_cxrom_1.cell13.data [7], _43100_);
  and (_05785_, _00478_, _00477_);
  or (_00479_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00480_, \oc8051_gm_cxrom_1.cell13.data [0], _00474_);
  nand (_00481_, _00480_, _00479_);
  nand (_00482_, _00481_, _43100_);
  or (_00483_, \oc8051_gm_cxrom_1.cell13.data [0], _43100_);
  and (_05792_, _00483_, _00482_);
  or (_00484_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00485_, \oc8051_gm_cxrom_1.cell13.data [1], _00474_);
  nand (_00486_, _00485_, _00484_);
  nand (_00487_, _00486_, _43100_);
  or (_00488_, \oc8051_gm_cxrom_1.cell13.data [1], _43100_);
  and (_05796_, _00488_, _00487_);
  or (_00489_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00490_, \oc8051_gm_cxrom_1.cell13.data [2], _00474_);
  nand (_00491_, _00490_, _00489_);
  nand (_00492_, _00491_, _43100_);
  or (_00493_, \oc8051_gm_cxrom_1.cell13.data [2], _43100_);
  and (_05800_, _00493_, _00492_);
  or (_00494_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00495_, \oc8051_gm_cxrom_1.cell13.data [3], _00474_);
  nand (_00496_, _00495_, _00494_);
  nand (_00497_, _00496_, _43100_);
  or (_00498_, \oc8051_gm_cxrom_1.cell13.data [3], _43100_);
  and (_05804_, _00498_, _00497_);
  or (_00499_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00500_, \oc8051_gm_cxrom_1.cell13.data [4], _00474_);
  nand (_00501_, _00500_, _00499_);
  nand (_00502_, _00501_, _43100_);
  or (_00503_, \oc8051_gm_cxrom_1.cell13.data [4], _43100_);
  and (_05808_, _00503_, _00502_);
  or (_00504_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00505_, \oc8051_gm_cxrom_1.cell13.data [5], _00474_);
  nand (_00506_, _00505_, _00504_);
  nand (_00507_, _00506_, _43100_);
  or (_00508_, \oc8051_gm_cxrom_1.cell13.data [5], _43100_);
  and (_05812_, _00508_, _00507_);
  or (_00509_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00510_, \oc8051_gm_cxrom_1.cell13.data [6], _00474_);
  nand (_00511_, _00510_, _00509_);
  nand (_00512_, _00511_, _43100_);
  or (_00513_, \oc8051_gm_cxrom_1.cell13.data [6], _43100_);
  and (_05816_, _00513_, _00512_);
  or (_00514_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_00515_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_00516_, _00515_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_00517_, _00516_, _00514_);
  nand (_00518_, _00517_, _43100_);
  or (_00519_, \oc8051_gm_cxrom_1.cell14.data [7], _43100_);
  and (_05838_, _00519_, _00518_);
  or (_00520_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00521_, \oc8051_gm_cxrom_1.cell14.data [0], _00515_);
  nand (_00522_, _00521_, _00520_);
  nand (_00523_, _00522_, _43100_);
  or (_00524_, \oc8051_gm_cxrom_1.cell14.data [0], _43100_);
  and (_05845_, _00524_, _00523_);
  or (_00525_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00526_, \oc8051_gm_cxrom_1.cell14.data [1], _00515_);
  nand (_00527_, _00526_, _00525_);
  nand (_00528_, _00527_, _43100_);
  or (_00529_, \oc8051_gm_cxrom_1.cell14.data [1], _43100_);
  and (_05849_, _00529_, _00528_);
  or (_00530_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00531_, \oc8051_gm_cxrom_1.cell14.data [2], _00515_);
  nand (_00532_, _00531_, _00530_);
  nand (_00533_, _00532_, _43100_);
  or (_00534_, \oc8051_gm_cxrom_1.cell14.data [2], _43100_);
  and (_05853_, _00534_, _00533_);
  or (_00535_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00536_, \oc8051_gm_cxrom_1.cell14.data [3], _00515_);
  nand (_00537_, _00536_, _00535_);
  nand (_00538_, _00537_, _43100_);
  or (_00539_, \oc8051_gm_cxrom_1.cell14.data [3], _43100_);
  and (_05857_, _00539_, _00538_);
  or (_00540_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00541_, \oc8051_gm_cxrom_1.cell14.data [4], _00515_);
  nand (_00542_, _00541_, _00540_);
  nand (_00543_, _00542_, _43100_);
  or (_00545_, \oc8051_gm_cxrom_1.cell14.data [4], _43100_);
  and (_05861_, _00545_, _00543_);
  or (_00547_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00548_, \oc8051_gm_cxrom_1.cell14.data [5], _00515_);
  nand (_00550_, _00548_, _00547_);
  nand (_00551_, _00550_, _43100_);
  or (_00553_, \oc8051_gm_cxrom_1.cell14.data [5], _43100_);
  and (_05865_, _00553_, _00551_);
  or (_00555_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00556_, \oc8051_gm_cxrom_1.cell14.data [6], _00515_);
  nand (_00558_, _00556_, _00555_);
  nand (_00559_, _00558_, _43100_);
  or (_00561_, \oc8051_gm_cxrom_1.cell14.data [6], _43100_);
  and (_05869_, _00561_, _00559_);
  or (_00563_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_00564_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_00566_, _00564_, \oc8051_gm_cxrom_1.cell15.data [7]);
  and (_00567_, _00566_, _00563_);
  or (_00569_, _00567_, rst);
  or (_00570_, \oc8051_gm_cxrom_1.cell15.data [7], _43100_);
  and (_05891_, _00570_, _00569_);
  or (_00572_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00574_, \oc8051_gm_cxrom_1.cell15.data [0], _00564_);
  and (_00575_, _00574_, _00572_);
  or (_00577_, _00575_, rst);
  or (_00578_, \oc8051_gm_cxrom_1.cell15.data [0], _43100_);
  and (_05898_, _00578_, _00577_);
  or (_00580_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00582_, \oc8051_gm_cxrom_1.cell15.data [1], _00564_);
  and (_00583_, _00582_, _00580_);
  or (_00585_, _00583_, rst);
  or (_00586_, \oc8051_gm_cxrom_1.cell15.data [1], _43100_);
  and (_05902_, _00586_, _00585_);
  or (_00588_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00590_, \oc8051_gm_cxrom_1.cell15.data [2], _00564_);
  and (_00591_, _00590_, _00588_);
  or (_00593_, _00591_, rst);
  or (_00594_, \oc8051_gm_cxrom_1.cell15.data [2], _43100_);
  and (_05906_, _00594_, _00593_);
  or (_00595_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00596_, \oc8051_gm_cxrom_1.cell15.data [3], _00564_);
  and (_00597_, _00596_, _00595_);
  or (_00598_, _00597_, rst);
  or (_00599_, \oc8051_gm_cxrom_1.cell15.data [3], _43100_);
  and (_05910_, _00599_, _00598_);
  or (_00600_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00601_, \oc8051_gm_cxrom_1.cell15.data [4], _00564_);
  and (_00602_, _00601_, _00600_);
  or (_00603_, _00602_, rst);
  or (_00604_, \oc8051_gm_cxrom_1.cell15.data [4], _43100_);
  and (_05914_, _00604_, _00603_);
  or (_00605_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00606_, \oc8051_gm_cxrom_1.cell15.data [5], _00564_);
  and (_00607_, _00606_, _00605_);
  or (_00608_, _00607_, rst);
  or (_00609_, \oc8051_gm_cxrom_1.cell15.data [5], _43100_);
  and (_05918_, _00609_, _00608_);
  or (_00610_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00611_, \oc8051_gm_cxrom_1.cell15.data [6], _00564_);
  and (_00612_, _00611_, _00610_);
  or (_00613_, _00612_, rst);
  or (_00614_, \oc8051_gm_cxrom_1.cell15.data [6], _43100_);
  and (_05922_, _00614_, _00613_);
  nor (_09697_, _38475_, rst);
  and (_00615_, _36509_, _43100_);
  nand (_00616_, _00615_, _38483_);
  nor (_00617_, _38467_, _38439_);
  or (_09700_, _00617_, _00616_);
  not (_00618_, _37164_);
  and (_00619_, _37654_, _37426_);
  and (_00620_, _00619_, _00618_);
  and (_00621_, _38215_, _38410_);
  and (_00622_, _00621_, _38432_);
  and (_00623_, _00622_, _37951_);
  and (_00624_, _00623_, _00620_);
  not (_00625_, _37426_);
  and (_00626_, _37654_, _00625_);
  not (_00627_, _36890_);
  not (_00628_, _38432_);
  nor (_00629_, _00628_, _38410_);
  not (_00630_, _37951_);
  nor (_00631_, _00630_, _38215_);
  and (_00632_, _00631_, _00629_);
  and (_00633_, _00632_, _00627_);
  and (_00634_, _00622_, _00630_);
  and (_00635_, _00634_, _37164_);
  or (_00636_, _00635_, _00633_);
  and (_00637_, _00636_, _00626_);
  or (_00638_, _00637_, _00624_);
  not (_00639_, _38215_);
  and (_00640_, _00629_, _00639_);
  and (_00641_, _00640_, _00630_);
  and (_00642_, _37164_, _36890_);
  nor (_00643_, _37654_, _37426_);
  and (_00644_, _00643_, _00642_);
  and (_00645_, _00644_, _00641_);
  and (_00646_, _00619_, _37164_);
  and (_00647_, _00646_, _00623_);
  or (_00648_, _00647_, _00645_);
  and (_00649_, _37164_, _00627_);
  and (_00650_, _00649_, _00626_);
  and (_00651_, _38432_, _38410_);
  and (_00652_, _00631_, _00651_);
  and (_00653_, _00652_, _00650_);
  not (_00654_, _00651_);
  nor (_00655_, _37164_, _00627_);
  and (_00656_, _00655_, _00626_);
  and (_00657_, _00656_, _00654_);
  or (_00658_, _00657_, _00653_);
  or (_00659_, _00658_, _00648_);
  not (_00660_, _00652_);
  nor (_00661_, _37164_, _36890_);
  and (_00662_, _00661_, _00619_);
  and (_00663_, _00642_, _00619_);
  nor (_00664_, _00663_, _00662_);
  nor (_00665_, _00664_, _00660_);
  and (_00666_, _00643_, _00618_);
  and (_00667_, _00627_, _38432_);
  and (_00668_, _00667_, _00621_);
  or (_00669_, _00668_, _00652_);
  and (_00670_, _00669_, _00666_);
  or (_00671_, _00670_, _00665_);
  or (_00672_, _00671_, _00659_);
  not (_00673_, _37654_);
  and (_00674_, _00673_, _37426_);
  and (_00675_, _00674_, _00661_);
  nor (_00676_, _00675_, _00630_);
  nor (_00677_, _00654_, _38215_);
  not (_00678_, _00677_);
  nor (_00679_, _00678_, _00676_);
  not (_00680_, _00679_);
  and (_00681_, _00655_, _00619_);
  and (_00682_, _00652_, _00681_);
  and (_00683_, _00674_, _00649_);
  and (_00684_, _00683_, _00652_);
  nor (_00685_, _00684_, _00682_);
  and (_00686_, _00685_, _00680_);
  and (_00687_, _36890_, _38432_);
  and (_00688_, _00687_, _00621_);
  and (_00689_, _00688_, _00666_);
  and (_00690_, _00644_, _00628_);
  or (_00691_, _00690_, _00689_);
  and (_00692_, _00674_, _00655_);
  and (_00693_, _00692_, _00634_);
  and (_00694_, _00674_, _36890_);
  and (_00695_, _00694_, _00652_);
  or (_00696_, _00695_, _00693_);
  nor (_00697_, _00696_, _00691_);
  nand (_00698_, _00697_, _00686_);
  or (_00699_, _00698_, _00672_);
  or (_00700_, _00699_, _00638_);
  and (_00701_, _00700_, _36520_);
  not (_00702_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_00703_, _36498_, _18201_);
  and (_00704_, _00703_, _38464_);
  nor (_00705_, _00704_, _00702_);
  or (_00706_, _00705_, rst);
  or (_09703_, _00706_, _00701_);
  nand (_00707_, _37426_, _36444_);
  or (_00708_, _36444_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_00709_, _00708_, _43100_);
  and (_09706_, _00709_, _00707_);
  and (_00710_, \oc8051_top_1.oc8051_sfr1.wait_data , _43100_);
  and (_00711_, _00710_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00712_, _38457_, _38484_);
  and (_00713_, _38440_, _38448_);
  and (_00714_, _00713_, _36967_);
  or (_00715_, _00714_, _00712_);
  and (_00716_, _38453_, _38467_);
  or (_00717_, _00716_, _38468_);
  or (_00718_, _00717_, _38543_);
  and (_00719_, _38520_, _38439_);
  and (_00720_, _38440_, _38517_);
  or (_00721_, _00720_, _00719_);
  nor (_00722_, _00721_, _00718_);
  nand (_00723_, _00722_, _38561_);
  or (_00724_, _00723_, _00715_);
  and (_00725_, _00724_, _00615_);
  or (_09709_, _00725_, _00711_);
  and (_00726_, _36967_, _38437_);
  and (_00727_, _00726_, _38516_);
  or (_00728_, _00727_, _38599_);
  not (_00729_, _38270_);
  and (_00730_, _00729_, _38455_);
  and (_00731_, _00730_, _38517_);
  or (_00732_, _00731_, _00728_);
  and (_00733_, _38467_, _38449_);
  or (_00734_, _00733_, _38441_);
  or (_00735_, _00734_, _00732_);
  and (_00736_, _00735_, _36509_);
  and (_00737_, _38570_, _00702_);
  not (_00738_, _38460_);
  and (_00739_, _00738_, _00737_);
  and (_00740_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00741_, _00740_, _00739_);
  or (_00742_, _00741_, _00736_);
  and (_09712_, _00742_, _43100_);
  and (_00743_, _00710_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_00744_, _38457_, _38508_);
  nor (_00745_, _38520_, _38508_);
  nor (_00746_, _00745_, _38490_);
  or (_00747_, _00746_, _00744_);
  and (_00748_, _00730_, _38530_);
  or (_00749_, _00748_, _00747_);
  nor (_00750_, _00745_, _38454_);
  and (_00751_, _36956_, _38437_);
  and (_00752_, _00751_, _38507_);
  nor (_00753_, _00752_, _00750_);
  not (_00754_, _00753_);
  and (_00755_, _38457_, _36956_);
  and (_00756_, _00755_, _37731_);
  and (_00757_, _38491_, _38437_);
  or (_00758_, _00757_, _38591_);
  or (_00759_, _00758_, _00756_);
  or (_00760_, _00759_, _00734_);
  or (_00761_, _00760_, _00754_);
  or (_00762_, _00761_, _00749_);
  and (_00763_, _00762_, _00615_);
  or (_09715_, _00763_, _00743_);
  and (_00764_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00765_, _38551_, _36509_);
  or (_00766_, _00765_, _00764_);
  or (_00767_, _00766_, _00739_);
  and (_09718_, _00767_, _43100_);
  and (_00768_, _38530_, _38504_);
  and (_00769_, _38438_, _38480_);
  and (_00770_, _00769_, _36956_);
  or (_00771_, _00770_, _00768_);
  or (_00772_, _00771_, _00714_);
  and (_00773_, _00771_, _38466_);
  or (_00774_, _00773_, _36455_);
  and (_00775_, _00774_, _00772_);
  not (_00776_, _38484_);
  nor (_00777_, _00617_, _00776_);
  nor (_00778_, _00777_, _00713_);
  not (_00779_, _00778_);
  and (_00780_, _00779_, _00737_);
  or (_00781_, _00780_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00782_, _00781_, _00775_);
  or (_00783_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18201_);
  and (_00784_, _00783_, _43100_);
  and (_09721_, _00784_, _00782_);
  and (_00785_, _00710_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_00786_, _00751_, _38516_);
  or (_00787_, _00752_, _00786_);
  or (_00788_, _38530_, _38517_);
  and (_00789_, _00788_, _38487_);
  or (_00790_, _00789_, _00787_);
  and (_00791_, _38504_, _37742_);
  or (_00792_, _00748_, _00719_);
  or (_00793_, _00792_, _00791_);
  or (_00794_, _00727_, _38518_);
  or (_00795_, _38441_, _38536_);
  or (_00796_, _00795_, _00794_);
  or (_00797_, _00796_, _00793_);
  or (_00798_, _00797_, _00790_);
  and (_00799_, _00798_, _00615_);
  or (_09724_, _00799_, _00785_);
  and (_00800_, _00710_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_00801_, _00730_, _38514_);
  and (_00802_, _38440_, _38496_);
  or (_00803_, _00802_, _38532_);
  nor (_00804_, _00803_, _00801_);
  nand (_00805_, _00804_, _00753_);
  nor (_00806_, _37219_, _37720_);
  and (_00807_, _00806_, _38488_);
  or (_00808_, _00807_, _38603_);
  and (_00809_, _38520_, _38487_);
  or (_00810_, _00809_, _00808_);
  or (_00811_, _38535_, _38528_);
  and (_00812_, _38457_, _38527_);
  or (_00813_, _00812_, _00731_);
  or (_00814_, _00813_, _00811_);
  or (_00815_, _00814_, _00810_);
  or (_00816_, _00815_, _00805_);
  and (_00817_, _00726_, _00806_);
  and (_00818_, _00726_, _38444_);
  or (_00819_, _00818_, _00817_);
  nor (_00820_, _38589_, _38563_);
  nand (_00821_, _00820_, _38541_);
  or (_00822_, _00821_, _00819_);
  or (_00823_, _00822_, _00749_);
  or (_00824_, _00823_, _00816_);
  and (_00825_, _00824_, _00615_);
  or (_09727_, _00825_, _00800_);
  and (_00826_, _00730_, _38497_);
  or (_00827_, _00826_, _38600_);
  and (_00828_, _00751_, _38447_);
  and (_00829_, _00828_, _37470_);
  or (_00830_, _00829_, _38583_);
  and (_00831_, _38497_, _38437_);
  or (_00832_, _00831_, _00830_);
  or (_00833_, _00832_, _00827_);
  and (_00834_, _00730_, _38449_);
  or (_00835_, _00834_, _00833_);
  and (_00836_, _00835_, _36509_);
  nand (_00837_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_00838_, _00837_, _38472_);
  or (_00839_, _00838_, _00836_);
  and (_09730_, _00839_, _43100_);
  or (_00840_, _38521_, _38518_);
  not (_00841_, _38564_);
  or (_00842_, _00746_, _00841_);
  or (_00843_, _00842_, _00840_);
  and (_00844_, _37219_, _37709_);
  and (_00845_, _00844_, _36956_);
  and (_00846_, _00845_, _38481_);
  or (_00847_, _00846_, _38531_);
  or (_00848_, _00847_, _38528_);
  or (_00849_, _00848_, _00768_);
  nand (_00850_, _38552_, _38544_);
  or (_00851_, _00850_, _00849_);
  or (_00852_, _00851_, _00843_);
  and (_00853_, _00726_, _38448_);
  or (_00854_, _00853_, _00770_);
  and (_00855_, _00751_, _00844_);
  or (_00856_, _00855_, _38510_);
  or (_00857_, _00856_, _00728_);
  or (_00858_, _00857_, _00854_);
  and (_00859_, _00845_, _38487_);
  or (_00860_, _00859_, _38589_);
  or (_00861_, _00860_, _38489_);
  or (_00862_, _38586_, _38548_);
  or (_00863_, _00862_, _00861_);
  or (_00864_, _00863_, _00858_);
  or (_00865_, _00864_, _00754_);
  or (_00866_, _00865_, _00852_);
  and (_00867_, _00866_, _36509_);
  or (_00868_, _00773_, _00739_);
  and (_00869_, _38466_, _38559_);
  or (_00870_, _00869_, _00868_);
  and (_00871_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00872_, _00871_, _00870_);
  or (_00873_, _00872_, _00867_);
  and (_09733_, _00873_, _43100_);
  nor (_09792_, _38612_, rst);
  nor (_09794_, _38575_, rst);
  nand (_09797_, _00779_, _00615_);
  nand (_00874_, _00713_, _00615_);
  not (_00875_, _38467_);
  or (_00876_, _00616_, _00875_);
  and (_09800_, _00876_, _00874_);
  or (_00877_, _00638_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_00878_, _00877_, _00704_);
  nor (_00879_, _00703_, _38464_);
  or (_00880_, _00879_, rst);
  or (_09803_, _00880_, _00878_);
  nand (_00881_, _37951_, _36444_);
  or (_00882_, _36444_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_00883_, _00882_, _43100_);
  and (_09806_, _00883_, _00881_);
  not (_00884_, _36444_);
  or (_00885_, _38215_, _00884_);
  or (_00886_, _36444_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_00887_, _00886_, _43100_);
  and (_09809_, _00887_, _00885_);
  nand (_00888_, _38410_, _36444_);
  or (_00889_, _36444_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_00890_, _00889_, _43100_);
  and (_09812_, _00890_, _00888_);
  nand (_00891_, _38432_, _36444_);
  or (_00892_, _36444_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_00893_, _00892_, _43100_);
  and (_09815_, _00893_, _00891_);
  or (_00894_, _36890_, _00884_);
  or (_00895_, _36444_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_00896_, _00895_, _43100_);
  and (_09818_, _00896_, _00894_);
  nand (_00897_, _37164_, _36444_);
  or (_00898_, _36444_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_00899_, _00898_, _43100_);
  and (_09821_, _00899_, _00897_);
  nand (_00900_, _37654_, _36444_);
  or (_00901_, _36444_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_00902_, _00901_, _43100_);
  and (_09824_, _00902_, _00900_);
  or (_00903_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _18201_);
  and (_00904_, _00903_, _43100_);
  and (_00905_, _00904_, _00781_);
  and (_00906_, _38449_, _38487_);
  or (_00907_, _00826_, _00906_);
  and (_00908_, _00726_, _38499_);
  or (_00909_, _00834_, _00908_);
  or (_00910_, _00909_, _00907_);
  or (_00911_, _38441_, _38593_);
  or (_00912_, _00911_, _00910_);
  and (_00913_, _38499_, _38437_);
  and (_00914_, _00913_, _36956_);
  or (_00915_, _00914_, _00831_);
  or (_00916_, _38520_, _38507_);
  and (_00917_, _00916_, _38457_);
  or (_00918_, _00917_, _00915_);
  or (_00919_, _00918_, _00912_);
  and (_00920_, _00730_, _38500_);
  or (_00921_, _00920_, _00830_);
  and (_00922_, _38457_, _38445_);
  and (_00923_, _00730_, _38484_);
  or (_00924_, _00923_, _00922_);
  or (_00925_, _00924_, _00921_);
  or (_00926_, _00802_, _38603_);
  or (_00928_, _00818_, _00801_);
  or (_00929_, _00928_, _00926_);
  or (_00930_, _00929_, _00925_);
  or (_00931_, _00733_, _38540_);
  or (_00932_, _00931_, _00812_);
  and (_00933_, _38500_, _38487_);
  and (_00934_, _00726_, _38483_);
  and (_00935_, _00755_, _38483_);
  or (_00936_, _00935_, _00934_);
  or (_00937_, _00936_, _00933_);
  or (_00938_, _00937_, _00932_);
  or (_00939_, _00938_, _00930_);
  or (_00940_, _00939_, _00919_);
  and (_00941_, _00940_, _00615_);
  or (_09827_, _00941_, _00905_);
  and (_00942_, _00710_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not (_00943_, _38519_);
  or (_00944_, _00819_, _00943_);
  or (_00945_, _38527_, _38514_);
  and (_00946_, _00945_, _38504_);
  not (_00947_, _38457_);
  nor (_00948_, _00947_, _38501_);
  or (_00949_, _00948_, _00946_);
  or (_00950_, _00949_, _00944_);
  or (_00951_, _00932_, _00810_);
  and (_00952_, _38457_, _38514_);
  and (_00953_, _37219_, _37720_);
  and (_00954_, _00751_, _00953_);
  and (_00955_, _00954_, _37470_);
  nor (_00956_, _00955_, _38588_);
  not (_00958_, _00956_);
  or (_00959_, _00958_, _00756_);
  or (_00960_, _00959_, _00952_);
  or (_00961_, _00960_, _00715_);
  or (_00962_, _00961_, _00951_);
  or (_00963_, _00962_, _00950_);
  and (_00964_, _00963_, _00615_);
  or (_34277_, _00964_, _00942_);
  or (_00965_, _00862_, _00854_);
  or (_00966_, _00965_, _00852_);
  and (_00967_, _00966_, _36509_);
  and (_00968_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00969_, _00968_, _00870_);
  or (_00970_, _00969_, _00967_);
  and (_34279_, _00970_, _43100_);
  and (_00971_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00972_, _00971_, _00868_);
  and (_00973_, _00972_, _43100_);
  and (_00974_, _38562_, _36967_);
  or (_00975_, _00974_, _38599_);
  or (_00977_, _00975_, _00861_);
  or (_00978_, _00977_, _00771_);
  and (_00979_, _00978_, _00615_);
  or (_34282_, _00979_, _00973_);
  or (_00980_, _00713_, _38459_);
  and (_00981_, _00826_, _36956_);
  or (_00982_, _00981_, _00920_);
  or (_00983_, _00982_, _00980_);
  or (_00984_, _00830_, _38582_);
  or (_00985_, _00915_, _00802_);
  or (_00986_, _00985_, _00984_);
  or (_00987_, _00986_, _00983_);
  and (_00988_, _38457_, _38517_);
  or (_00989_, _00935_, _38458_);
  or (_00990_, _00989_, _00988_);
  and (_00991_, _00730_, _38491_);
  or (_00992_, _00991_, _00834_);
  or (_00993_, _00992_, _00712_);
  or (_00994_, _00993_, _00917_);
  or (_00995_, _00994_, _00990_);
  or (_00996_, _00855_, _00906_);
  or (_00997_, _00996_, _00859_);
  or (_00998_, _00812_, _38446_);
  or (_00999_, _00922_, _00952_);
  or (_01000_, _00999_, _00998_);
  or (_01001_, _01000_, _00997_);
  and (_01002_, _00826_, _36967_);
  and (_01003_, _38504_, _38500_);
  and (_01004_, _00846_, _37470_);
  or (_01005_, _01004_, _01003_);
  or (_01006_, _01005_, _01002_);
  or (_01007_, _01006_, _00771_);
  or (_01008_, _01007_, _01001_);
  or (_01009_, _01008_, _00995_);
  or (_01010_, _01009_, _00987_);
  and (_01011_, _01010_, _36509_);
  and (_01012_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01013_, _00780_, _38473_);
  or (_01014_, _01013_, _01012_);
  or (_01015_, _01014_, _01011_);
  and (_34284_, _01015_, _43100_);
  and (_01016_, _00859_, _37470_);
  or (_01017_, _38459_, _00906_);
  or (_01018_, _01017_, _38548_);
  or (_01019_, _01018_, _01016_);
  or (_01020_, _01019_, _00984_);
  or (_01021_, _01020_, _00985_);
  and (_01022_, _00751_, _38483_);
  or (_01023_, _00846_, _00733_);
  nor (_01024_, _01023_, _01022_);
  nand (_01025_, _01024_, _38451_);
  and (_01026_, _00945_, _38440_);
  or (_01027_, _01026_, _38502_);
  or (_01028_, _01027_, _01025_);
  or (_01029_, _01028_, _00995_);
  or (_01030_, _01029_, _01021_);
  and (_01031_, _01030_, _36509_);
  and (_01032_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01033_, _01032_, _01013_);
  or (_01034_, _01033_, _01031_);
  and (_34286_, _01034_, _43100_);
  and (_01035_, _00710_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not (_01036_, _42525_);
  or (_01037_, _00834_, _01036_);
  and (_01038_, _38440_, _38520_);
  and (_01039_, _38440_, _38507_);
  and (_01040_, _01039_, _36956_);
  or (_01041_, _01040_, _01038_);
  or (_01042_, _01041_, _00790_);
  or (_01043_, _01042_, _01037_);
  not (_01044_, _42524_);
  or (_01045_, _00795_, _01044_);
  and (_01046_, _38457_, _38520_);
  or (_01047_, _01046_, _00748_);
  or (_01048_, _01047_, _00840_);
  or (_01049_, _01048_, _01045_);
  or (_01050_, _00829_, _00727_);
  and (_01051_, _38581_, _38497_);
  and (_01052_, _38440_, _38491_);
  or (_01053_, _01052_, _01051_);
  or (_01054_, _01053_, _01050_);
  and (_01055_, _38554_, _38437_);
  or (_01056_, _01055_, _00906_);
  or (_01057_, _01056_, _38550_);
  and (_01058_, _38440_, _38554_);
  or (_01059_, _01058_, _00981_);
  or (_01060_, _01059_, _01057_);
  or (_01061_, _01060_, _01054_);
  or (_01062_, _01061_, _01049_);
  or (_01063_, _01062_, _01043_);
  and (_01064_, _01063_, _00615_);
  or (_34288_, _01064_, _01035_);
  or (_01065_, _00809_, _00807_);
  or (_01066_, _01065_, _01002_);
  or (_01067_, _01066_, _00814_);
  or (_01068_, _01067_, _00983_);
  or (_01069_, _01058_, _01046_);
  or (_01070_, _01040_, _00915_);
  or (_01071_, _01070_, _01069_);
  nand (_01072_, _38585_, _38549_);
  or (_01073_, _00817_, _38441_);
  or (_01074_, _38446_, _38540_);
  or (_01075_, _01074_, _01073_);
  or (_01076_, _01075_, _01072_);
  or (_01077_, _01076_, _01071_);
  or (_01078_, _01077_, _01068_);
  and (_01079_, _01078_, _00615_);
  and (_01080_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_01081_, _38459_, _36466_);
  or (_01082_, _01081_, _01080_);
  and (_01083_, _01082_, _43100_);
  or (_34290_, _01083_, _01079_);
  or (_01084_, _00933_, _00914_);
  nor (_01085_, _00757_, _38539_);
  nand (_01086_, _01085_, _38590_);
  or (_01087_, _01086_, _00993_);
  or (_01088_, _01087_, _01084_);
  nor (_01089_, _00920_, _38548_);
  not (_01090_, _01089_);
  nor (_01091_, _01090_, _38547_);
  or (_01092_, _00731_, _38602_);
  and (_01093_, _38440_, _38497_);
  or (_01094_, _01093_, _01050_);
  nor (_01095_, _01094_, _01092_);
  nand (_01096_, _01095_, _01091_);
  or (_01097_, _01096_, _01088_);
  or (_01098_, _00935_, _38542_);
  or (_01099_, _01098_, _01052_);
  or (_01100_, _01099_, _00754_);
  or (_01101_, _01100_, _00749_);
  or (_01102_, _01101_, _01097_);
  and (_01103_, _01102_, _36509_);
  and (_01104_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01105_, _01104_, _38470_);
  or (_01106_, _01105_, _01103_);
  and (_34292_, _01106_, _43100_);
  or (_01107_, _01047_, _00794_);
  or (_01108_, _01090_, _01084_);
  or (_01109_, _01108_, _01107_);
  or (_01110_, _38599_, _38589_);
  nor (_01111_, _01110_, _01039_);
  nand (_01112_, _01111_, _42525_);
  or (_01113_, _01112_, _00747_);
  or (_01114_, _01113_, _01109_);
  or (_01115_, _01114_, _01100_);
  and (_01116_, _01115_, _00615_);
  and (_01117_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01118_, _01117_, _38471_);
  and (_01119_, _01118_, _43100_);
  or (_34294_, _01119_, _01116_);
  and (_01120_, _00710_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_01121_, _00720_, _38522_);
  nand (_01122_, _01121_, _42524_);
  not (_01123_, _38438_);
  or (_01124_, _38440_, _01123_);
  and (_01125_, _01124_, _38491_);
  or (_01126_, _01125_, _01069_);
  or (_01127_, _01126_, _01122_);
  or (_01128_, _01041_, _00833_);
  or (_01129_, _01128_, _01037_);
  or (_01130_, _01129_, _01127_);
  and (_01131_, _01130_, _00615_);
  or (_34296_, _01131_, _01120_);
  nor (_39173_, _37426_, rst);
  nor (_39174_, _42516_, rst);
  and (_01132_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_01133_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_01134_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_01135_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_01136_, _01135_, _01134_);
  and (_01137_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01138_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_01139_, _01138_, _01137_);
  and (_01140_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_01141_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_01142_, _01141_, _01140_);
  and (_01143_, _01142_, _01139_);
  and (_01144_, _01143_, _01136_);
  nor (_01145_, _01144_, _36694_);
  nor (_01146_, _01145_, _01133_);
  nor (_01147_, _01146_, _42500_);
  nor (_01148_, _01147_, _01132_);
  nor (_39176_, _01148_, rst);
  nor (_39186_, _37951_, rst);
  and (_39188_, _38215_, _43100_);
  nor (_39189_, _38410_, rst);
  nor (_39190_, _38432_, rst);
  and (_39191_, _36890_, _43100_);
  nor (_39192_, _37164_, rst);
  nor (_39193_, _37654_, rst);
  nor (_39194_, _42682_, rst);
  nor (_39195_, _42611_, rst);
  nor (_39197_, _42803_, rst);
  nor (_39198_, _42646_, rst);
  nor (_39199_, _42551_, rst);
  nor (_39200_, _42777_, rst);
  nor (_39201_, _42739_, rst);
  and (_01149_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_01150_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_01151_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_01152_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_01153_, _01152_, _01151_);
  and (_01154_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_01155_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_01156_, _01155_, _01154_);
  and (_01157_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_01158_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_01159_, _01158_, _01157_);
  and (_01160_, _01159_, _01156_);
  and (_01161_, _01160_, _01153_);
  nor (_01162_, _01161_, _36694_);
  nor (_01163_, _01162_, _01150_);
  nor (_01164_, _01163_, _42500_);
  nor (_01165_, _01164_, _01149_);
  nor (_39203_, _01165_, rst);
  and (_01166_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_01167_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_01168_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_01169_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_01170_, _01169_, _01168_);
  and (_01171_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_01172_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_01173_, _01172_, _01171_);
  and (_01174_, _01173_, _01170_);
  and (_01175_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_01176_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_01177_, _01176_, _01175_);
  and (_01178_, _01177_, _01174_);
  nor (_01179_, _01178_, _36694_);
  nor (_01180_, _01179_, _01167_);
  nor (_01181_, _01180_, _42500_);
  nor (_01182_, _01181_, _01166_);
  nor (_39204_, _01182_, rst);
  and (_01183_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_01184_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_01185_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_01186_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01187_, _01186_, _01185_);
  and (_01188_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_01189_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_01190_, _01189_, _01188_);
  and (_01191_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_01192_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_01193_, _01192_, _01191_);
  and (_01194_, _01193_, _01190_);
  and (_01195_, _01194_, _01187_);
  nor (_01196_, _01195_, _36694_);
  nor (_01197_, _01196_, _01184_);
  nor (_01198_, _01197_, _42500_);
  nor (_01199_, _01198_, _01183_);
  nor (_39205_, _01199_, rst);
  and (_01200_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_01201_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_01202_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_01203_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_01204_, _01203_, _01202_);
  and (_01205_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_01206_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_01207_, _01206_, _01205_);
  and (_01208_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_01209_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_01210_, _01209_, _01208_);
  and (_01212_, _01210_, _01207_);
  and (_01214_, _01212_, _01204_);
  nor (_01216_, _01214_, _36694_);
  nor (_01218_, _01216_, _01201_);
  nor (_01220_, _01218_, _42500_);
  nor (_01222_, _01220_, _01200_);
  nor (_39206_, _01222_, rst);
  and (_01225_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_01227_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_01229_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_01231_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_01233_, _01231_, _01229_);
  and (_01235_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_01237_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_01239_, _01237_, _01235_);
  and (_01241_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_01243_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_01245_, _01243_, _01241_);
  and (_01247_, _01245_, _01239_);
  and (_01249_, _01247_, _01233_);
  nor (_01251_, _01249_, _36694_);
  nor (_01253_, _01251_, _01227_);
  nor (_01255_, _01253_, _42500_);
  nor (_01257_, _01255_, _01225_);
  nor (_39207_, _01257_, rst);
  and (_01260_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_01262_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_01264_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_01266_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_01268_, _01266_, _01264_);
  and (_01270_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_01272_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_01274_, _01272_, _01270_);
  and (_01276_, _01274_, _01268_);
  and (_01278_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_01280_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_01282_, _01280_, _01278_);
  and (_01284_, _01282_, _01276_);
  nor (_01286_, _01284_, _36694_);
  nor (_01288_, _01286_, _01262_);
  nor (_01290_, _01288_, _42500_);
  nor (_01292_, _01290_, _01260_);
  nor (_39209_, _01292_, rst);
  and (_01295_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_01297_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_01299_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_01301_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_01303_, _01301_, _01299_);
  and (_01305_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_01306_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_01307_, _01306_, _01305_);
  and (_01308_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_01309_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_01310_, _01309_, _01308_);
  and (_01311_, _01310_, _01307_);
  and (_01312_, _01311_, _01303_);
  nor (_01313_, _01312_, _36694_);
  nor (_01314_, _01313_, _01297_);
  nor (_01315_, _01314_, _42500_);
  nor (_01316_, _01315_, _01295_);
  nor (_39210_, _01316_, rst);
  and (_01317_, _36520_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_01318_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_01319_, _01317_, _38760_);
  and (_01320_, _01319_, _43100_);
  and (_39234_, _01320_, _01318_);
  not (_01321_, _01317_);
  or (_01322_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_01323_, _36520_, _43100_);
  and (_00000_, _01323_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _43100_);
  or (_01325_, _01324_, _00000_);
  and (_39235_, _01325_, _01322_);
  nor (_39273_, _42521_, rst);
  and (_39275_, _42559_, _43100_);
  and (_39276_, _42495_, _43100_);
  nor (_01326_, _38561_, _38570_);
  nor (_01327_, _42665_, _27650_);
  and (_01328_, _42665_, _27650_);
  nor (_01329_, _01328_, _01327_);
  nor (_01330_, _42579_, _27825_);
  and (_01331_, _42579_, _27825_);
  nor (_01332_, _01331_, _01330_);
  nor (_01333_, _01332_, _01329_);
  nor (_01334_, _42787_, _27343_);
  and (_01335_, _42787_, _27343_);
  nor (_01336_, _01335_, _01334_);
  nor (_01337_, _42743_, _27211_);
  and (_01338_, _42743_, _27211_);
  nor (_01339_, _01338_, _01337_);
  nor (_01340_, _01339_, _01336_);
  and (_01341_, _01340_, _01333_);
  and (_01342_, _01341_, _42858_);
  nor (_01343_, _31308_, _40112_);
  and (_01344_, _01343_, _01342_);
  and (_01345_, _01344_, _01326_);
  not (_01346_, _01345_);
  not (_01347_, _00786_);
  nor (_01348_, _00991_, _38536_);
  and (_01349_, _01348_, _01347_);
  and (_01350_, _01349_, _00956_);
  nor (_01351_, _01326_, _38469_);
  or (_01352_, _28571_, _28209_);
  nor (_01353_, _01352_, _28538_);
  and (_01354_, _01353_, _31460_);
  nand (_01355_, _01354_, _33725_);
  nor (_01356_, _01355_, _34573_);
  and (_01357_, _01356_, _01351_);
  and (_01358_, _01357_, _35748_);
  and (_01359_, _01358_, _29196_);
  not (_01360_, _01359_);
  and (_01361_, _01326_, _28944_);
  not (_01362_, _01361_);
  nor (_01363_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_01364_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01365_, _01364_, _01363_);
  nor (_01366_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_01367_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01368_, _01367_, _01366_);
  and (_01369_, _01368_, _01365_);
  and (_01370_, _01369_, _38610_);
  not (_01371_, _38469_);
  nor (_01372_, _01326_, _38498_);
  nor (_01373_, _01372_, _01371_);
  and (_01374_, _01373_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_01375_, _01374_, _01370_);
  and (_01376_, _01375_, _01362_);
  and (_01377_, _01376_, _01360_);
  not (_01378_, _38500_);
  nor (_01379_, _38554_, _38445_);
  and (_01380_, _01379_, _01378_);
  nor (_01381_, _01380_, _00875_);
  not (_01382_, _01381_);
  and (_01383_, _01382_, _01377_);
  and (_01384_, _01383_, _01350_);
  and (_01385_, _38468_, _36967_);
  or (_01386_, _01385_, _38559_);
  or (_01387_, _01386_, _01377_);
  nor (_01388_, _01387_, _38558_);
  or (_01389_, _01388_, _01384_);
  nor (_01390_, _00729_, _38414_);
  and (_01391_, _38006_, _38454_);
  and (_01392_, _01391_, _01390_);
  and (_01393_, _01392_, _38445_);
  nor (_01394_, _01393_, _00716_);
  and (_01395_, _01394_, _01389_);
  and (_01396_, _01395_, _38506_);
  nor (_01397_, _01396_, _42532_);
  and (_01398_, _38507_, _38504_);
  nor (_01399_, _01398_, _00769_);
  nor (_01400_, _01399_, _36466_);
  nor (_01401_, _01400_, _38572_);
  not (_01402_, _01401_);
  nor (_01403_, _01402_, _01397_);
  nor (_01404_, _39115_, _39106_);
  and (_01405_, _01404_, _39170_);
  not (_01406_, _01405_);
  and (_01407_, _01406_, _01373_);
  not (_01408_, _39409_);
  and (_01409_, _01408_, _38610_);
  nor (_01410_, _01409_, _01407_);
  not (_01411_, _01410_);
  nor (_01412_, _01411_, _01403_);
  nor (_01413_, _42617_, _26860_);
  and (_01414_, _42617_, _26860_);
  nor (_01415_, _01414_, _01413_);
  and (_01416_, _42701_, _32582_);
  nor (_01417_, _42701_, _32582_);
  or (_01418_, _01417_, _01416_);
  nor (_01419_, _01418_, _01415_);
  nor (_01420_, _42823_, _26740_);
  and (_01421_, _42823_, _26740_);
  nor (_01422_, _01421_, _01420_);
  nor (_01423_, _01422_, _39432_);
  and (_01424_, _01423_, _01419_);
  and (_01425_, _01424_, _01342_);
  nor (_01426_, _27496_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_01427_, _01426_, _01425_);
  not (_01428_, _01427_);
  and (_01429_, _01428_, _01412_);
  and (_01430_, _01429_, _01346_);
  nor (_01431_, _38572_, rst);
  and (_39280_, _01431_, _01430_);
  and (_39281_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _43100_);
  and (_39282_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _43100_);
  not (_01432_, _38572_);
  nor (_01433_, _01432_, _30574_);
  not (_01434_, _38845_);
  and (_01435_, _38446_, _38466_);
  and (_01436_, _01435_, _01434_);
  not (_01437_, _38468_);
  and (_01438_, _00956_, _38561_);
  and (_01439_, _01438_, _01437_);
  and (_01440_, _01439_, _01394_);
  and (_01441_, _01440_, _01349_);
  nor (_01442_, _01441_, _42532_);
  nor (_01443_, _01435_, _01400_);
  not (_01444_, _01443_);
  and (_01445_, _01438_, _01348_);
  nor (_01446_, _01445_, _42532_);
  and (_01447_, _01398_, _36455_);
  not (_01448_, _01447_);
  and (_01449_, _38467_, _38497_);
  and (_01450_, _01449_, _36455_);
  nor (_01451_, _01450_, _38572_);
  and (_01452_, _01451_, _01448_);
  not (_01453_, _01452_);
  nor (_01454_, _01453_, _01446_);
  nand (_01455_, _01454_, _01444_);
  nor (_01456_, _01455_, _01442_);
  and (_01457_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01458_, _01457_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01459_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01460_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01461_, _01460_, _01459_);
  and (_01462_, _01461_, _01458_);
  and (_01463_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01464_, _01463_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01465_, _01464_, _01462_);
  and (_01466_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01467_, _01466_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01468_, _01467_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01469_, _01468_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_01470_, _01469_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_01471_, _01469_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_01472_, _01471_, _01470_);
  and (_01473_, _01472_, _01456_);
  and (_01474_, _01447_, _42517_);
  or (_01475_, _01474_, _01473_);
  nor (_01476_, _01444_, _01442_);
  and (_01477_, _01476_, _01454_);
  and (_01478_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_01479_, _01478_, _01475_);
  nor (_01480_, _01479_, _01436_);
  nand (_01481_, _01480_, _01430_);
  or (_01482_, _01481_, _01433_);
  and (_01483_, _01454_, _42516_);
  not (_01484_, _01148_);
  nor (_01485_, _01454_, _01484_);
  nor (_01486_, _01485_, _01483_);
  and (_01487_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_01488_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01489_, _01454_, _42739_);
  not (_01490_, _01316_);
  nor (_01491_, _01454_, _01490_);
  nor (_01492_, _01491_, _01489_);
  and (_01493_, _01492_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_01494_, _01492_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_01495_, _01494_, _01493_);
  and (_01496_, _01454_, _42777_);
  not (_01497_, _01292_);
  nor (_01498_, _01454_, _01497_);
  nor (_01499_, _01498_, _01496_);
  and (_01500_, _01499_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_01501_, _01499_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_01502_, _01454_, _42551_);
  not (_01503_, _01257_);
  nor (_01504_, _01454_, _01503_);
  nor (_01505_, _01504_, _01502_);
  nand (_01506_, _01505_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01507_, _01454_, _42646_);
  not (_01508_, _01222_);
  nor (_01509_, _01454_, _01508_);
  nor (_01510_, _01509_, _01507_);
  and (_01511_, _01510_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_01512_, _01510_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01513_, _01454_, _42803_);
  not (_01514_, _01199_);
  nor (_01515_, _01454_, _01514_);
  nor (_01516_, _01515_, _01513_);
  and (_01517_, _01516_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01518_, _01454_, _42611_);
  not (_01519_, _01182_);
  nor (_01520_, _01454_, _01519_);
  nor (_01521_, _01520_, _01518_);
  and (_01522_, _01521_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01523_, _01454_, _42682_);
  not (_01524_, _01165_);
  nor (_01525_, _01454_, _01524_);
  nor (_01526_, _01525_, _01523_);
  and (_01527_, _01526_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_01528_, _01521_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_01529_, _01528_, _01522_);
  and (_01530_, _01529_, _01527_);
  nor (_01531_, _01530_, _01522_);
  not (_01532_, _01531_);
  nor (_01533_, _01516_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_01534_, _01533_, _01517_);
  and (_01535_, _01534_, _01532_);
  nor (_01536_, _01535_, _01517_);
  nor (_01537_, _01536_, _01512_);
  or (_01538_, _01537_, _01511_);
  or (_01539_, _01505_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01540_, _01539_, _01506_);
  nand (_01541_, _01540_, _01538_);
  and (_01542_, _01541_, _01506_);
  nor (_01543_, _01542_, _01501_);
  or (_01544_, _01543_, _01500_);
  and (_01545_, _01544_, _01495_);
  nor (_01546_, _01545_, _01493_);
  nor (_01547_, _01546_, _01488_);
  or (_01548_, _01547_, _01487_);
  and (_01549_, _01548_, _01464_);
  and (_01550_, _01549_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01551_, _01550_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01552_, _01551_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_01553_, _01552_, _01486_);
  not (_01554_, _01486_);
  nor (_01555_, _01548_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01556_, _01555_, _38782_);
  and (_01557_, _01556_, _38787_);
  and (_01558_, _01557_, _38772_);
  nor (_01559_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01560_, _01559_, _01558_);
  nor (_01561_, _01560_, _01554_);
  nor (_01562_, _01561_, _01553_);
  or (_01563_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_01564_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01565_, _01564_, _01563_);
  and (_01566_, _01565_, _01562_);
  or (_01567_, _01566_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_01568_, _01566_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_01569_, _01568_, _01567_);
  and (_01570_, _38497_, _36455_);
  and (_01571_, _01570_, _38467_);
  or (_01572_, _01571_, _01442_);
  and (_01573_, _01572_, _01455_);
  and (_01574_, _01573_, _01569_);
  or (_01575_, _01574_, _01482_);
  and (_01576_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01577_, _36564_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01578_, _01577_, _42500_);
  nor (_01579_, _01578_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_01580_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_01581_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_01582_, _01581_, _01580_);
  not (_01583_, _01582_);
  nor (_01584_, _01583_, _01579_);
  and (_01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_01586_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01587_, _01586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01588_, _01587_, _01584_);
  and (_01589_, _01588_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01590_, _01589_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01591_, _01590_, _01576_);
  and (_01592_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01593_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_01594_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01595_, _01594_, _01593_);
  or (_01596_, _01595_, _01430_);
  and (_01597_, _01596_, _43100_);
  and (_39283_, _01597_, _01575_);
  and (_01598_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _43100_);
  and (_01599_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_01600_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_01601_, _36509_, _01600_);
  not (_01602_, _01601_);
  not (_01603_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_01604_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_01605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_01607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01609_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_01610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_01611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_01612_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_01613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01614_, _01613_, _01612_);
  and (_01615_, _01614_, _01611_);
  and (_01616_, _01615_, _01610_);
  and (_01617_, _01616_, _01609_);
  and (_01618_, _01617_, _01608_);
  and (_01619_, _01618_, _01607_);
  and (_01620_, _01619_, _01606_);
  and (_01621_, _01620_, _01605_);
  and (_01622_, _01621_, _01604_);
  nor (_01623_, _01622_, _01603_);
  and (_01624_, _01622_, _01603_);
  nor (_01625_, _01624_, _01623_);
  nor (_01626_, _01621_, _01604_);
  nor (_01627_, _01626_, _01622_);
  and (_01628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01631_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01632_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_01634_, _01632_, _01629_);
  and (_01635_, _01634_, _01631_);
  nor (_01637_, _01635_, _01629_);
  nor (_01638_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01640_, _01638_, _01628_);
  not (_01641_, _01640_);
  nor (_01643_, _01641_, _01637_);
  nor (_01644_, _01643_, _01628_);
  not (_01646_, _01644_);
  and (_01647_, _01646_, _01619_);
  and (_01649_, _01647_, _01606_);
  and (_01650_, _01649_, _01605_);
  not (_01652_, _01650_);
  nor (_01653_, _01652_, _01627_);
  and (_01655_, _01652_, _01627_);
  or (_01656_, _01655_, _01653_);
  not (_01658_, _01656_);
  and (_01659_, _01644_, _01621_);
  and (_01661_, _01644_, _01620_);
  nor (_01662_, _01661_, _01605_);
  nor (_01663_, _01662_, _01659_);
  not (_01664_, _01663_);
  and (_01665_, _01644_, _01619_);
  nor (_01666_, _01665_, _01606_);
  nor (_01667_, _01666_, _01661_);
  not (_01668_, _01667_);
  and (_01669_, _01644_, _01617_);
  and (_01670_, _01669_, _01608_);
  nor (_01671_, _01670_, _01607_);
  nor (_01672_, _01671_, _01665_);
  not (_01673_, _01672_);
  nor (_01674_, _01669_, _01608_);
  nor (_01675_, _01674_, _01670_);
  not (_01676_, _01675_);
  not (_01677_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_01678_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01679_, _01644_, _01616_);
  and (_01680_, _01679_, _01678_);
  nor (_01681_, _01680_, _01677_);
  nor (_01682_, _01681_, _01669_);
  not (_01683_, _01682_);
  and (_01684_, _01644_, _01614_);
  and (_01685_, _01684_, _01611_);
  nor (_01686_, _01685_, _01610_);
  nor (_01687_, _01686_, _01679_);
  not (_01688_, _01687_);
  nor (_01689_, _01684_, _01611_);
  nor (_01690_, _01689_, _01685_);
  not (_01691_, _01690_);
  and (_01692_, _01644_, _01613_);
  nor (_01693_, _01692_, _01612_);
  nor (_01694_, _01693_, _01684_);
  not (_01695_, _01694_);
  not (_01696_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01697_, _01644_, _01696_);
  nor (_01698_, _01644_, _01696_);
  nor (_01699_, _01698_, _01697_);
  not (_01700_, _01699_);
  nor (_01701_, _00695_, _00653_);
  not (_01702_, _00690_);
  and (_01703_, _01702_, _00686_);
  and (_01704_, _01703_, _01701_);
  nand (_01705_, _00646_, _00641_);
  and (_01706_, _00656_, _00641_);
  and (_01707_, _00674_, _00642_);
  and (_01708_, _01707_, _00634_);
  nor (_01709_, _01708_, _01706_);
  and (_01710_, _01709_, _01705_);
  and (_01711_, _00661_, _00626_);
  and (_01712_, _00642_, _00626_);
  or (_01713_, _01712_, _01711_);
  and (_01714_, _01713_, _00623_);
  not (_01715_, _00641_);
  nor (_01716_, _00692_, _00650_);
  nor (_01717_, _01716_, _01715_);
  nor (_01718_, _01717_, _01714_);
  and (_01719_, _01718_, _01710_);
  not (_01720_, _00623_);
  and (_01721_, _00643_, _00649_);
  nor (_01722_, _01721_, _00656_);
  or (_01723_, _01722_, _01720_);
  nand (_01724_, _00641_, _00620_);
  and (_01725_, _01724_, _01723_);
  and (_01726_, _00643_, _00655_);
  nor (_01727_, _01726_, _00683_);
  nor (_01728_, _01727_, _01715_);
  nor (_01729_, _01728_, _00647_);
  and (_01730_, _01729_, _01725_);
  and (_01731_, _01730_, _01719_);
  and (_01732_, _01731_, _01704_);
  not (_01733_, _00665_);
  and (_01734_, _00656_, _00632_);
  nor (_01735_, _01734_, _00645_);
  and (_01736_, _01735_, _01733_);
  not (_01737_, _01707_);
  nor (_01738_, _00640_, _00623_);
  nor (_01739_, _01738_, _01737_);
  and (_01740_, _00643_, _37164_);
  nor (_01741_, _01740_, _01711_);
  nor (_01742_, _01741_, _00660_);
  nor (_01743_, _01742_, _01739_);
  and (_01744_, _01743_, _01736_);
  nand (_01745_, _00633_, _00620_);
  and (_01746_, _00674_, _00618_);
  nor (_01747_, _00639_, _38410_);
  and (_01748_, _01747_, _00687_);
  and (_01749_, _01748_, _01746_);
  and (_01750_, _00650_, _00623_);
  and (_01751_, _00681_, _00632_);
  or (_01752_, _01751_, _01750_);
  nor (_01753_, _01752_, _01749_);
  and (_01754_, _01753_, _01745_);
  and (_01755_, _00643_, _00661_);
  nand (_01756_, _01755_, _00641_);
  and (_01757_, _00652_, _01712_);
  and (_01758_, _00692_, _00632_);
  nor (_01759_, _01758_, _01757_);
  and (_01760_, _01759_, _01756_);
  and (_01761_, _01721_, _00641_);
  and (_01762_, _00656_, _00652_);
  nor (_01763_, _01762_, _01761_);
  nor (_01764_, _01747_, _00628_);
  not (_01765_, _01764_);
  and (_01766_, _01765_, _00656_);
  and (_01767_, _00683_, _00634_);
  nor (_01768_, _01767_, _01766_);
  and (_01769_, _01768_, _01763_);
  and (_01770_, _01769_, _01760_);
  and (_01771_, _01770_, _01754_);
  and (_01772_, _01771_, _01744_);
  and (_01773_, _01772_, _01732_);
  and (_01774_, _00650_, _00628_);
  and (_01775_, _01747_, _00626_);
  and (_01776_, _01775_, _00667_);
  nor (_01777_, _00692_, _01711_);
  nor (_01778_, _01777_, _38432_);
  or (_01779_, _01778_, _01776_);
  nor (_01780_, _01779_, _01774_);
  nor (_01781_, _00675_, _01712_);
  not (_01782_, _01781_);
  and (_01783_, _01782_, _00640_);
  and (_01784_, _00683_, _00632_);
  nor (_01785_, _01784_, _00623_);
  not (_01786_, _00683_);
  nor (_01787_, _00692_, _00644_);
  and (_01788_, _01787_, _01786_);
  nor (_01789_, _01788_, _01785_);
  and (_01790_, _00675_, _00622_);
  or (_01791_, _01790_, _01789_);
  nor (_01792_, _01791_, _01783_);
  and (_01793_, _01792_, _01780_);
  and (_01794_, _01793_, _01773_);
  nor (_01795_, _01634_, _01631_);
  nor (_01796_, _01795_, _01635_);
  not (_01797_, _01796_);
  nor (_01798_, _01797_, _01794_);
  and (_01799_, _00675_, _00634_);
  nor (_01800_, _01767_, _01799_);
  nor (_01801_, _00682_, _00647_);
  nor (_01802_, _01717_, _01757_);
  and (_01803_, _01802_, _01801_);
  and (_01804_, _01803_, _01800_);
  not (_01805_, _01766_);
  and (_01806_, _01709_, _01736_);
  and (_01807_, _01806_, _01805_);
  and (_01808_, _01807_, _01804_);
  not (_01809_, _01808_);
  nor (_01810_, _01809_, _01794_);
  not (_01811_, _01810_);
  nor (_01812_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01813_, _01812_, _01631_);
  and (_01814_, _01813_, _01811_);
  and (_01815_, _01797_, _01794_);
  nor (_01816_, _01815_, _01798_);
  and (_01817_, _01816_, _01814_);
  nor (_01818_, _01817_, _01798_);
  not (_01819_, _01818_);
  and (_01820_, _01641_, _01637_);
  nor (_01821_, _01820_, _01643_);
  and (_01822_, _01821_, _01819_);
  and (_01823_, _01822_, _01700_);
  not (_01824_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_01825_, _01697_, _01824_);
  or (_01826_, _01825_, _01692_);
  and (_01827_, _01826_, _01823_);
  and (_01828_, _01827_, _01695_);
  and (_01829_, _01828_, _01691_);
  and (_01830_, _01829_, _01688_);
  nor (_01831_, _01679_, _01678_);
  or (_01832_, _01831_, _01680_);
  and (_01833_, _01832_, _01830_);
  and (_01834_, _01833_, _01683_);
  and (_01835_, _01834_, _01676_);
  and (_01836_, _01835_, _01673_);
  and (_01837_, _01836_, _01668_);
  and (_01838_, _01837_, _01664_);
  and (_01839_, _01838_, _01658_);
  nor (_01840_, _01839_, _01653_);
  not (_01841_, _01840_);
  nor (_01842_, _01841_, _01625_);
  and (_01843_, _01841_, _01625_);
  or (_01844_, _01843_, _01842_);
  or (_01845_, _01844_, _01602_);
  or (_01846_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_01847_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_01848_, _01847_, _01846_);
  and (_01849_, _01848_, _01845_);
  or (_39285_, _01849_, _01599_);
  nor (_01850_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_39286_, _01850_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_39287_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _43100_);
  not (_01851_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor (_01852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_01853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01854_, _01853_, _01852_);
  not (_01855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_01856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_01857_, _01856_, _01855_);
  and (_01858_, _01857_, _01854_);
  and (_01859_, _01858_, _01851_);
  and (_01860_, \oc8051_top_1.oc8051_rom1.ea_int , _36477_);
  nand (_01861_, _01860_, _36509_);
  nand (_01862_, _01861_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_01863_, _01862_, _01859_);
  and (_39288_, _01863_, _43100_);
  and (_01864_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_01865_, _01864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_39290_, _01865_, _43100_);
  nor (_01866_, _01579_, _42500_);
  nor (_01867_, _01794_, _36760_);
  nor (_01868_, _01810_, _36629_);
  and (_01869_, _01794_, _36760_);
  nor (_01870_, _01869_, _01867_);
  and (_01871_, _01870_, _01868_);
  nor (_01872_, _01871_, _01867_);
  nor (_01873_, _01872_, _42500_);
  and (_01874_, _01873_, _36553_);
  nor (_01875_, _01873_, _36553_);
  nor (_01876_, _01875_, _01874_);
  nor (_01877_, _01876_, _01866_);
  and (_01878_, _36770_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_01879_, _01878_, _01866_);
  nor (_01880_, _01879_, _01808_);
  or (_01881_, _01880_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01882_, _01881_, _01877_);
  and (_39291_, _01882_, _43100_);
  nor (_01883_, _36825_, _38149_);
  and (_01884_, _37612_, _37382_);
  and (_01885_, _01884_, _01883_);
  nand (_01886_, _01323_, _38406_);
  nor (_01887_, _01886_, _37907_);
  not (_01888_, _38428_);
  and (_01889_, _37121_, _01888_);
  and (_01890_, _01889_, _01887_);
  and (_39294_, _01890_, _01885_);
  nor (_01891_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_01892_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_01893_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_39297_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _43100_);
  and (_01894_, _39297_, _01893_);
  or (_39295_, _01894_, _01892_);
  not (_01895_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01896_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01897_, _01896_, _01895_);
  and (_01898_, _01896_, _01895_);
  nor (_01899_, _01898_, _01897_);
  not (_01900_, _01899_);
  and (_01901_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01902_, _01901_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01903_, _01901_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01904_, _01903_, _01902_);
  or (_01905_, _01904_, _01896_);
  and (_01906_, _01905_, _01900_);
  nor (_01907_, _01897_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01908_, _01897_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_01909_, _01908_, _01907_);
  or (_01910_, _01902_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_39299_, _01910_, _43100_);
  and (_01911_, _39299_, _01909_);
  and (_39298_, _01911_, _01906_);
  not (_01912_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_01913_, _01579_, _01912_);
  and (_01914_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_01915_, _01913_);
  and (_01916_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_01917_, _01916_, _01914_);
  and (_39300_, _01917_, _43100_);
  and (_01918_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01919_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_01920_, _01919_, _01918_);
  and (_39301_, _01920_, _43100_);
  and (_01921_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_01922_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_01923_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _01922_);
  and (_01924_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_01925_, _01924_, _01921_);
  and (_39302_, _01925_, _43100_);
  and (_01926_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_01927_, _01926_, _01923_);
  and (_39303_, _01927_, _43100_);
  or (_01928_, _01922_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_39305_, _01928_, _43100_);
  not (_01929_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_01930_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01931_, _01930_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_01932_, _01922_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_01933_, _01932_, _43100_);
  and (_39306_, _01933_, _01931_);
  or (_01934_, _01922_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_39307_, _01934_, _43100_);
  nor (_01935_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_01936_, _01935_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_01937_, _01936_, _43100_);
  and (_01938_, _39297_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_39308_, _01938_, _01937_);
  and (_01939_, _01912_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_01940_, _01939_, _01936_);
  and (_39309_, _01940_, _43100_);
  nand (_01941_, _01936_, _38845_);
  or (_01942_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_01943_, _01942_, _43100_);
  and (_39310_, _01943_, _01941_);
  nand (_01944_, _38477_, _43100_);
  nor (_39311_, _01944_, _38614_);
  or (_01945_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_01946_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_01947_, _01317_, _01946_);
  and (_01948_, _01947_, _43100_);
  and (_39347_, _01948_, _01945_);
  or (_01949_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_01950_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_01951_, _01317_, _01950_);
  and (_01952_, _01951_, _43100_);
  and (_39348_, _01952_, _01949_);
  or (_01953_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_01954_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_01955_, _01317_, _01954_);
  and (_01956_, _01955_, _43100_);
  and (_39349_, _01956_, _01953_);
  or (_01957_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_01958_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_01959_, _01317_, _01958_);
  and (_01960_, _01959_, _43100_);
  and (_39350_, _01960_, _01957_);
  or (_01961_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_01962_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_01963_, _01317_, _01962_);
  and (_01964_, _01963_, _43100_);
  and (_39351_, _01964_, _01961_);
  or (_01965_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_01966_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_01967_, _01317_, _01966_);
  and (_01968_, _01967_, _43100_);
  and (_39353_, _01968_, _01965_);
  or (_01969_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_01970_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01971_, _01970_, _43100_);
  and (_39354_, _01971_, _01969_);
  or (_01972_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_01973_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_01974_, _01317_, _01973_);
  and (_01975_, _01974_, _43100_);
  and (_39355_, _01975_, _01972_);
  or (_01976_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_01977_, _01317_, _38776_);
  and (_01978_, _01977_, _43100_);
  and (_39356_, _01978_, _01976_);
  or (_01979_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_01980_, _01317_, _38782_);
  and (_01981_, _01980_, _43100_);
  and (_39357_, _01981_, _01979_);
  or (_01982_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_01983_, _01317_, _38787_);
  and (_01984_, _01983_, _43100_);
  and (_39358_, _01984_, _01982_);
  or (_01985_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_01986_, _01317_, _38772_);
  and (_01987_, _01986_, _43100_);
  and (_39359_, _01987_, _01985_);
  or (_01988_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_01989_, _01317_, _38793_);
  and (_01990_, _01989_, _43100_);
  and (_39360_, _01990_, _01988_);
  or (_01991_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_01992_, _01317_, _38768_);
  and (_01993_, _01992_, _43100_);
  and (_39361_, _01993_, _01991_);
  or (_01994_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_01995_, _01317_, _38764_);
  and (_01996_, _01995_, _43100_);
  and (_39362_, _01996_, _01994_);
  and (_01997_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_01998_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_01999_, _01998_, _01997_);
  and (_39367_, _01999_, _43100_);
  and (_02000_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_02001_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_02002_, _02001_, _02000_);
  and (_39368_, _02002_, _43100_);
  and (_02003_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_02004_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_02005_, _02004_, _02003_);
  and (_39369_, _02005_, _43100_);
  and (_02006_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_02007_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_02008_, _02007_, _02006_);
  and (_39370_, _02008_, _43100_);
  and (_02009_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_02010_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or (_02011_, _02010_, _02009_);
  and (_39371_, _02011_, _43100_);
  and (_02012_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_02013_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or (_02014_, _02013_, _02012_);
  and (_39372_, _02014_, _43100_);
  and (_02015_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_02016_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or (_02017_, _02016_, _02015_);
  and (_39373_, _02017_, _43100_);
  and (_02018_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_02019_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or (_02020_, _02019_, _02018_);
  and (_39374_, _02020_, _43100_);
  and (_02021_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_02022_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or (_02023_, _02022_, _02021_);
  and (_39375_, _02023_, _43100_);
  and (_02024_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_02025_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or (_02026_, _02025_, _02024_);
  and (_39376_, _02026_, _43100_);
  and (_02027_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_02028_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or (_02029_, _02028_, _02027_);
  and (_39378_, _02029_, _43100_);
  and (_02030_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_02031_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or (_02032_, _02031_, _02030_);
  and (_39379_, _02032_, _43100_);
  and (_02033_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_02034_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or (_02035_, _02034_, _02033_);
  and (_39380_, _02035_, _43100_);
  and (_02036_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_02037_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or (_02038_, _02037_, _02036_);
  and (_39381_, _02038_, _43100_);
  and (_02039_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_02040_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or (_02041_, _02040_, _02039_);
  and (_39382_, _02041_, _43100_);
  and (_39558_, _38006_, _43100_);
  and (_39559_, _38270_, _43100_);
  and (_39560_, _38414_, _43100_);
  nor (_39561_, _42476_, rst);
  and (_02042_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02043_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_02044_, _02043_, _02042_);
  and (_39562_, _02044_, _43100_);
  and (_02045_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_02046_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_02047_, _02046_, _02045_);
  and (_39563_, _02047_, _43100_);
  and (_02048_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02049_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_02050_, _02049_, _02048_);
  and (_39564_, _02050_, _43100_);
  and (_02051_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02052_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_02053_, _02052_, _02051_);
  and (_39565_, _02053_, _43100_);
  and (_02054_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02055_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_02056_, _02055_, _02054_);
  and (_39567_, _02056_, _43100_);
  and (_02057_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02058_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_02059_, _02058_, _02057_);
  and (_39568_, _02059_, _43100_);
  and (_02060_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02061_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_02062_, _02061_, _02060_);
  and (_39569_, _02062_, _43100_);
  and (_02063_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02064_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_02065_, _02064_, _02063_);
  and (_39570_, _02065_, _43100_);
  and (_02066_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_02067_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_02068_, _02067_, _02066_);
  and (_39571_, _02068_, _43100_);
  and (_02069_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_02070_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_02071_, _02070_, _02069_);
  and (_39572_, _02071_, _43100_);
  and (_02072_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_02073_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_02074_, _02073_, _02072_);
  and (_39573_, _02074_, _43100_);
  and (_02075_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_02076_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_02077_, _02076_, _02075_);
  and (_39574_, _02077_, _43100_);
  and (_02078_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_02079_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_02080_, _02079_, _02078_);
  and (_39575_, _02080_, _43100_);
  and (_02081_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_02082_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_02083_, _02082_, _02081_);
  and (_39576_, _02083_, _43100_);
  and (_02084_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_02085_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_02086_, _02085_, _02084_);
  and (_39578_, _02086_, _43100_);
  and (_02087_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_02088_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_02089_, _02088_, _02087_);
  and (_39579_, _02089_, _43100_);
  and (_02090_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_02091_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_02092_, _02091_, _02090_);
  and (_39580_, _02092_, _43100_);
  and (_02093_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_02094_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_02095_, _02094_, _02093_);
  and (_39581_, _02095_, _43100_);
  and (_02096_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_02097_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_02098_, _02097_, _02096_);
  and (_39582_, _02098_, _43100_);
  and (_02099_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_02100_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_02101_, _02100_, _02099_);
  and (_39583_, _02101_, _43100_);
  and (_02102_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_02103_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_02104_, _02103_, _02102_);
  and (_39584_, _02104_, _43100_);
  and (_02105_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_02106_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_02107_, _02106_, _02105_);
  and (_39585_, _02107_, _43100_);
  and (_02108_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_02109_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_02110_, _02109_, _02108_);
  and (_39586_, _02110_, _43100_);
  and (_02111_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_02113_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_02115_, _02113_, _02111_);
  and (_39587_, _02115_, _43100_);
  and (_02118_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_02120_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_02122_, _02120_, _02118_);
  and (_39589_, _02122_, _43100_);
  and (_02125_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_02127_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_02129_, _02127_, _02125_);
  and (_39590_, _02129_, _43100_);
  and (_02132_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_02134_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_02136_, _02134_, _02132_);
  and (_39591_, _02136_, _43100_);
  and (_02139_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_02141_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_02143_, _02141_, _02139_);
  and (_39592_, _02143_, _43100_);
  and (_02146_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_02148_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_02150_, _02148_, _02146_);
  and (_39593_, _02150_, _43100_);
  and (_02153_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_02155_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_02157_, _02155_, _02153_);
  and (_39594_, _02157_, _43100_);
  and (_02160_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_02162_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_02164_, _02162_, _02160_);
  and (_39595_, _02164_, _43100_);
  nor (_39596_, _42697_, rst);
  nor (_39598_, _42591_, rst);
  nor (_39599_, _42815_, rst);
  nor (_39600_, _42661_, rst);
  nor (_39601_, _42575_, rst);
  and (_39602_, _42762_, _43100_);
  nor (_39604_, _42720_, rst);
  and (_39620_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _43100_);
  and (_39621_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _43100_);
  and (_39622_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _43100_);
  and (_39623_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _43100_);
  and (_39624_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _43100_);
  and (_39626_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _43100_);
  and (_39627_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _43100_);
  or (_02170_, _01477_, _01435_);
  and (_02171_, _02170_, _31809_);
  or (_02172_, _01526_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_02173_, _01527_);
  nor (_02174_, _01450_, _01442_);
  not (_02175_, _02174_);
  and (_02176_, _02175_, _01455_);
  and (_02177_, _02176_, _02173_);
  and (_02178_, _02177_, _02172_);
  and (_02179_, _01456_, _42683_);
  and (_02180_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_02181_, _02180_, _02179_);
  and (_02182_, _01447_, _01524_);
  or (_02183_, _02182_, _02181_);
  nor (_02184_, _02183_, _02178_);
  nand (_02185_, _02184_, _01430_);
  or (_02186_, _02185_, _02171_);
  or (_02187_, _01430_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_02188_, _02187_, _43100_);
  and (_39628_, _02188_, _02186_);
  and (_02189_, _02170_, _32506_);
  or (_02190_, _01529_, _01527_);
  not (_02191_, _01530_);
  and (_02192_, _02176_, _02191_);
  and (_02193_, _02192_, _02190_);
  and (_02194_, _01456_, _42612_);
  and (_02195_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_02196_, _02195_, _02194_);
  and (_02197_, _01447_, _01519_);
  or (_02198_, _02197_, _02196_);
  nor (_02199_, _02198_, _02193_);
  nand (_02200_, _02199_, _01430_);
  or (_02201_, _02200_, _02189_);
  or (_02202_, _01430_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_02203_, _02202_, _43100_);
  and (_39629_, _02203_, _02201_);
  and (_02204_, _02170_, _33213_);
  or (_02205_, _01534_, _01532_);
  not (_02206_, _01535_);
  and (_02207_, _02176_, _02206_);
  and (_02208_, _02207_, _02205_);
  and (_02209_, _01456_, _42804_);
  and (_02210_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_02211_, _02210_, _02209_);
  and (_02212_, _01447_, _01514_);
  or (_02213_, _02212_, _02211_);
  nor (_02214_, _02213_, _02208_);
  nand (_02215_, _02214_, _01430_);
  or (_02216_, _02215_, _02204_);
  not (_02217_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02218_, _01579_, _02217_);
  and (_02219_, _01579_, _02217_);
  nor (_02220_, _02219_, _02218_);
  or (_02221_, _02220_, _01430_);
  and (_02222_, _02221_, _43100_);
  and (_39630_, _02222_, _02216_);
  and (_02223_, _02170_, _33964_);
  or (_02224_, _01512_, _01511_);
  or (_02225_, _02224_, _01536_);
  nand (_02226_, _02224_, _01536_);
  and (_02227_, _02226_, _02176_);
  and (_02228_, _02227_, _02225_);
  and (_02229_, _01456_, _42647_);
  and (_02230_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_02231_, _02230_, _02229_);
  and (_02232_, _01447_, _01508_);
  or (_02233_, _02232_, _02231_);
  nor (_02234_, _02233_, _02228_);
  nand (_02235_, _02234_, _01430_);
  or (_02236_, _02235_, _02223_);
  and (_02237_, _02218_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02238_, _02218_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02239_, _02238_, _02237_);
  or (_02240_, _02239_, _01430_);
  and (_02241_, _02240_, _43100_);
  and (_39631_, _02241_, _02236_);
  and (_02242_, _02170_, _34704_);
  or (_02243_, _01540_, _01538_);
  and (_02244_, _02176_, _01541_);
  and (_02245_, _02244_, _02243_);
  and (_02246_, _01456_, _42552_);
  and (_02247_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_02248_, _02247_, _02246_);
  and (_02249_, _01447_, _01503_);
  or (_02250_, _02249_, _02248_);
  nor (_02251_, _02250_, _02245_);
  nand (_02252_, _02251_, _01430_);
  or (_02253_, _02252_, _02242_);
  and (_02254_, _02237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02255_, _02237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02256_, _02255_, _02254_);
  or (_02257_, _02256_, _01430_);
  and (_02258_, _02257_, _43100_);
  and (_39632_, _02258_, _02253_);
  and (_02259_, _02170_, _35531_);
  and (_02260_, _01456_, _42778_);
  and (_02261_, _01447_, _01497_);
  and (_02262_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_02263_, _02262_, _02261_);
  or (_02264_, _02263_, _02260_);
  or (_02265_, _01501_, _01500_);
  or (_02266_, _02265_, _01542_);
  nand (_02267_, _02265_, _01542_);
  and (_02268_, _02267_, _02176_);
  and (_02269_, _02268_, _02266_);
  nor (_02270_, _02269_, _02264_);
  nand (_02271_, _02270_, _01430_);
  or (_02272_, _02271_, _02259_);
  nor (_02273_, _02254_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02274_, _02273_, _01584_);
  or (_02275_, _02274_, _01430_);
  and (_02276_, _02275_, _43100_);
  and (_39633_, _02276_, _02272_);
  nor (_02277_, _01584_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02278_, _01584_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_02279_, _02278_, _02277_);
  or (_02280_, _02279_, _01430_);
  and (_02281_, _02280_, _43100_);
  and (_02282_, _02170_, _36249_);
  or (_02283_, _01544_, _01495_);
  not (_02284_, _01545_);
  and (_02285_, _02176_, _02284_);
  and (_02286_, _02285_, _02283_);
  and (_02287_, _01456_, _42740_);
  and (_02288_, _01447_, _01490_);
  and (_02289_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_02290_, _02289_, _02288_);
  or (_02291_, _02290_, _02287_);
  nor (_02292_, _02291_, _02286_);
  nand (_02293_, _02292_, _01430_);
  or (_02294_, _02293_, _02282_);
  and (_39634_, _02294_, _02281_);
  and (_02295_, _02170_, _30585_);
  or (_02296_, _01487_, _01488_);
  or (_02297_, _02296_, _01546_);
  nand (_02298_, _02296_, _01546_);
  and (_02299_, _02298_, _02176_);
  and (_02300_, _02299_, _02297_);
  and (_02301_, _01456_, _42517_);
  and (_02302_, _01447_, _01484_);
  and (_02303_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_02304_, _02303_, _02302_);
  nor (_02305_, _02304_, _02301_);
  nand (_02306_, _02305_, _01430_);
  or (_02307_, _02306_, _02300_);
  or (_02308_, _02307_, _02295_);
  nor (_02309_, _02278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_02310_, _02278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_02311_, _02310_, _02309_);
  or (_02312_, _02311_, _01430_);
  and (_02313_, _02312_, _43100_);
  and (_39635_, _02313_, _02308_);
  nor (_02314_, _01432_, _31808_);
  not (_02315_, _38882_);
  and (_02316_, _01435_, _02315_);
  and (_02317_, _01548_, _38776_);
  nor (_02318_, _01548_, _38776_);
  nor (_02319_, _02318_, _02317_);
  nor (_02320_, _02319_, _01486_);
  and (_02321_, _02319_, _01486_);
  or (_02322_, _02321_, _02320_);
  and (_02323_, _02322_, _02176_);
  nand (_02324_, _01447_, _42683_);
  and (_02325_, _01456_, _00618_);
  and (_02326_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_02327_, _02326_, _02325_);
  and (_02328_, _02327_, _02324_);
  nand (_02329_, _02328_, _01430_);
  or (_02330_, _02329_, _02323_);
  or (_02331_, _02330_, _02316_);
  or (_02332_, _02331_, _02314_);
  or (_02333_, _02310_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_02334_, _01586_, _01584_);
  and (_02335_, _02334_, _02333_);
  or (_02336_, _02335_, _01430_);
  and (_02337_, _02336_, _43100_);
  and (_39636_, _02337_, _02332_);
  nor (_02338_, _01432_, _32495_);
  and (_02339_, _01548_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02340_, _02339_, _01554_);
  and (_02341_, _01555_, _01486_);
  nor (_02342_, _02341_, _02340_);
  nand (_02343_, _02342_, _38782_);
  or (_02344_, _02342_, _38782_);
  and (_02345_, _02344_, _02176_);
  and (_02346_, _02345_, _02343_);
  not (_02347_, _38916_);
  and (_02348_, _01435_, _02347_);
  and (_02349_, _01456_, _00673_);
  and (_02350_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_02351_, _01447_, _42612_);
  or (_02352_, _02351_, _02350_);
  or (_02353_, _02352_, _02349_);
  nor (_02354_, _02353_, _02348_);
  nand (_02355_, _02354_, _01430_);
  or (_02356_, _02355_, _02346_);
  or (_02357_, _02356_, _02338_);
  nand (_02358_, _02334_, _01677_);
  or (_02360_, _02334_, _01677_);
  and (_02361_, _02360_, _02358_);
  or (_02362_, _02361_, _01430_);
  and (_02363_, _02362_, _43100_);
  and (_39637_, _02363_, _02357_);
  nor (_02364_, _01432_, _33202_);
  and (_02365_, _01556_, _01486_);
  and (_02366_, _02340_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_02367_, _02366_, _02365_);
  nor (_02368_, _02367_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_02369_, _02367_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_02370_, _02369_, _02368_);
  and (_02371_, _02370_, _02176_);
  not (_02372_, _38947_);
  and (_02373_, _01435_, _02372_);
  and (_02374_, _01456_, _00625_);
  and (_02375_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_02376_, _01447_, _42804_);
  or (_02377_, _02376_, _02375_);
  or (_02378_, _02377_, _02374_);
  nor (_02379_, _02378_, _02373_);
  nand (_02380_, _02379_, _01430_);
  or (_02381_, _02380_, _02371_);
  or (_02382_, _02381_, _02364_);
  nor (_02383_, _01588_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_02384_, _02383_, _01589_);
  or (_02385_, _02384_, _01430_);
  and (_02386_, _02385_, _43100_);
  and (_39638_, _02386_, _02382_);
  nor (_02387_, _01432_, _33953_);
  and (_02388_, _01549_, _01554_);
  and (_02389_, _01557_, _01486_);
  nor (_02390_, _02389_, _02388_);
  nand (_02391_, _02390_, _38772_);
  or (_02392_, _02390_, _38772_);
  and (_02393_, _02392_, _02176_);
  and (_02394_, _02393_, _02391_);
  not (_02395_, _38976_);
  and (_02396_, _01435_, _02395_);
  and (_02397_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02398_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_02399_, _02398_, _01466_);
  and (_02400_, _02399_, _01456_);
  and (_02401_, _01447_, _42647_);
  or (_02402_, _02401_, _02400_);
  or (_02403_, _02402_, _02397_);
  nor (_02404_, _02403_, _02396_);
  nand (_02405_, _02404_, _01430_);
  or (_02406_, _02405_, _02394_);
  or (_02407_, _02406_, _02387_);
  nor (_02408_, _01589_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02409_, _02408_, _01590_);
  or (_02410_, _02409_, _01430_);
  and (_02411_, _02410_, _43100_);
  and (_39639_, _02411_, _02407_);
  nor (_02412_, _01432_, _34693_);
  and (_02413_, _01550_, _01554_);
  and (_02414_, _01558_, _01486_);
  nor (_02415_, _02414_, _02413_);
  nand (_02416_, _02415_, _38793_);
  or (_02417_, _02415_, _38793_);
  and (_02418_, _02417_, _02176_);
  and (_02419_, _02418_, _02416_);
  not (_02420_, _39007_);
  nand (_02421_, _01435_, _02420_);
  nor (_02422_, _01466_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_02423_, _02422_, _01467_);
  and (_02424_, _02423_, _01456_);
  and (_02425_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_02426_, _01447_, _42552_);
  or (_02427_, _02426_, _02425_);
  nor (_02428_, _02427_, _02424_);
  and (_02429_, _02428_, _02421_);
  nand (_02430_, _02429_, _01430_);
  or (_02431_, _02430_, _02419_);
  or (_02432_, _02431_, _02412_);
  nor (_02433_, _01590_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_02434_, _01590_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_02435_, _02434_, _02433_);
  or (_02436_, _02435_, _01430_);
  and (_02437_, _02436_, _43100_);
  and (_39640_, _02437_, _02432_);
  nor (_02438_, _01432_, _35520_);
  and (_02439_, _01551_, _01554_);
  and (_02440_, _02414_, _38793_);
  nor (_02441_, _02440_, _02439_);
  nand (_02442_, _02441_, _38768_);
  or (_02443_, _02441_, _38768_);
  and (_02444_, _02443_, _02176_);
  and (_02445_, _02444_, _02442_);
  not (_02446_, _39041_);
  nand (_02447_, _01435_, _02446_);
  nor (_02448_, _01467_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_02449_, _02448_, _01468_);
  and (_02450_, _02449_, _01456_);
  and (_02451_, _01447_, _42778_);
  or (_02452_, _02451_, _02450_);
  and (_02453_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_02454_, _02453_, _02452_);
  and (_02455_, _02454_, _02447_);
  nand (_02456_, _02455_, _01430_);
  or (_02457_, _02456_, _02445_);
  or (_02458_, _02457_, _02438_);
  or (_02459_, _02434_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_02460_, _02434_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_02461_, _02460_, _02459_);
  or (_02462_, _02461_, _01430_);
  and (_02463_, _02462_, _43100_);
  and (_39641_, _02463_, _02458_);
  nor (_02464_, _01432_, _36239_);
  nor (_02465_, _01562_, _38764_);
  and (_02466_, _01562_, _38764_);
  or (_02467_, _02466_, _02465_);
  and (_02468_, _02467_, _02176_);
  not (_02469_, _39071_);
  nand (_02470_, _01435_, _02469_);
  nor (_02471_, _01468_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_02472_, _02471_, _01469_);
  and (_02473_, _02472_, _01456_);
  and (_02474_, _01447_, _42740_);
  or (_02475_, _02474_, _02473_);
  and (_02476_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_02477_, _02476_, _02475_);
  and (_02478_, _02477_, _02470_);
  nand (_02479_, _02478_, _01430_);
  or (_02480_, _02479_, _02468_);
  or (_02481_, _02480_, _02464_);
  nor (_02482_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_02483_, _02482_, _01592_);
  or (_02484_, _02483_, _01430_);
  and (_02485_, _02484_, _43100_);
  and (_39642_, _02485_, _02481_);
  and (_02486_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_02487_, _01813_, _01811_);
  nor (_02488_, _02487_, _01814_);
  or (_02489_, _02488_, _01602_);
  or (_02490_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_02491_, _02490_, _01847_);
  and (_02492_, _02491_, _02489_);
  or (_39643_, _02492_, _02486_);
  nor (_02493_, _01816_, _01814_);
  nor (_02494_, _02493_, _01817_);
  or (_02495_, _02494_, _01602_);
  or (_02496_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_02497_, _02496_, _01847_);
  and (_02498_, _02497_, _02495_);
  and (_02499_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39644_, _02499_, _02498_);
  or (_02500_, _01821_, _01819_);
  nor (_02501_, _01602_, _01822_);
  and (_02502_, _02501_, _02500_);
  nor (_02503_, _01601_, _01954_);
  or (_02504_, _02503_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02505_, _02504_, _02502_);
  or (_02506_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _36477_);
  and (_02507_, _02506_, _43100_);
  and (_39645_, _02507_, _02505_);
  and (_02508_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02509_, _01822_, _01700_);
  nor (_02510_, _02509_, _01823_);
  or (_02511_, _02510_, _01602_);
  or (_02512_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_02513_, _02512_, _01847_);
  and (_02514_, _02513_, _02511_);
  or (_39647_, _02514_, _02508_);
  and (_02515_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02516_, _01826_, _01823_);
  nor (_02517_, _02516_, _01827_);
  or (_02518_, _02517_, _01602_);
  or (_02519_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_02520_, _02519_, _01847_);
  and (_02521_, _02520_, _02518_);
  or (_39648_, _02521_, _02515_);
  and (_02522_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02523_, _01827_, _01695_);
  nor (_02524_, _02523_, _01828_);
  or (_02525_, _02524_, _01602_);
  or (_02526_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_02527_, _02526_, _01847_);
  and (_02528_, _02527_, _02525_);
  or (_39649_, _02528_, _02522_);
  nor (_02529_, _01828_, _01691_);
  nor (_02530_, _02529_, _01829_);
  or (_02531_, _02530_, _01602_);
  or (_02532_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_02533_, _02532_, _01847_);
  and (_02534_, _02533_, _02531_);
  and (_02535_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39650_, _02535_, _02534_);
  nor (_02536_, _01829_, _01688_);
  nor (_02537_, _02536_, _01830_);
  or (_02538_, _02537_, _01602_);
  or (_02539_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_02540_, _02539_, _01847_);
  and (_02541_, _02540_, _02538_);
  and (_02542_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_39651_, _02542_, _02541_);
  and (_02543_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_02544_, _01832_, _01830_);
  nor (_02545_, _02544_, _01833_);
  or (_02547_, _02545_, _01602_);
  or (_02548_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02549_, _02548_, _01847_);
  and (_02550_, _02549_, _02547_);
  or (_39652_, _02550_, _02543_);
  nor (_02551_, _01833_, _01683_);
  nor (_02552_, _02551_, _01834_);
  or (_02553_, _02552_, _01602_);
  or (_02554_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_02555_, _02554_, _01847_);
  and (_02556_, _02555_, _02553_);
  and (_02557_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_39653_, _02557_, _02556_);
  or (_02558_, _01834_, _01676_);
  nor (_02559_, _01602_, _01835_);
  and (_02560_, _02559_, _02558_);
  nor (_02561_, _01601_, _38787_);
  or (_02562_, _02561_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02563_, _02562_, _02560_);
  or (_02564_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _36477_);
  and (_02565_, _02564_, _43100_);
  and (_39654_, _02565_, _02563_);
  nor (_02566_, _01835_, _01673_);
  nor (_02568_, _02566_, _01836_);
  or (_02569_, _02568_, _01602_);
  or (_02570_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_02571_, _02570_, _01847_);
  and (_02572_, _02571_, _02569_);
  and (_02573_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_39655_, _02573_, _02572_);
  and (_02574_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_02575_, _01836_, _01668_);
  nor (_02576_, _02575_, _01837_);
  or (_02577_, _02576_, _01602_);
  or (_02579_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_02580_, _02579_, _01847_);
  and (_02581_, _02580_, _02577_);
  or (_39656_, _02581_, _02574_);
  nor (_02582_, _01837_, _01664_);
  nor (_02583_, _02582_, _01838_);
  or (_02584_, _02583_, _01602_);
  or (_02585_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_02586_, _02585_, _01847_);
  and (_02587_, _02586_, _02584_);
  and (_02588_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_39658_, _02588_, _02587_);
  nor (_02589_, _01838_, _01658_);
  nor (_02590_, _02589_, _01839_);
  or (_02591_, _02590_, _01602_);
  or (_02592_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02593_, _02592_, _01847_);
  and (_02594_, _02593_, _02591_);
  and (_02595_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_39659_, _02595_, _02594_);
  and (_02596_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_02597_, _02596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_39660_, _02597_, _43100_);
  and (_02598_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_02599_, _02598_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_39661_, _02599_, _43100_);
  and (_02600_, _01858_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_02601_, _02600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_39662_, _02601_, _43100_);
  and (_02602_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_02603_, _02602_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39663_, _02603_, _43100_);
  and (_02604_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_02605_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_39664_, _02605_, _43100_);
  and (_02606_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_02607_, _02606_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_39665_, _02607_, _43100_);
  and (_02608_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_02609_, _02608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_39666_, _02609_, _43100_);
  nor (_02610_, _01810_, _42500_);
  nand (_02611_, _02610_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_02612_, _02610_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_02613_, _02612_, _01847_);
  and (_39667_, _02613_, _02611_);
  nor (_02614_, _01870_, _01868_);
  nor (_02615_, _02614_, _01871_);
  or (_02616_, _02615_, _42500_);
  or (_02617_, _36509_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_02618_, _02617_, _01847_);
  and (_39669_, _02618_, _02616_);
  and (_02619_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_02620_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_02621_, _02620_, _39297_);
  or (_39685_, _02621_, _02619_);
  and (_02622_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_02623_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_02624_, _02623_, _39297_);
  or (_39686_, _02624_, _02622_);
  and (_02625_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_02626_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_02627_, _02626_, _39297_);
  or (_39687_, _02627_, _02625_);
  and (_02628_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_02629_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_02630_, _02629_, _39297_);
  or (_39688_, _02630_, _02628_);
  and (_02631_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_02632_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_02633_, _02632_, _39297_);
  or (_39689_, _02633_, _02631_);
  and (_02634_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_02635_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_02636_, _02635_, _39297_);
  or (_39691_, _02636_, _02634_);
  and (_02637_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_02638_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_02639_, _02638_, _39297_);
  or (_39692_, _02639_, _02637_);
  and (_39693_, _01899_, _43100_);
  nor (_39694_, _01909_, rst);
  and (_39695_, _01905_, _43100_);
  and (_02640_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02641_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_02642_, _02641_, _02640_);
  and (_39696_, _02642_, _43100_);
  and (_02643_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_02644_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_02645_, _02644_, _02643_);
  and (_39697_, _02645_, _43100_);
  and (_02646_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02647_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_02648_, _02647_, _02646_);
  and (_39698_, _02648_, _43100_);
  and (_02649_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02650_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_02651_, _02650_, _02649_);
  and (_39699_, _02651_, _43100_);
  and (_02652_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02653_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_02654_, _02653_, _02652_);
  and (_39700_, _02654_, _43100_);
  and (_02655_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02656_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_02657_, _02656_, _02655_);
  and (_39702_, _02657_, _43100_);
  and (_02658_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02659_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_02660_, _02659_, _02658_);
  and (_39703_, _02660_, _43100_);
  and (_02661_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02662_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_02663_, _02662_, _02661_);
  and (_39704_, _02663_, _43100_);
  and (_02664_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_02665_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_02666_, _02665_, _02664_);
  and (_39705_, _02666_, _43100_);
  and (_02667_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_02668_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_02669_, _02668_, _02667_);
  and (_39706_, _02669_, _43100_);
  and (_02670_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_02671_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_02672_, _02671_, _02670_);
  and (_39707_, _02672_, _43100_);
  and (_02673_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_02674_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_02675_, _02674_, _02673_);
  and (_39708_, _02675_, _43100_);
  and (_02676_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_02677_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_02678_, _02677_, _02676_);
  and (_39709_, _02678_, _43100_);
  and (_02679_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_02680_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_02681_, _02680_, _02679_);
  and (_39710_, _02681_, _43100_);
  and (_02682_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_02683_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_02684_, _02683_, _02682_);
  and (_39711_, _02684_, _43100_);
  and (_02685_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_02686_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_02687_, _02686_, _02685_);
  and (_39713_, _02687_, _43100_);
  and (_02688_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_02689_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_02690_, _02689_, _02688_);
  and (_39714_, _02690_, _43100_);
  and (_02691_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_02692_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_02693_, _02692_, _02691_);
  and (_39715_, _02693_, _43100_);
  and (_02694_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_02695_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_02696_, _02695_, _02694_);
  and (_39716_, _02696_, _43100_);
  and (_02697_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_02698_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_02699_, _02698_, _02697_);
  and (_39717_, _02699_, _43100_);
  and (_02700_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_02701_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_02702_, _02701_, _02700_);
  and (_39718_, _02702_, _43100_);
  and (_02704_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_02705_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_02706_, _02705_, _02704_);
  and (_39719_, _02706_, _43100_);
  and (_02707_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_02708_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_02709_, _02708_, _02707_);
  and (_39720_, _02709_, _43100_);
  and (_02710_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_02711_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_02712_, _02711_, _02710_);
  and (_39721_, _02712_, _43100_);
  and (_02713_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_02714_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_02715_, _02714_, _02713_);
  and (_39722_, _02715_, _43100_);
  and (_02716_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_02717_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_02718_, _02717_, _02716_);
  and (_39724_, _02718_, _43100_);
  and (_02719_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_02720_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_02721_, _02720_, _02719_);
  and (_39725_, _02721_, _43100_);
  and (_02722_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_02723_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_02724_, _02723_, _02722_);
  and (_39726_, _02724_, _43100_);
  and (_02725_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_02726_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_02727_, _02726_, _02725_);
  and (_39727_, _02727_, _43100_);
  and (_02728_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_02729_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_02730_, _02729_, _02728_);
  and (_39728_, _02730_, _43100_);
  and (_02731_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_02732_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_02733_, _02732_, _02731_);
  and (_39729_, _02733_, _43100_);
  and (_02734_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02735_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_02736_, _02735_, _02734_);
  and (_39730_, _02736_, _43100_);
  and (_02737_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02738_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_02739_, _02738_, _02737_);
  and (_39731_, _02739_, _43100_);
  and (_02740_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02741_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_02742_, _02741_, _02740_);
  and (_39732_, _02742_, _43100_);
  and (_02743_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02744_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_02745_, _02744_, _02743_);
  and (_39733_, _02745_, _43100_);
  and (_02746_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02747_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_02748_, _02747_, _02746_);
  and (_39735_, _02748_, _43100_);
  and (_02749_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02750_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_02751_, _02750_, _02749_);
  and (_39736_, _02751_, _43100_);
  and (_02752_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02753_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_02754_, _02753_, _02752_);
  and (_39737_, _02754_, _43100_);
  and (_02755_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02756_, _42697_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02757_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_02758_, _02757_, _01922_);
  and (_02759_, _02758_, _02756_);
  or (_02760_, _02759_, _02755_);
  and (_39738_, _02760_, _43100_);
  and (_02761_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02762_, _42591_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02763_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_02764_, _02763_, _01922_);
  and (_02765_, _02764_, _02762_);
  or (_02766_, _02765_, _02761_);
  and (_39739_, _02766_, _43100_);
  and (_02767_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02768_, _42815_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02769_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_02770_, _02769_, _01922_);
  and (_02771_, _02770_, _02768_);
  or (_02772_, _02771_, _02767_);
  and (_39740_, _02772_, _43100_);
  and (_02773_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02774_, _42661_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02775_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_02776_, _02775_, _01922_);
  and (_02777_, _02776_, _02774_);
  or (_02778_, _02777_, _02773_);
  and (_39741_, _02778_, _43100_);
  and (_02779_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02780_, _42575_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02781_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_02782_, _02781_, _01922_);
  and (_02783_, _02782_, _02780_);
  or (_02784_, _02783_, _02779_);
  and (_39742_, _02784_, _43100_);
  and (_02785_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02786_, _42762_, _01929_);
  or (_02787_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_02788_, _02787_, _01922_);
  and (_02789_, _02788_, _02786_);
  or (_02790_, _02789_, _02785_);
  and (_39743_, _02790_, _43100_);
  and (_02791_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02792_, _42720_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02793_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_02794_, _02793_, _01922_);
  and (_02795_, _02794_, _02792_);
  or (_02796_, _02795_, _02791_);
  and (_39744_, _02796_, _43100_);
  and (_02797_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02798_, _42495_, _01929_);
  or (_02799_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_02800_, _02799_, _01922_);
  and (_02801_, _02800_, _02798_);
  or (_02803_, _02801_, _02797_);
  and (_39746_, _02803_, _43100_);
  and (_02804_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_02805_, _02804_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02806_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _01922_);
  and (_02808_, _02806_, _43100_);
  and (_39747_, _02808_, _02805_);
  and (_02809_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_02810_, _02809_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02811_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _01922_);
  and (_02813_, _02811_, _43100_);
  and (_39748_, _02813_, _02810_);
  and (_02814_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_02815_, _02814_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02816_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _01922_);
  and (_02818_, _02816_, _43100_);
  and (_39749_, _02818_, _02815_);
  and (_02819_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_02820_, _02819_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02821_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _01922_);
  and (_02823_, _02821_, _43100_);
  and (_39750_, _02823_, _02820_);
  and (_02824_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_02825_, _02824_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02826_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _01922_);
  and (_02828_, _02826_, _43100_);
  and (_39751_, _02828_, _02825_);
  and (_02829_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_02830_, _02829_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02831_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _01922_);
  and (_02833_, _02831_, _43100_);
  and (_39752_, _02833_, _02830_);
  and (_02835_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_02836_, _02835_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02837_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _01922_);
  and (_02838_, _02837_, _43100_);
  and (_39753_, _02838_, _02836_);
  nand (_02840_, _01936_, _31808_);
  or (_02841_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_02843_, _02841_, _43100_);
  and (_39754_, _02843_, _02840_);
  nand (_02844_, _01936_, _32495_);
  or (_02846_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_02847_, _02846_, _43100_);
  and (_39755_, _02847_, _02844_);
  nand (_02849_, _01936_, _33202_);
  or (_02850_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_02852_, _02850_, _43100_);
  and (_39757_, _02852_, _02849_);
  nand (_02854_, _01936_, _33953_);
  or (_02855_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_02857_, _02855_, _43100_);
  and (_39758_, _02857_, _02854_);
  nand (_02858_, _01936_, _34693_);
  or (_02860_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_02861_, _02860_, _43100_);
  and (_39759_, _02861_, _02858_);
  nand (_02863_, _01936_, _35520_);
  or (_02864_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_02866_, _02864_, _43100_);
  and (_39760_, _02866_, _02863_);
  nand (_02867_, _01936_, _36239_);
  or (_02868_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_02869_, _02868_, _43100_);
  and (_39761_, _02869_, _02867_);
  nand (_02870_, _01936_, _30574_);
  or (_02872_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_02874_, _02872_, _43100_);
  and (_39762_, _02874_, _02870_);
  nand (_02876_, _01936_, _38882_);
  or (_02877_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_02878_, _02877_, _43100_);
  and (_39763_, _02878_, _02876_);
  nand (_02880_, _01936_, _38916_);
  or (_02881_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_02883_, _02881_, _43100_);
  and (_39764_, _02883_, _02880_);
  nand (_02885_, _01936_, _38947_);
  or (_02887_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_02888_, _02887_, _43100_);
  and (_39765_, _02888_, _02885_);
  nand (_02890_, _01936_, _38976_);
  or (_02891_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_02892_, _02891_, _43100_);
  and (_39766_, _02892_, _02890_);
  nand (_02894_, _01936_, _39007_);
  or (_02896_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_02898_, _02896_, _43100_);
  and (_39768_, _02898_, _02894_);
  nand (_02899_, _01936_, _39041_);
  or (_02900_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_02902_, _02900_, _43100_);
  and (_39769_, _02902_, _02899_);
  nand (_02903_, _01936_, _39071_);
  or (_02905_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_02906_, _02905_, _43100_);
  and (_39770_, _02906_, _02903_);
  nor (_39980_, _42534_, rst);
  and (_02908_, _39237_, _27496_);
  and (_02909_, _02908_, _42467_);
  nand (_02911_, _02909_, _38704_);
  or (_02912_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_02913_, _02912_, _43100_);
  and (_39981_, _02913_, _02911_);
  and (_02915_, _39497_, _27496_);
  not (_02916_, _02915_);
  nor (_02918_, _02916_, _38704_);
  not (_02920_, _42467_);
  and (_02921_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_02923_, _02921_, _02920_);
  or (_02924_, _02923_, _02918_);
  or (_02926_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_02927_, _02926_, _43100_);
  and (_39982_, _02927_, _02924_);
  and (_02928_, _27003_, _27661_);
  and (_02929_, _02928_, _27496_);
  not (_02930_, _02929_);
  nor (_02932_, _02930_, _38704_);
  and (_02934_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or (_02935_, _02934_, _02920_);
  or (_02936_, _02935_, _02932_);
  or (_02938_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_02939_, _02938_, _43100_);
  and (_39983_, _02939_, _02936_);
  and (_02941_, _41582_, _27496_);
  not (_02942_, _02941_);
  nor (_02943_, _02942_, _38704_);
  and (_02946_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_02947_, _02946_, _02920_);
  or (_02948_, _02947_, _02943_);
  or (_02950_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_02951_, _02950_, _43100_);
  and (_39985_, _02951_, _02948_);
  nand (_02953_, _02909_, _38682_);
  or (_02954_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_02955_, _02954_, _43100_);
  and (_40013_, _02955_, _02953_);
  nand (_02958_, _02909_, _38672_);
  or (_02960_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_02961_, _02960_, _43100_);
  and (_40014_, _02961_, _02958_);
  nand (_02962_, _02909_, _38665_);
  or (_02964_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_02965_, _02964_, _43100_);
  and (_40015_, _02965_, _02962_);
  nand (_02967_, _02909_, _38658_);
  or (_02968_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_02970_, _02968_, _43100_);
  and (_40016_, _02970_, _02967_);
  nand (_02972_, _02909_, _38650_);
  or (_02973_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_02975_, _02973_, _43100_);
  and (_40017_, _02975_, _02972_);
  nand (_02976_, _02909_, _38642_);
  or (_02978_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_02979_, _02978_, _43100_);
  and (_40018_, _02979_, _02976_);
  nand (_02982_, _02909_, _38635_);
  or (_02983_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_02984_, _02983_, _43100_);
  and (_40019_, _02984_, _02982_);
  nor (_02986_, _02916_, _38682_);
  and (_02988_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_02989_, _02988_, _02920_);
  or (_02990_, _02989_, _02986_);
  or (_02991_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_02993_, _02991_, _43100_);
  and (_40021_, _02993_, _02990_);
  nor (_02995_, _02916_, _38672_);
  and (_02997_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_02998_, _02997_, _02920_);
  or (_02999_, _02998_, _02995_);
  or (_03001_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_03002_, _03001_, _43100_);
  and (_40022_, _03002_, _02999_);
  nor (_03004_, _02916_, _38665_);
  and (_03005_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_03007_, _03005_, _02920_);
  or (_03009_, _03007_, _03004_);
  or (_03010_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_03011_, _03010_, _43100_);
  and (_40023_, _03011_, _03009_);
  nor (_03013_, _02916_, _38658_);
  and (_03014_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_03016_, _03014_, _02920_);
  or (_03017_, _03016_, _03013_);
  or (_03019_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_03021_, _03019_, _43100_);
  and (_40024_, _03021_, _03017_);
  nor (_03022_, _02916_, _38650_);
  and (_03024_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_03025_, _03024_, _02920_);
  or (_03026_, _03025_, _03022_);
  or (_03028_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_03029_, _03028_, _43100_);
  and (_40025_, _03029_, _03026_);
  nor (_03031_, _02916_, _38642_);
  and (_03032_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_03033_, _03032_, _02920_);
  or (_03035_, _03033_, _03031_);
  or (_03036_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_03037_, _03036_, _43100_);
  and (_40026_, _03037_, _03035_);
  nor (_03039_, _02916_, _38635_);
  and (_03040_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_03042_, _03040_, _02920_);
  or (_03043_, _03042_, _03039_);
  or (_03044_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_03046_, _03044_, _43100_);
  and (_40027_, _03046_, _03043_);
  or (_03048_, _02929_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand (_03049_, _02929_, _38682_);
  and (_03050_, _03049_, _03048_);
  or (_03051_, _03050_, _02920_);
  or (_03052_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_03053_, _03052_, _43100_);
  and (_40028_, _03053_, _03051_);
  nor (_03055_, _02930_, _38672_);
  and (_03056_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_03057_, _03056_, _02920_);
  or (_03059_, _03057_, _03055_);
  or (_03060_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_03061_, _03060_, _43100_);
  and (_40029_, _03061_, _03059_);
  nor (_03063_, _02930_, _38665_);
  and (_03064_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or (_03066_, _03064_, _02920_);
  or (_03067_, _03066_, _03063_);
  or (_03068_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_03070_, _03068_, _43100_);
  and (_40030_, _03070_, _03067_);
  not (_03071_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_03073_, _02929_, _42467_);
  nor (_03074_, _03073_, _03071_);
  and (_03075_, _03073_, _40346_);
  or (_03077_, _03075_, _03074_);
  and (_40032_, _03077_, _43100_);
  nor (_03079_, _02930_, _38650_);
  and (_03080_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or (_03081_, _03080_, _02920_);
  or (_03082_, _03081_, _03079_);
  or (_03084_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_03085_, _03084_, _43100_);
  and (_40033_, _03085_, _03082_);
  nor (_03087_, _02930_, _38642_);
  and (_03088_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_03089_, _03088_, _02920_);
  or (_03091_, _03089_, _03087_);
  or (_03092_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_03093_, _03092_, _43100_);
  and (_40034_, _03093_, _03091_);
  nor (_03095_, _02930_, _38635_);
  and (_03096_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_03098_, _03096_, _02920_);
  or (_03099_, _03098_, _03095_);
  or (_03100_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_03102_, _03100_, _43100_);
  and (_40035_, _03102_, _03099_);
  and (_03103_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_03105_, _02942_, _38682_);
  or (_03106_, _03105_, _02920_);
  or (_03108_, _03106_, _03103_);
  or (_03109_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_03110_, _03109_, _43100_);
  and (_40036_, _03110_, _03108_);
  nor (_03112_, _02942_, _38672_);
  and (_03113_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_03114_, _03113_, _02920_);
  or (_03116_, _03114_, _03112_);
  or (_03117_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_03118_, _03117_, _43100_);
  and (_40037_, _03118_, _03116_);
  nor (_03120_, _02942_, _38665_);
  and (_03121_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_03123_, _03121_, _02920_);
  or (_03124_, _03123_, _03120_);
  or (_03125_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_03128_, _03125_, _43100_);
  and (_40038_, _03128_, _03124_);
  nor (_03129_, _02942_, _38658_);
  and (_03131_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_03132_, _03131_, _02920_);
  or (_03133_, _03132_, _03129_);
  or (_03135_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_03136_, _03135_, _43100_);
  and (_40039_, _03136_, _03133_);
  nor (_03138_, _02942_, _38650_);
  and (_03139_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or (_03140_, _03139_, _02920_);
  or (_03142_, _03140_, _03138_);
  or (_03143_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_03144_, _03143_, _43100_);
  and (_40040_, _03144_, _03142_);
  nor (_03146_, _02942_, _38642_);
  and (_03147_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_03149_, _03147_, _02920_);
  or (_03150_, _03149_, _03146_);
  or (_03151_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_03153_, _03151_, _43100_);
  and (_40041_, _03153_, _03150_);
  nor (_03154_, _02942_, _38635_);
  and (_03156_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_03157_, _03156_, _02920_);
  or (_03158_, _03157_, _03154_);
  or (_03160_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_03161_, _03160_, _43100_);
  and (_40043_, _03161_, _03158_);
  not (_03163_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_03164_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_03166_, _03164_, _03163_);
  and (_03167_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _43100_);
  and (_40070_, _03167_, _03166_);
  nor (_03168_, _03166_, rst);
  nand (_03169_, _03164_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03171_, _03164_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03172_, _03171_, _03169_);
  and (_40072_, _03172_, _03168_);
  nor (_03174_, _42743_, _42787_);
  not (_03175_, _42521_);
  and (_03176_, _42579_, _03175_);
  and (_03178_, _03176_, _03174_);
  and (_03179_, _03178_, _42665_);
  and (_03180_, _03179_, _39236_);
  nor (_03182_, _03180_, _01344_);
  nor (_03183_, _42743_, _42788_);
  nor (_03184_, _42666_, _42579_);
  and (_03186_, _03184_, _03175_);
  and (_03187_, _03186_, _03183_);
  not (_03188_, _42823_);
  nor (_03190_, _39326_, _39314_);
  and (_03191_, _39326_, _39314_);
  nor (_03192_, _03191_, _03190_);
  nor (_03194_, _39383_, _39338_);
  and (_03195_, _39383_, _39338_);
  nor (_03197_, _03195_, _03194_);
  nor (_03198_, _03197_, _03192_);
  and (_03199_, _03197_, _03192_);
  or (_03200_, _03199_, _03198_);
  and (_03202_, _39407_, _39395_);
  nor (_03203_, _39407_, _39395_);
  nor (_03204_, _03203_, _03202_);
  nor (_03206_, _39419_, _39260_);
  and (_03207_, _39419_, _39260_);
  nor (_03208_, _03207_, _03206_);
  or (_03210_, _03208_, _03204_);
  nand (_03211_, _03208_, _03204_);
  and (_03212_, _03211_, _03210_);
  nor (_03214_, _03212_, _03200_);
  and (_03215_, _03212_, _03200_);
  nor (_03216_, _03215_, _03214_);
  or (_03218_, _03216_, _03188_);
  and (_03219_, _42701_, _42617_);
  or (_03220_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03222_, _03220_, _03219_);
  and (_03223_, _03222_, _03218_);
  nor (_03224_, _42701_, _42617_);
  and (_03226_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  not (_03227_, _42701_);
  and (_03229_, _03227_, _42617_);
  and (_03230_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_03231_, _03230_, _03226_);
  and (_03232_, _03231_, _03188_);
  or (_03234_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_03235_, _03227_, _42617_);
  or (_03236_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_03238_, _03236_, _03235_);
  and (_03239_, _03238_, _03234_);
  and (_03240_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_03242_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_03243_, _03242_, _03240_);
  and (_03244_, _03243_, _42823_);
  or (_03246_, _03244_, _03239_);
  or (_03247_, _03246_, _03232_);
  or (_03248_, _03247_, _03223_);
  and (_03250_, _03248_, _03187_);
  nor (_03251_, _03187_, _28636_);
  and (_03252_, _42743_, _03175_);
  nand (_03254_, _03252_, _42666_);
  not (_03255_, _03183_);
  nand (_03256_, _03186_, _03255_);
  and (_03258_, _03256_, _03254_);
  and (_03259_, _03258_, _03251_);
  and (_03261_, _03176_, _42666_);
  and (_03262_, _03261_, _03183_);
  nor (_03263_, _03262_, _03179_);
  and (_03264_, _42743_, _42787_);
  and (_03266_, _03264_, _03176_);
  and (_03267_, _03266_, _42665_);
  and (_03268_, _42743_, _42788_);
  and (_03270_, _03268_, _03176_);
  and (_03271_, _03270_, _42665_);
  nor (_03272_, _03271_, _03267_);
  and (_03274_, _03272_, _03263_);
  and (_03275_, _03274_, _03259_);
  and (_03276_, _01425_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  nor (_03278_, _00818_, _38521_);
  and (_03279_, _38443_, _38488_);
  nor (_03280_, _03279_, _00933_);
  and (_03282_, _03280_, _03278_);
  not (_03283_, _38515_);
  nor (_03284_, _00913_, _38509_);
  and (_03286_, _03284_, _03283_);
  and (_03287_, _03286_, _00820_);
  and (_03288_, _03287_, _03282_);
  and (_03290_, _01091_, _00753_);
  and (_03291_, _03290_, _03288_);
  and (_03292_, _03291_, _38546_);
  nor (_03293_, _03292_, _36466_);
  or (_03294_, _03293_, p2_in[5]);
  not (_03295_, _03293_);
  or (_03296_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03297_, _03296_, _03294_);
  and (_03298_, _03297_, _03188_);
  or (_03299_, _03293_, p2_in[1]);
  or (_03300_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_03301_, _03300_, _03299_);
  and (_03302_, _03301_, _42823_);
  or (_03303_, _03302_, _03298_);
  and (_03304_, _03303_, _03229_);
  or (_03305_, _03293_, p2_in[2]);
  or (_03306_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03307_, _03306_, _03305_);
  or (_03308_, _03307_, _03188_);
  or (_03309_, _03293_, p2_in[6]);
  or (_03310_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03311_, _03310_, _03309_);
  or (_03312_, _03311_, _42823_);
  and (_03313_, _03312_, _03235_);
  and (_03314_, _03313_, _03308_);
  or (_03315_, _03293_, p2_in[4]);
  or (_03316_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_03317_, _03316_, _03315_);
  and (_03318_, _03317_, _03188_);
  nor (_03319_, _03293_, p2_in[0]);
  and (_03320_, _03293_, _39860_);
  nor (_03321_, _03320_, _03319_);
  and (_03322_, _03321_, _42823_);
  or (_03323_, _03322_, _03318_);
  and (_03324_, _03323_, _03219_);
  or (_03325_, _03293_, p2_in[3]);
  or (_03326_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03327_, _03326_, _03325_);
  or (_03328_, _03327_, _03188_);
  or (_03329_, _03293_, p2_in[7]);
  or (_03330_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_03331_, _03330_, _03329_);
  or (_03332_, _03331_, _42823_);
  and (_03333_, _03332_, _03224_);
  and (_03334_, _03333_, _03328_);
  or (_03335_, _03334_, _03324_);
  or (_03336_, _03335_, _03314_);
  or (_03337_, _03336_, _03304_);
  and (_03338_, _03337_, _03271_);
  and (_03339_, _03219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03340_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_03341_, _03340_, _03339_);
  and (_03342_, _03235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_03343_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_03344_, _03343_, _03342_);
  or (_03345_, _03344_, _03341_);
  and (_03346_, _03345_, _03188_);
  and (_03347_, _03219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_03348_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03349_, _03348_, _03347_);
  and (_03350_, _03235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_03351_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_03352_, _03351_, _03350_);
  or (_03353_, _03352_, _03349_);
  and (_03354_, _03353_, _42823_);
  or (_03355_, _03354_, _03346_);
  and (_03356_, _03355_, _03262_);
  or (_03357_, _03356_, _03338_);
  or (_03358_, _03357_, _03276_);
  or (_03359_, _03358_, _03275_);
  nor (_03360_, _42823_, _40899_);
  and (_03361_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_03362_, _03361_, _03360_);
  and (_03364_, _03362_, _03219_);
  or (_03365_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_03366_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03367_, _03366_, _03224_);
  and (_03368_, _03367_, _03365_);
  or (_03369_, _03368_, _03364_);
  and (_03370_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03371_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_03372_, _03371_, _03370_);
  and (_03373_, _03372_, _03235_);
  or (_03374_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_03375_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_03376_, _03375_, _03229_);
  and (_03377_, _03376_, _03374_);
  or (_03378_, _03377_, _03373_);
  or (_03379_, _03378_, _03369_);
  and (_03380_, _03379_, _03268_);
  and (_03381_, _03219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_03382_, _03235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_03383_, _03382_, _03381_);
  and (_03384_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_03385_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_03386_, _03385_, _03384_);
  or (_03387_, _03386_, _03383_);
  and (_03388_, _03387_, _42823_);
  and (_03389_, _03219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_03390_, _03235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_03391_, _03390_, _03389_);
  and (_03392_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03393_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03394_, _03393_, _03392_);
  or (_03395_, _03394_, _03391_);
  and (_03396_, _03395_, _03188_);
  or (_03397_, _03396_, _03388_);
  and (_03398_, _03397_, _03264_);
  or (_03399_, _03398_, _03380_);
  and (_03400_, _03399_, _03261_);
  and (_03401_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03402_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_03403_, _03402_, _03401_);
  and (_03404_, _03403_, _03188_);
  and (_03405_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_03406_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03407_, _03406_, _03405_);
  and (_03408_, _03407_, _03219_);
  and (_03409_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_03410_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03411_, _03410_, _03409_);
  and (_03412_, _03411_, _03235_);
  or (_03413_, _03412_, _03408_);
  and (_03414_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_03415_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03416_, _03415_, _03414_);
  and (_03417_, _03416_, _42823_);
  or (_03418_, _03417_, _03413_);
  or (_03419_, _03418_, _03404_);
  and (_03420_, _03419_, _03179_);
  or (_03421_, _42665_, _42521_);
  nor (_03422_, _03421_, _42579_);
  and (_03423_, _03422_, _03264_);
  nor (_03424_, _42823_, _41473_);
  and (_03425_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_03426_, _03425_, _03424_);
  and (_03427_, _03426_, _03224_);
  or (_03428_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand (_03429_, _42823_, _41490_);
  and (_03430_, _03429_, _03219_);
  and (_03431_, _03430_, _03428_);
  or (_03432_, _03431_, _03427_);
  nor (_03433_, _42823_, _41899_);
  and (_03434_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03435_, _03434_, _03433_);
  and (_03436_, _03435_, _03229_);
  nand (_03437_, _42823_, _41924_);
  or (_03438_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_03439_, _03438_, _03235_);
  and (_03440_, _03439_, _03437_);
  or (_03441_, _03440_, _03436_);
  or (_03442_, _03441_, _03432_);
  and (_03443_, _03442_, _03423_);
  or (_03444_, _03293_, p0_in[5]);
  or (_03445_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03446_, _03445_, _03444_);
  and (_03447_, _03446_, _03188_);
  or (_03448_, _03293_, p0_in[1]);
  or (_03449_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03450_, _03449_, _03448_);
  and (_03451_, _03450_, _42823_);
  or (_03452_, _03451_, _03447_);
  and (_03453_, _03452_, _03229_);
  or (_03454_, _03293_, p0_in[2]);
  nand (_03455_, _03293_, _39510_);
  and (_03456_, _03455_, _03454_);
  or (_03457_, _03456_, _03188_);
  or (_03458_, _03293_, p0_in[6]);
  or (_03459_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03460_, _03459_, _03458_);
  or (_03461_, _03460_, _42823_);
  and (_03462_, _03461_, _03235_);
  and (_03463_, _03462_, _03457_);
  or (_03464_, _03293_, p0_in[4]);
  or (_03465_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_03466_, _03465_, _03464_);
  and (_03467_, _03466_, _03188_);
  nor (_03468_, _03293_, p0_in[0]);
  and (_03469_, _03293_, _39493_);
  nor (_03470_, _03469_, _03468_);
  and (_03471_, _03470_, _42823_);
  or (_03472_, _03471_, _03467_);
  and (_03473_, _03472_, _03219_);
  or (_03474_, _03293_, p0_in[3]);
  or (_03475_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03476_, _03475_, _03474_);
  or (_03477_, _03476_, _03188_);
  or (_03478_, _03293_, p0_in[7]);
  or (_03479_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03480_, _03479_, _03478_);
  or (_03481_, _03480_, _42823_);
  and (_03482_, _03481_, _03224_);
  and (_03483_, _03482_, _03477_);
  or (_03484_, _03483_, _03473_);
  or (_03485_, _03484_, _03463_);
  or (_03486_, _03485_, _03453_);
  and (_03487_, _03486_, _03267_);
  or (_03488_, _03487_, _03443_);
  or (_03489_, _03488_, _03420_);
  or (_03490_, _03489_, _03400_);
  and (_03491_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_03492_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03493_, _03492_, _03491_);
  and (_03494_, _03493_, _03224_);
  or (_03495_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nand (_03496_, _42823_, _40918_);
  and (_03497_, _03496_, _03219_);
  and (_03498_, _03497_, _03495_);
  or (_03499_, _03498_, _03494_);
  nor (_03500_, _42823_, _40930_);
  and (_03501_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_03502_, _03501_, _03500_);
  and (_03503_, _03502_, _03229_);
  nand (_03504_, _42823_, _40923_);
  or (_03505_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03506_, _03505_, _03235_);
  and (_03507_, _03506_, _03504_);
  or (_03508_, _03507_, _03503_);
  or (_03509_, _03508_, _03499_);
  and (_03510_, _03509_, _03422_);
  or (_03511_, _03293_, p3_in[7]);
  or (_03512_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_03513_, _03512_, _03511_);
  and (_03514_, _03513_, _03188_);
  or (_03515_, _03293_, p3_in[3]);
  or (_03516_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03517_, _03516_, _03515_);
  and (_03518_, _03517_, _42823_);
  or (_03519_, _03518_, _03514_);
  and (_03520_, _03519_, _03224_);
  nor (_03521_, _03293_, p3_in[0]);
  and (_03522_, _03293_, _39947_);
  nor (_03523_, _03522_, _03521_);
  or (_03524_, _03523_, _03188_);
  or (_03525_, _03293_, p3_in[4]);
  or (_03526_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_03527_, _03526_, _03525_);
  or (_03528_, _03527_, _42823_);
  and (_03529_, _03528_, _03219_);
  and (_03530_, _03529_, _03524_);
  or (_03531_, _03530_, _03520_);
  or (_03532_, _03293_, p3_in[6]);
  or (_03533_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03534_, _03533_, _03532_);
  and (_03535_, _03534_, _03188_);
  or (_03536_, _03293_, p3_in[2]);
  or (_03537_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03538_, _03537_, _03536_);
  and (_03539_, _03538_, _42823_);
  or (_03540_, _03539_, _03535_);
  and (_03541_, _03540_, _03235_);
  or (_03542_, _03293_, p3_in[1]);
  or (_03543_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03544_, _03543_, _03542_);
  or (_03545_, _03544_, _03188_);
  or (_03546_, _03293_, p3_in[5]);
  or (_03547_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03548_, _03547_, _03546_);
  or (_03549_, _03548_, _42823_);
  and (_03550_, _03549_, _03229_);
  and (_03551_, _03550_, _03545_);
  or (_03552_, _03551_, _03541_);
  or (_03553_, _03552_, _03531_);
  and (_03554_, _03553_, _03186_);
  or (_03555_, _03554_, _03510_);
  and (_03556_, _03555_, _03268_);
  nor (_03557_, _42823_, _30661_);
  and (_03558_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_03559_, _03558_, _03557_);
  and (_03560_, _03559_, _03224_);
  or (_03561_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_03562_, _42823_, _31831_);
  and (_03563_, _03562_, _03219_);
  and (_03565_, _03563_, _03561_);
  or (_03566_, _03565_, _03560_);
  nor (_03567_, _42823_, _35553_);
  and (_03568_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_03569_, _03568_, _03567_);
  and (_03570_, _03569_, _03229_);
  nand (_03571_, _42823_, _33235_);
  or (_03572_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_03573_, _03572_, _03235_);
  and (_03574_, _03573_, _03571_);
  or (_03575_, _03574_, _03570_);
  or (_03576_, _03575_, _03566_);
  and (_03577_, _03576_, _03174_);
  or (_03578_, _03293_, p1_in[5]);
  or (_03579_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03580_, _03579_, _03578_);
  and (_03581_, _03580_, _03188_);
  or (_03582_, _03293_, p1_in[1]);
  or (_03583_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03584_, _03583_, _03582_);
  and (_03585_, _03584_, _42823_);
  or (_03586_, _03585_, _03581_);
  and (_03587_, _03586_, _03229_);
  or (_03588_, _03293_, p1_in[2]);
  or (_03589_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03590_, _03589_, _03588_);
  or (_03591_, _03590_, _03188_);
  or (_03592_, _03293_, p1_in[6]);
  or (_03593_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03594_, _03593_, _03592_);
  or (_03595_, _03594_, _42823_);
  and (_03596_, _03595_, _03235_);
  and (_03597_, _03596_, _03591_);
  or (_03598_, _03293_, p1_in[4]);
  or (_03599_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03600_, _03599_, _03598_);
  and (_03601_, _03600_, _03188_);
  nor (_03602_, _03293_, p1_in[0]);
  and (_03603_, _03293_, _39779_);
  nor (_03604_, _03603_, _03602_);
  and (_03605_, _03604_, _42823_);
  or (_03606_, _03605_, _03601_);
  and (_03607_, _03606_, _03219_);
  or (_03608_, _03293_, p1_in[3]);
  or (_03609_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03610_, _03609_, _03608_);
  or (_03611_, _03610_, _03188_);
  or (_03612_, _03293_, p1_in[7]);
  or (_03613_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_03614_, _03613_, _03612_);
  or (_03615_, _03614_, _42823_);
  and (_03616_, _03615_, _03224_);
  and (_03617_, _03616_, _03611_);
  or (_03618_, _03617_, _03607_);
  or (_03619_, _03618_, _03597_);
  or (_03620_, _03619_, _03587_);
  and (_03621_, _03620_, _03264_);
  or (_03622_, _03621_, _03577_);
  and (_03623_, _03622_, _03186_);
  or (_03624_, _03623_, _03556_);
  or (_03625_, _03624_, _03490_);
  or (_03626_, _03625_, _03359_);
  or (_03627_, _03626_, _03250_);
  nand (_03628_, _03276_, _31265_);
  nand (_03629_, _03628_, _03627_);
  nand (_03630_, _03629_, _03182_);
  and (_03631_, _03219_, _38683_);
  or (_03632_, _03631_, _03188_);
  and (_03633_, _03224_, _40346_);
  and (_03634_, _03229_, _41428_);
  and (_03635_, _03235_, _40334_);
  or (_03636_, _03635_, _03634_);
  or (_03637_, _03636_, _03633_);
  or (_03638_, _03637_, _03632_);
  and (_03639_, _03219_, _40357_);
  or (_03640_, _03639_, _42823_);
  and (_03641_, _03224_, _40145_);
  and (_03642_, _03229_, _40370_);
  and (_03643_, _03235_, _40383_);
  or (_03644_, _03643_, _03642_);
  or (_03645_, _03644_, _03641_);
  or (_03646_, _03645_, _03640_);
  and (_03647_, _03646_, _03638_);
  or (_03648_, _03647_, _03182_);
  and (_03649_, _03648_, _43100_);
  and (_40073_, _03649_, _03630_);
  and (_03650_, _42665_, _42823_);
  and (_03651_, _03650_, _03219_);
  and (_03652_, _03651_, _03178_);
  and (_03653_, _03652_, _39231_);
  nor (_03654_, _42788_, _42579_);
  nor (_03655_, _42743_, _42521_);
  and (_03656_, _03651_, _03655_);
  and (_03657_, _03656_, _03654_);
  and (_03658_, _03657_, _39106_);
  nor (_03659_, _03658_, _03653_);
  and (_03660_, _03650_, _03224_);
  and (_03661_, _03660_, _03266_);
  nand (_03662_, _03661_, _38755_);
  and (_03663_, _03662_, _03659_);
  nor (_03664_, _03663_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_03665_, _03664_);
  and (_03666_, _03652_, _39236_);
  not (_03667_, _39247_);
  and (_03668_, _03224_, _03188_);
  nor (_03669_, _03668_, _03667_);
  and (_03670_, _03669_, _01342_);
  nor (_03671_, _03670_, _03666_);
  and (_03672_, _03671_, _01428_);
  and (_03673_, _03672_, _03665_);
  and (_03674_, _03266_, _03235_);
  and (_03675_, _03674_, _03650_);
  and (_03676_, _03675_, _38755_);
  or (_03677_, _03676_, rst);
  nor (_40074_, _03677_, _03673_);
  nand (_03678_, _03676_, _30574_);
  and (_03679_, _03183_, _03176_);
  nor (_03680_, _42665_, _42823_);
  and (_03681_, _03680_, _03219_);
  and (_03682_, _03681_, _03679_);
  and (_03683_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_03684_, _42666_, _42823_);
  and (_03685_, _03684_, _03219_);
  and (_03686_, _03685_, _03679_);
  and (_03687_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_03688_, _03687_, _03683_);
  and (_03689_, _03684_, _03235_);
  and (_03690_, _03689_, _03679_);
  and (_03691_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_03692_, _03680_, _03229_);
  and (_03693_, _03692_, _03679_);
  and (_03694_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_03695_, _03694_, _03691_);
  or (_03696_, _03695_, _03688_);
  and (_03697_, _03684_, _03224_);
  and (_03698_, _03697_, _03679_);
  and (_03699_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_03700_, _03685_, _03266_);
  and (_03701_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_03702_, _03701_, _03699_);
  and (_03703_, _03685_, _03270_);
  and (_03704_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03705_, _03668_, _42665_);
  nor (_03706_, _42787_, _42579_);
  and (_03707_, _03706_, _03252_);
  and (_03708_, _03707_, _03705_);
  and (_03709_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_03710_, _03709_, _03704_);
  or (_03711_, _03710_, _03702_);
  or (_03712_, _03711_, _03696_);
  and (_03713_, _03684_, _03229_);
  and (_03714_, _03713_, _03266_);
  and (_03715_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_03716_, _03697_, _03266_);
  and (_03717_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or (_03718_, _03717_, _03715_);
  and (_03719_, _03692_, _03266_);
  and (_03720_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_03721_, _03689_, _03266_);
  and (_03722_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_03723_, _03722_, _03720_);
  or (_03724_, _03723_, _03718_);
  and (_03725_, _03654_, _03252_);
  and (_03726_, _03725_, _03713_);
  and (_03727_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_03728_, _03725_, _03685_);
  and (_03729_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_03730_, _03729_, _03727_);
  and (_03731_, _03681_, _03266_);
  and (_03732_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_03733_, _03668_, _03267_);
  and (_03734_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_03735_, _03734_, _03732_);
  or (_03736_, _03735_, _03730_);
  or (_03737_, _03736_, _03724_);
  or (_03738_, _03737_, _03712_);
  and (_03739_, _03266_, _03229_);
  and (_03740_, _03739_, _03650_);
  and (_03741_, _03740_, _38706_);
  and (_03742_, _03706_, _03656_);
  and (_03743_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_03744_, _03743_, _03741_);
  and (_03745_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_03746_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_03747_, _03746_, _03745_);
  or (_03748_, _03747_, _03744_);
  and (_03749_, _03651_, _03270_);
  and (_03750_, _03749_, _03331_);
  and (_03751_, _03707_, _03651_);
  and (_03752_, _03751_, _03513_);
  or (_03753_, _03752_, _03750_);
  and (_03754_, _03651_, _03266_);
  and (_03755_, _03754_, _03480_);
  and (_03756_, _03725_, _03651_);
  and (_03757_, _03756_, _03614_);
  or (_03758_, _03757_, _03755_);
  or (_03759_, _03758_, _03753_);
  or (_03760_, _03759_, _03748_);
  and (_03761_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03762_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03764_, _03762_, _03761_);
  or (_03765_, _03764_, _03760_);
  or (_03766_, _03765_, _03738_);
  and (_03767_, _03651_, _03252_);
  or (_03768_, _03742_, _03767_);
  or (_03769_, _03768_, _03740_);
  and (_03770_, _03266_, _03224_);
  nand (_03771_, _03684_, _03770_);
  nor (_03772_, _03726_, _03731_);
  nor (_03773_, _03719_, _03728_);
  and (_03774_, _03773_, _03772_);
  nand (_03775_, _03774_, _03771_);
  or (_03776_, _03775_, _03769_);
  or (_03777_, _03708_, _03652_);
  or (_03778_, _03733_, _03657_);
  or (_03779_, _03778_, _03777_);
  and (_03780_, _03770_, _03650_);
  or (_03781_, _03698_, _03690_);
  or (_03782_, _03693_, _03700_);
  or (_03783_, _03782_, _03781_);
  or (_03784_, _03783_, _03780_);
  or (_03785_, _03784_, _03779_);
  nand (_03786_, _03684_, _03674_);
  nor (_03787_, _03703_, _03714_);
  nand (_03788_, _03787_, _03786_);
  and (_03789_, _03262_, _03219_);
  or (_03790_, _03789_, _03675_);
  or (_03791_, _03790_, _03788_);
  or (_03792_, _03791_, _03785_);
  or (_03793_, _03792_, _03776_);
  nand (_03794_, _03793_, _03673_);
  and (_03795_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_03796_, _03795_, _03766_);
  or (_03797_, _03673_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_03798_, _03797_, _03796_);
  or (_03799_, _03798_, _03676_);
  and (_03800_, _03799_, _43100_);
  and (_40075_, _03800_, _03678_);
  nor (_40156_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_03801_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_03802_, _03164_, rst);
  and (_40157_, _03802_, _03801_);
  nor (_03803_, _03164_, _03163_);
  or (_03804_, _03803_, _03166_);
  and (_03805_, _03169_, _43100_);
  and (_40158_, _03805_, _03804_);
  not (_03806_, _03673_);
  nand (_03807_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_03808_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_03809_, _03808_, _03807_);
  nand (_03810_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_03811_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_03812_, _03811_, _03810_);
  and (_03813_, _03812_, _03809_);
  nand (_03814_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_03815_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_03816_, _03815_, _03814_);
  nand (_03817_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_03818_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_03819_, _03818_, _03817_);
  and (_03820_, _03819_, _03816_);
  and (_03821_, _03820_, _03813_);
  nand (_03822_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_03823_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_03824_, _03823_, _03822_);
  nand (_03825_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_03826_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_03827_, _03826_, _03825_);
  and (_03828_, _03827_, _03824_);
  nand (_03829_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand (_03830_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_03831_, _03830_, _03829_);
  nand (_03832_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_03833_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_03834_, _03833_, _03832_);
  and (_03835_, _03834_, _03831_);
  and (_03836_, _03835_, _03828_);
  and (_03837_, _03836_, _03821_);
  nand (_03838_, _03740_, _42686_);
  nand (_03839_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_03840_, _03839_, _03838_);
  nand (_03841_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_03842_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_03843_, _03842_, _03841_);
  and (_03844_, _03843_, _03840_);
  nand (_03845_, _03749_, _03321_);
  nand (_03846_, _03751_, _03523_);
  and (_03847_, _03846_, _03845_);
  nand (_03848_, _03756_, _03604_);
  nand (_03849_, _03754_, _03470_);
  and (_03850_, _03849_, _03848_);
  and (_03851_, _03850_, _03847_);
  and (_03852_, _03851_, _03844_);
  nand (_03853_, _03657_, _03216_);
  nand (_03854_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_03855_, _03854_, _03853_);
  and (_03856_, _03855_, _03852_);
  and (_03857_, _03856_, _03837_);
  nor (_03858_, _03857_, _03806_);
  and (_03859_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or (_03860_, _03859_, _03676_);
  or (_03861_, _03860_, _03858_);
  nand (_03862_, _03676_, _31808_);
  and (_03863_, _03862_, _43100_);
  and (_40159_, _03863_, _03861_);
  nand (_03864_, _03676_, _32495_);
  and (_03865_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_03866_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_03867_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03868_, _03867_, _03866_);
  and (_03869_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_03870_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_03871_, _03870_, _03869_);
  or (_03872_, _03871_, _03868_);
  and (_03873_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_03874_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_03875_, _03874_, _03873_);
  and (_03876_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_03877_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_03878_, _03877_, _03876_);
  or (_03879_, _03878_, _03875_);
  or (_03880_, _03879_, _03872_);
  and (_03881_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_03882_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_03883_, _03882_, _03881_);
  and (_03884_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_03885_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_03886_, _03885_, _03884_);
  or (_03887_, _03886_, _03883_);
  and (_03888_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_03889_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03890_, _03889_, _03888_);
  and (_03891_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_03892_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_03893_, _03892_, _03891_);
  or (_03894_, _03893_, _03890_);
  or (_03895_, _03894_, _03887_);
  or (_03896_, _03895_, _03880_);
  and (_03897_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_03898_, _03740_, _42595_);
  or (_03899_, _03898_, _03897_);
  and (_03900_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_03901_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_03902_, _03901_, _03900_);
  or (_03903_, _03902_, _03899_);
  and (_03904_, _03749_, _03301_);
  and (_03905_, _03751_, _03544_);
  or (_03906_, _03905_, _03904_);
  and (_03907_, _03756_, _03584_);
  and (_03908_, _03754_, _03450_);
  or (_03909_, _03908_, _03907_);
  or (_03910_, _03909_, _03906_);
  or (_03911_, _03910_, _03903_);
  and (_03912_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_03913_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_03914_, _03913_, _03912_);
  or (_03915_, _03914_, _03911_);
  or (_03916_, _03915_, _03896_);
  and (_03917_, _03916_, _03673_);
  or (_03918_, _03917_, _03865_);
  or (_03919_, _03918_, _03676_);
  and (_03920_, _03919_, _43100_);
  and (_40161_, _03920_, _03864_);
  nand (_03921_, _03676_, _33202_);
  and (_03922_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_03923_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_03924_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_03925_, _03924_, _03923_);
  and (_03926_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_03927_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_03928_, _03927_, _03926_);
  or (_03929_, _03928_, _03925_);
  and (_03930_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_03931_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_03932_, _03931_, _03930_);
  and (_03933_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_03934_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03935_, _03934_, _03933_);
  or (_03936_, _03935_, _03932_);
  or (_03937_, _03936_, _03929_);
  and (_03938_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_03939_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_03940_, _03939_, _03938_);
  and (_03941_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_03942_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_03943_, _03942_, _03941_);
  or (_03944_, _03943_, _03940_);
  and (_03945_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_03946_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_03947_, _03946_, _03945_);
  and (_03948_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_03949_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_03950_, _03949_, _03948_);
  or (_03951_, _03950_, _03947_);
  or (_03952_, _03951_, _03944_);
  or (_03953_, _03952_, _03937_);
  and (_03954_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_03955_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03956_, _03955_, _03954_);
  and (_03957_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_03959_, _03740_, _42819_);
  or (_03960_, _03959_, _03957_);
  and (_03961_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_03962_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_03963_, _03962_, _03961_);
  or (_03964_, _03963_, _03960_);
  and (_03965_, _03749_, _03307_);
  and (_03966_, _03751_, _03538_);
  or (_03967_, _03966_, _03965_);
  and (_03968_, _03754_, _03456_);
  and (_03969_, _03756_, _03590_);
  or (_03970_, _03969_, _03968_);
  or (_03971_, _03970_, _03967_);
  or (_03972_, _03971_, _03964_);
  or (_03973_, _03972_, _03956_);
  or (_03974_, _03973_, _03953_);
  and (_03975_, _03974_, _03673_);
  or (_03976_, _03975_, _03922_);
  or (_03977_, _03976_, _03676_);
  and (_03978_, _03977_, _43100_);
  and (_40162_, _03978_, _03921_);
  nand (_03979_, _03676_, _33953_);
  and (_03980_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_03981_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_03982_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_03983_, _03982_, _03981_);
  and (_03984_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_03985_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_03986_, _03985_, _03984_);
  or (_03987_, _03986_, _03983_);
  and (_03988_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_03989_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_03990_, _03989_, _03988_);
  and (_03991_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03992_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03993_, _03992_, _03991_);
  or (_03994_, _03993_, _03990_);
  or (_03995_, _03994_, _03987_);
  and (_03996_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_03997_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_03998_, _03997_, _03996_);
  and (_03999_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_04000_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_04001_, _04000_, _03999_);
  or (_04002_, _04001_, _03998_);
  and (_04003_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_04004_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_04005_, _04004_, _04003_);
  and (_04006_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_04007_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_04008_, _04007_, _04006_);
  or (_04009_, _04008_, _04005_);
  or (_04010_, _04009_, _04002_);
  or (_04011_, _04010_, _03995_);
  and (_04012_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_04013_, _03740_, _42650_);
  or (_04014_, _04013_, _04012_);
  and (_04015_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_04016_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_04017_, _04016_, _04015_);
  or (_04018_, _04017_, _04014_);
  and (_04019_, _03749_, _03327_);
  and (_04020_, _03751_, _03517_);
  or (_04021_, _04020_, _04019_);
  and (_04022_, _03756_, _03610_);
  and (_04023_, _03754_, _03476_);
  or (_04024_, _04023_, _04022_);
  or (_04025_, _04024_, _04021_);
  or (_04026_, _04025_, _04018_);
  and (_04027_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_04028_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_04029_, _04028_, _04027_);
  or (_04030_, _04029_, _04026_);
  or (_04031_, _04030_, _04011_);
  and (_04032_, _04031_, _03673_);
  or (_04033_, _04032_, _03980_);
  or (_04034_, _04033_, _03676_);
  and (_04035_, _04034_, _43100_);
  and (_40163_, _04035_, _03979_);
  nand (_04036_, _03676_, _34693_);
  and (_04037_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_04038_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_04039_, _04038_, _04037_);
  and (_04040_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_04041_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_04042_, _04041_, _04040_);
  or (_04043_, _04042_, _04039_);
  and (_04044_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_04045_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_04046_, _04045_, _04044_);
  and (_04047_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_04048_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_04049_, _04048_, _04047_);
  or (_04050_, _04049_, _04046_);
  or (_04051_, _04050_, _04043_);
  and (_04052_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_04053_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or (_04054_, _04053_, _04052_);
  and (_04055_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_04056_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_04058_, _04056_, _04055_);
  or (_04059_, _04058_, _04054_);
  and (_04060_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_04061_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_04062_, _04061_, _04060_);
  and (_04063_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_04064_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_04065_, _04064_, _04063_);
  or (_04066_, _04065_, _04062_);
  or (_04067_, _04066_, _04059_);
  or (_04068_, _04067_, _04051_);
  and (_04069_, _03740_, _42563_);
  and (_04070_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_04071_, _04070_, _04069_);
  and (_04072_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_04073_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_04074_, _04073_, _04072_);
  or (_04075_, _04074_, _04071_);
  and (_04076_, _03749_, _03317_);
  and (_04077_, _03751_, _03527_);
  or (_04078_, _04077_, _04076_);
  and (_04079_, _03756_, _03600_);
  and (_04080_, _03754_, _03466_);
  or (_04081_, _04080_, _04079_);
  or (_04082_, _04081_, _04078_);
  or (_04083_, _04082_, _04075_);
  and (_04084_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_04085_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_04086_, _04085_, _04084_);
  or (_04087_, _04086_, _04083_);
  or (_04088_, _04087_, _04068_);
  and (_04089_, _04088_, _03673_);
  and (_04090_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_04091_, _04090_, _03676_);
  or (_04092_, _04091_, _04089_);
  and (_04093_, _04092_, _43100_);
  and (_40164_, _04093_, _04036_);
  nand (_04094_, _03676_, _35520_);
  and (_04095_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_04096_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_04097_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_04098_, _04097_, _04096_);
  and (_04099_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_04100_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_04101_, _04100_, _04099_);
  or (_04102_, _04101_, _04098_);
  and (_04103_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04104_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_04105_, _04104_, _04103_);
  and (_04106_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_04107_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_04108_, _04107_, _04106_);
  or (_04109_, _04108_, _04105_);
  or (_04110_, _04109_, _04102_);
  and (_04111_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_04112_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_04113_, _04112_, _04111_);
  and (_04114_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_04115_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_04116_, _04115_, _04114_);
  or (_04117_, _04116_, _04113_);
  and (_04118_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_04119_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_04120_, _04119_, _04118_);
  and (_04121_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_04122_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_04123_, _04122_, _04121_);
  or (_04124_, _04123_, _04120_);
  or (_04125_, _04124_, _04117_);
  or (_04126_, _04125_, _04110_);
  and (_04127_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_04128_, _38744_);
  and (_04129_, _03740_, _04128_);
  or (_04130_, _04129_, _04127_);
  and (_04131_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_04132_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_04133_, _04132_, _04131_);
  or (_04134_, _04133_, _04130_);
  and (_04135_, _03749_, _03297_);
  and (_04136_, _03751_, _03548_);
  or (_04137_, _04136_, _04135_);
  and (_04138_, _03756_, _03580_);
  and (_04139_, _03754_, _03446_);
  or (_04140_, _04139_, _04138_);
  or (_04141_, _04140_, _04137_);
  or (_04142_, _04141_, _04134_);
  and (_04143_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_04144_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_04145_, _04144_, _04143_);
  or (_04146_, _04145_, _04142_);
  or (_04147_, _04146_, _04126_);
  and (_04148_, _04147_, _03673_);
  or (_04149_, _04148_, _04095_);
  or (_04150_, _04149_, _03676_);
  and (_04151_, _04150_, _43100_);
  and (_40165_, _04151_, _04094_);
  nand (_04152_, _03676_, _36239_);
  and (_04153_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_04154_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_04155_, _04154_, _04153_);
  and (_04157_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_04158_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_04159_, _04158_, _04157_);
  or (_04160_, _04159_, _04155_);
  and (_04161_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_04162_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_04163_, _04162_, _04161_);
  and (_04164_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_04165_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_04166_, _04165_, _04164_);
  or (_04167_, _04166_, _04163_);
  or (_04168_, _04167_, _04160_);
  and (_04169_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_04170_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_04171_, _04170_, _04169_);
  and (_04172_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_04173_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_04174_, _04173_, _04172_);
  or (_04175_, _04174_, _04171_);
  and (_04176_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_04177_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or (_04178_, _04177_, _04176_);
  and (_04179_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_04180_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_04181_, _04180_, _04179_);
  or (_04182_, _04181_, _04178_);
  or (_04183_, _04182_, _04175_);
  or (_04184_, _04183_, _04168_);
  and (_04185_, _03740_, _42724_);
  and (_04186_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_04187_, _04186_, _04185_);
  and (_04188_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_04189_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_04190_, _04189_, _04188_);
  or (_04191_, _04190_, _04187_);
  and (_04192_, _03749_, _03311_);
  and (_04193_, _03751_, _03534_);
  or (_04194_, _04193_, _04192_);
  and (_04195_, _03756_, _03594_);
  and (_04196_, _03754_, _03460_);
  or (_04197_, _04196_, _04195_);
  or (_04198_, _04197_, _04194_);
  or (_04199_, _04198_, _04191_);
  and (_04200_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_04201_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_04202_, _04201_, _04200_);
  or (_04203_, _04202_, _04199_);
  or (_04204_, _04203_, _04184_);
  and (_04205_, _04204_, _03673_);
  and (_04206_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or (_04207_, _04206_, _03676_);
  or (_04208_, _04207_, _04205_);
  and (_04209_, _04208_, _43100_);
  and (_40166_, _04209_, _04152_);
  and (_40237_, _42861_, _43100_);
  nor (_40241_, _42823_, rst);
  and (_40262_, _43005_, _43100_);
  nor (_40265_, _42701_, rst);
  nor (_40266_, _42617_, rst);
  not (_04210_, _00394_);
  nor (_04211_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_04212_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04213_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _04212_);
  nor (_04214_, _04213_, _04211_);
  nor (_04215_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04216_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _04212_);
  nor (_04217_, _04216_, _04215_);
  not (_04218_, _04217_);
  nor (_04219_, _04218_, _04214_);
  and (_04220_, _04217_, _04214_);
  nor (_04221_, _02220_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04222_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _04212_);
  nor (_04223_, _04222_, _04221_);
  and (_04224_, _04223_, _04220_);
  nor (_04225_, _04223_, _04220_);
  nor (_04226_, _04225_, _04224_);
  not (_04227_, _04226_);
  nor (_04228_, _02239_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04229_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _04212_);
  nor (_04230_, _04229_, _04228_);
  and (_04231_, _04230_, _04224_);
  nor (_04232_, _04230_, _04224_);
  nor (_04233_, _04232_, _04231_);
  and (_04234_, _04233_, _04227_);
  and (_04235_, _04234_, _04219_);
  and (_04236_, _04235_, _04210_);
  not (_04237_, _00312_);
  nor (_04238_, _04217_, _04214_);
  and (_04239_, _04238_, _04234_);
  and (_04240_, _04239_, _04237_);
  or (_04241_, _04240_, _04236_);
  not (_04242_, _00353_);
  and (_04243_, _04218_, _04214_);
  and (_04244_, _04243_, _04234_);
  and (_04245_, _04244_, _04242_);
  not (_04246_, _00035_);
  nor (_04247_, _04233_, _04226_);
  and (_04248_, _04247_, _04219_);
  and (_04249_, _04248_, _04246_);
  or (_04251_, _04249_, _04245_);
  or (_04252_, _04251_, _04241_);
  not (_04253_, _43980_);
  and (_04254_, _04247_, _04238_);
  and (_04255_, _04254_, _04253_);
  not (_04256_, _44021_);
  and (_04257_, _04247_, _04243_);
  and (_04258_, _04257_, _04256_);
  or (_04259_, _04258_, _04255_);
  not (_04260_, _00476_);
  and (_04261_, _04230_, _04226_);
  and (_04262_, _04261_, _04238_);
  and (_04263_, _04262_, _04260_);
  not (_04264_, _00230_);
  not (_04265_, _04230_);
  and (_04266_, _04265_, _04226_);
  and (_04267_, _04266_, _04219_);
  and (_04268_, _04267_, _04264_);
  or (_04269_, _04268_, _04263_);
  not (_04270_, _00517_);
  and (_04271_, _04261_, _04243_);
  and (_04272_, _04271_, _04270_);
  not (_04273_, _00117_);
  and (_04274_, _04266_, _04238_);
  and (_04275_, _04274_, _04273_);
  or (_04276_, _04275_, _04272_);
  or (_04277_, _04276_, _04269_);
  not (_04278_, _00076_);
  and (_04279_, _04232_, _04220_);
  and (_04280_, _04279_, _04278_);
  not (_04281_, _00271_);
  and (_04282_, _04265_, _04224_);
  and (_04283_, _04282_, _04281_);
  and (_04284_, _04223_, _04219_);
  and (_04285_, _04284_, _04230_);
  and (_04286_, _04285_, _00567_);
  not (_04287_, _43939_);
  and (_04288_, _04231_, _04287_);
  or (_04289_, _04288_, _04286_);
  or (_04290_, _04289_, _04283_);
  or (_04291_, _04290_, _04280_);
  not (_04292_, _00435_);
  and (_04293_, _04261_, _04220_);
  and (_04294_, _04293_, _04292_);
  not (_04295_, _00189_);
  and (_04296_, _04266_, _04243_);
  and (_04297_, _04296_, _04295_);
  or (_04298_, _04297_, _04294_);
  or (_04299_, _04298_, _04291_);
  or (_04300_, _04299_, _04277_);
  or (_04301_, _04300_, _04259_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _04301_, _04252_);
  and (_04302_, _04235_, _04292_);
  and (_04303_, _04239_, _04242_);
  or (_04304_, _04303_, _04302_);
  and (_04305_, _04244_, _04210_);
  and (_04306_, _04248_, _04278_);
  or (_04307_, _04306_, _04305_);
  or (_04308_, _04307_, _04304_);
  and (_04309_, _04296_, _04264_);
  and (_04310_, _04274_, _04295_);
  or (_04311_, _04310_, _04309_);
  and (_04312_, _04262_, _04270_);
  and (_04313_, _04267_, _04281_);
  or (_04314_, _04313_, _04312_);
  or (_04315_, _04314_, _04311_);
  and (_04316_, _04279_, _04273_);
  and (_04317_, _04231_, _04253_);
  and (_04318_, _04282_, _04237_);
  and (_04319_, _04285_, _04287_);
  or (_04320_, _04319_, _04318_);
  or (_04321_, _04320_, _04317_);
  or (_04322_, _04321_, _04316_);
  and (_04323_, _04271_, _00567_);
  and (_04324_, _04293_, _04260_);
  or (_04325_, _04324_, _04323_);
  or (_04326_, _04325_, _04322_);
  or (_04327_, _04326_, _04315_);
  and (_04328_, _04257_, _04246_);
  and (_04329_, _04254_, _04256_);
  or (_04330_, _04329_, _04328_);
  or (_04331_, _04330_, _04327_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _04331_, _04308_);
  and (_04332_, _04239_, _04210_);
  and (_04333_, _04248_, _04273_);
  or (_04334_, _04333_, _04332_);
  and (_04335_, _04244_, _04292_);
  and (_04336_, _04235_, _04260_);
  or (_04337_, _04336_, _04335_);
  or (_04338_, _04337_, _04334_);
  and (_04339_, _04254_, _04246_);
  and (_04340_, _04257_, _04278_);
  or (_04341_, _04340_, _04339_);
  and (_04342_, _04262_, _00567_);
  and (_04343_, _04267_, _04237_);
  or (_04344_, _04343_, _04342_);
  and (_04345_, _04293_, _04270_);
  and (_04346_, _04274_, _04264_);
  or (_04347_, _04346_, _04345_);
  or (_04348_, _04347_, _04344_);
  and (_04350_, _04279_, _04295_);
  and (_04351_, _04285_, _04253_);
  and (_04352_, _04282_, _04242_);
  and (_04353_, _04231_, _04256_);
  or (_04354_, _04353_, _04352_);
  or (_04355_, _04354_, _04351_);
  or (_04356_, _04355_, _04350_);
  and (_04357_, _04296_, _04281_);
  and (_04358_, _04271_, _04287_);
  or (_04359_, _04358_, _04357_);
  or (_04360_, _04359_, _04356_);
  or (_04361_, _04360_, _04348_);
  or (_04362_, _04361_, _04341_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _04362_, _04338_);
  and (_04363_, _04231_, _00567_);
  and (_04364_, _04248_, _04256_);
  and (_04365_, _04254_, _04287_);
  or (_04366_, _04365_, _04364_);
  and (_04367_, _04257_, _04253_);
  and (_04368_, _04267_, _04295_);
  and (_04369_, _04296_, _04273_);
  or (_04370_, _04369_, _04368_);
  and (_04371_, _04274_, _04278_);
  and (_04372_, _04279_, _04246_);
  or (_04373_, _04372_, _04371_);
  or (_04374_, _04373_, _04370_);
  or (_04375_, _04374_, _04367_);
  or (_04376_, _04375_, _04366_);
  and (_04377_, _04271_, _04260_);
  and (_04378_, _04285_, _04270_);
  or (_04379_, _04378_, _04377_);
  and (_04380_, _04293_, _04210_);
  and (_04381_, _04262_, _04292_);
  or (_04382_, _04381_, _04380_);
  or (_04383_, _04382_, _04379_);
  and (_04384_, _04235_, _04242_);
  and (_04385_, _04244_, _04237_);
  or (_04386_, _04385_, _04384_);
  and (_04387_, _04239_, _04281_);
  and (_04388_, _04282_, _04264_);
  or (_04389_, _04388_, _04387_);
  or (_04390_, _04389_, _04386_);
  or (_04391_, _04390_, _04383_);
  or (_04392_, _04391_, _04376_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _04392_, _04363_);
  not (_04393_, _00399_);
  and (_04394_, _04239_, _04393_);
  not (_04395_, _00440_);
  and (_04396_, _04244_, _04395_);
  or (_04397_, _04396_, _04394_);
  not (_04398_, _00481_);
  and (_04399_, _04235_, _04398_);
  not (_04400_, _00122_);
  and (_04401_, _04248_, _04400_);
  or (_04402_, _04401_, _04399_);
  or (_04403_, _04402_, _04397_);
  not (_04404_, _00081_);
  and (_04405_, _04257_, _04404_);
  not (_04406_, _00040_);
  and (_04407_, _04254_, _04406_);
  or (_04408_, _04407_, _04405_);
  not (_04409_, _00317_);
  and (_04410_, _04267_, _04409_);
  not (_04411_, _00276_);
  and (_04412_, _04296_, _04411_);
  or (_04413_, _04412_, _04410_);
  not (_04414_, _00235_);
  and (_04415_, _04274_, _04414_);
  not (_04416_, _43944_);
  and (_04417_, _04271_, _04416_);
  or (_04418_, _04417_, _04415_);
  or (_04419_, _04418_, _04413_);
  not (_04420_, _00194_);
  and (_04421_, _04279_, _04420_);
  not (_04422_, _44026_);
  and (_04423_, _04231_, _04422_);
  not (_04424_, _00358_);
  and (_04425_, _04282_, _04424_);
  not (_04426_, _43985_);
  and (_04427_, _04285_, _04426_);
  or (_04428_, _04427_, _04425_);
  or (_04429_, _04428_, _04423_);
  or (_04430_, _04429_, _04421_);
  and (_04431_, _04262_, _00575_);
  not (_04432_, _00522_);
  and (_04433_, _04293_, _04432_);
  or (_04434_, _04433_, _04431_);
  or (_04435_, _04434_, _04430_);
  or (_04436_, _04435_, _04419_);
  or (_04437_, _04436_, _04408_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _04437_, _04403_);
  not (_04438_, _00404_);
  and (_04439_, _04239_, _04438_);
  not (_04440_, _00445_);
  and (_04441_, _04244_, _04440_);
  or (_04442_, _04441_, _04439_);
  not (_04443_, _00486_);
  and (_04444_, _04235_, _04443_);
  not (_04445_, _00127_);
  and (_04446_, _04248_, _04445_);
  or (_04448_, _04446_, _04444_);
  or (_04449_, _04448_, _04442_);
  not (_04450_, _00086_);
  and (_04451_, _04257_, _04450_);
  not (_04452_, _00045_);
  and (_04453_, _04254_, _04452_);
  or (_04454_, _04453_, _04451_);
  not (_04455_, _00322_);
  and (_04456_, _04267_, _04455_);
  not (_04457_, _00281_);
  and (_04458_, _04296_, _04457_);
  or (_04459_, _04458_, _04456_);
  not (_04460_, _00240_);
  and (_04461_, _04274_, _04460_);
  not (_04462_, _43949_);
  and (_04463_, _04271_, _04462_);
  or (_04464_, _04463_, _04461_);
  or (_04465_, _04464_, _04459_);
  not (_04466_, _00199_);
  and (_04467_, _04279_, _04466_);
  not (_04468_, _00004_);
  and (_04469_, _04231_, _04468_);
  not (_04470_, _00363_);
  and (_04471_, _04282_, _04470_);
  not (_04472_, _43990_);
  and (_04473_, _04285_, _04472_);
  or (_04474_, _04473_, _04471_);
  or (_04475_, _04474_, _04469_);
  or (_04476_, _04475_, _04467_);
  and (_04477_, _04262_, _00583_);
  not (_04478_, _00527_);
  and (_04479_, _04293_, _04478_);
  or (_04480_, _04479_, _04477_);
  or (_04481_, _04480_, _04476_);
  or (_04482_, _04481_, _04465_);
  or (_04483_, _04482_, _04454_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _04483_, _04449_);
  not (_04484_, _00409_);
  and (_04485_, _04239_, _04484_);
  not (_04486_, _00450_);
  and (_04487_, _04244_, _04486_);
  or (_04488_, _04487_, _04485_);
  not (_04489_, _00491_);
  and (_04490_, _04235_, _04489_);
  not (_04491_, _00134_);
  and (_04492_, _04248_, _04491_);
  or (_04493_, _04492_, _04490_);
  or (_04494_, _04493_, _04488_);
  not (_04495_, _00091_);
  and (_04496_, _04257_, _04495_);
  not (_04497_, _00050_);
  and (_04498_, _04254_, _04497_);
  or (_04499_, _04498_, _04496_);
  not (_04500_, _00327_);
  and (_04501_, _04267_, _04500_);
  not (_04502_, _00286_);
  and (_04503_, _04296_, _04502_);
  or (_04504_, _04503_, _04501_);
  not (_04505_, _00245_);
  and (_04506_, _04274_, _04505_);
  not (_04507_, _43954_);
  and (_04508_, _04271_, _04507_);
  or (_04509_, _04508_, _04506_);
  or (_04510_, _04509_, _04504_);
  not (_04511_, _00204_);
  and (_04512_, _04279_, _04511_);
  not (_04513_, _00009_);
  and (_04514_, _04231_, _04513_);
  not (_04515_, _00368_);
  and (_04516_, _04282_, _04515_);
  not (_04517_, _43995_);
  and (_04518_, _04285_, _04517_);
  or (_04519_, _04518_, _04516_);
  or (_04520_, _04519_, _04514_);
  or (_04521_, _04520_, _04512_);
  and (_04522_, _04262_, _00591_);
  not (_04523_, _00532_);
  and (_04524_, _04293_, _04523_);
  or (_04525_, _04524_, _04522_);
  or (_04526_, _04525_, _04521_);
  or (_04527_, _04526_, _04510_);
  or (_04528_, _04527_, _04499_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _04528_, _04494_);
  not (_04529_, _00455_);
  and (_04530_, _04244_, _04529_);
  not (_04531_, _00145_);
  and (_04532_, _04248_, _04531_);
  or (_04533_, _04532_, _04530_);
  not (_04534_, _00414_);
  and (_04535_, _04239_, _04534_);
  not (_04536_, _00496_);
  and (_04537_, _04235_, _04536_);
  or (_04538_, _04537_, _04535_);
  or (_04539_, _04538_, _04533_);
  not (_04540_, _00096_);
  and (_04541_, _04257_, _04540_);
  not (_04542_, _00055_);
  and (_04543_, _04254_, _04542_);
  or (_04544_, _04543_, _04541_);
  not (_04545_, _00332_);
  and (_04547_, _04267_, _04545_);
  not (_04548_, _00291_);
  and (_04549_, _04296_, _04548_);
  or (_04550_, _04549_, _04547_);
  not (_04551_, _00537_);
  and (_04552_, _04293_, _04551_);
  not (_04553_, _43959_);
  and (_04554_, _04271_, _04553_);
  or (_04555_, _04554_, _04552_);
  or (_04556_, _04555_, _04550_);
  not (_04557_, _00209_);
  and (_04558_, _04279_, _04557_);
  not (_04559_, _00014_);
  and (_04560_, _04231_, _04559_);
  not (_04561_, _00373_);
  and (_04562_, _04282_, _04561_);
  not (_04563_, _44000_);
  and (_04564_, _04285_, _04563_);
  or (_04565_, _04564_, _04562_);
  or (_04566_, _04565_, _04560_);
  or (_04567_, _04566_, _04558_);
  and (_04568_, _04262_, _00597_);
  not (_04569_, _00250_);
  and (_04570_, _04274_, _04569_);
  or (_04571_, _04570_, _04568_);
  or (_04572_, _04571_, _04567_);
  or (_04573_, _04572_, _04556_);
  or (_04574_, _04573_, _04544_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _04574_, _04539_);
  not (_04575_, _00460_);
  and (_04576_, _04244_, _04575_);
  not (_04577_, _00156_);
  and (_04578_, _04248_, _04577_);
  or (_04579_, _04578_, _04576_);
  not (_04580_, _00419_);
  and (_04581_, _04239_, _04580_);
  not (_04582_, _00501_);
  and (_04583_, _04235_, _04582_);
  or (_04584_, _04583_, _04581_);
  or (_04585_, _04584_, _04579_);
  not (_04586_, _00101_);
  and (_04587_, _04257_, _04586_);
  not (_04588_, _00060_);
  and (_04589_, _04254_, _04588_);
  or (_04590_, _04589_, _04587_);
  not (_04591_, _00337_);
  and (_04592_, _04267_, _04591_);
  not (_04593_, _00296_);
  and (_04594_, _04296_, _04593_);
  or (_04595_, _04594_, _04592_);
  not (_04596_, _00542_);
  and (_04597_, _04293_, _04596_);
  not (_04598_, _43964_);
  and (_04599_, _04271_, _04598_);
  or (_04600_, _04599_, _04597_);
  or (_04601_, _04600_, _04595_);
  not (_04602_, _00214_);
  and (_04603_, _04279_, _04602_);
  not (_04604_, _00378_);
  and (_04605_, _04282_, _04604_);
  not (_04606_, _44005_);
  and (_04607_, _04285_, _04606_);
  not (_04608_, _00019_);
  and (_04609_, _04231_, _04608_);
  or (_04610_, _04609_, _04607_);
  or (_04611_, _04610_, _04605_);
  or (_04612_, _04611_, _04603_);
  and (_04613_, _04262_, _00602_);
  not (_04614_, _00255_);
  and (_04615_, _04274_, _04614_);
  or (_04616_, _04615_, _04613_);
  or (_04617_, _04616_, _04612_);
  or (_04618_, _04617_, _04601_);
  or (_04619_, _04618_, _04590_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _04619_, _04585_);
  not (_04620_, _00424_);
  and (_04621_, _04239_, _04620_);
  not (_04622_, _00465_);
  and (_04623_, _04244_, _04622_);
  or (_04624_, _04623_, _04621_);
  not (_04625_, _00506_);
  and (_04626_, _04235_, _04625_);
  not (_04627_, _00167_);
  and (_04628_, _04248_, _04627_);
  or (_04629_, _04628_, _04626_);
  or (_04630_, _04629_, _04624_);
  not (_04631_, _00106_);
  and (_04632_, _04257_, _04631_);
  not (_04633_, _00065_);
  and (_04634_, _04254_, _04633_);
  or (_04635_, _04634_, _04632_);
  not (_04636_, _00342_);
  and (_04637_, _04267_, _04636_);
  not (_04638_, _00301_);
  and (_04639_, _04296_, _04638_);
  or (_04640_, _04639_, _04637_);
  not (_04641_, _00260_);
  and (_04642_, _04274_, _04641_);
  not (_04643_, _43969_);
  and (_04644_, _04271_, _04643_);
  or (_04646_, _04644_, _04642_);
  or (_04647_, _04646_, _04640_);
  not (_04648_, _00219_);
  and (_04649_, _04279_, _04648_);
  not (_04650_, _00024_);
  and (_04651_, _04231_, _04650_);
  not (_04652_, _00383_);
  and (_04653_, _04282_, _04652_);
  not (_04654_, _44010_);
  and (_04655_, _04285_, _04654_);
  or (_04656_, _04655_, _04653_);
  or (_04657_, _04656_, _04651_);
  or (_04658_, _04657_, _04649_);
  and (_04659_, _04262_, _00607_);
  not (_04660_, _00550_);
  and (_04661_, _04293_, _04660_);
  or (_04662_, _04661_, _04659_);
  or (_04663_, _04662_, _04658_);
  or (_04664_, _04663_, _04647_);
  or (_04665_, _04664_, _04635_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _04665_, _04630_);
  not (_04666_, _00429_);
  and (_04667_, _04239_, _04666_);
  not (_04668_, _00470_);
  and (_04669_, _04244_, _04668_);
  or (_04670_, _04669_, _04667_);
  not (_04671_, _00511_);
  and (_04672_, _04235_, _04671_);
  not (_04673_, _00178_);
  and (_04674_, _04248_, _04673_);
  or (_04675_, _04674_, _04672_);
  or (_04676_, _04675_, _04670_);
  not (_04677_, _00111_);
  and (_04678_, _04257_, _04677_);
  not (_04679_, _00070_);
  and (_04680_, _04254_, _04679_);
  or (_04681_, _04680_, _04678_);
  not (_04682_, _00347_);
  and (_04683_, _04267_, _04682_);
  not (_04684_, _00306_);
  and (_04685_, _04296_, _04684_);
  or (_04686_, _04685_, _04683_);
  not (_04687_, _00265_);
  and (_04688_, _04274_, _04687_);
  not (_04689_, _43974_);
  and (_04690_, _04271_, _04689_);
  or (_04691_, _04690_, _04688_);
  or (_04692_, _04691_, _04686_);
  not (_04693_, _00224_);
  and (_04694_, _04279_, _04693_);
  not (_04695_, _00029_);
  and (_04696_, _04231_, _04695_);
  not (_04697_, _00388_);
  and (_04698_, _04282_, _04697_);
  not (_04699_, _44015_);
  and (_04700_, _04285_, _04699_);
  or (_04701_, _04700_, _04698_);
  or (_04702_, _04701_, _04696_);
  or (_04703_, _04702_, _04694_);
  and (_04704_, _04262_, _00612_);
  not (_04705_, _00558_);
  and (_04706_, _04293_, _04705_);
  or (_04707_, _04706_, _04704_);
  or (_04708_, _04707_, _04703_);
  or (_04709_, _04708_, _04692_);
  or (_04710_, _04709_, _04681_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _04710_, _04676_);
  and (_04711_, _04235_, _04395_);
  and (_04712_, _04244_, _04393_);
  or (_04713_, _04712_, _04711_);
  and (_04714_, _04239_, _04424_);
  and (_04715_, _04248_, _04404_);
  or (_04716_, _04715_, _04714_);
  or (_04717_, _04716_, _04713_);
  and (_04718_, _04296_, _04414_);
  and (_04719_, _04274_, _04420_);
  or (_04720_, _04719_, _04718_);
  and (_04721_, _04262_, _04432_);
  and (_04722_, _04267_, _04411_);
  or (_04723_, _04722_, _04721_);
  or (_04724_, _04723_, _04720_);
  and (_04725_, _04279_, _04400_);
  and (_04726_, _04231_, _04426_);
  and (_04727_, _04282_, _04409_);
  and (_04728_, _04285_, _04416_);
  or (_04729_, _04728_, _04727_);
  or (_04730_, _04729_, _04726_);
  or (_04731_, _04730_, _04725_);
  and (_04732_, _04271_, _00575_);
  and (_04733_, _04293_, _04398_);
  or (_04734_, _04733_, _04732_);
  or (_04735_, _04734_, _04731_);
  or (_04736_, _04735_, _04724_);
  and (_04737_, _04257_, _04406_);
  and (_04738_, _04254_, _04422_);
  or (_04739_, _04738_, _04737_);
  or (_04740_, _04739_, _04736_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _04740_, _04717_);
  and (_04741_, _04244_, _04438_);
  and (_04742_, _04239_, _04470_);
  or (_04743_, _04742_, _04741_);
  and (_04744_, _04235_, _04440_);
  and (_04745_, _04248_, _04450_);
  or (_04746_, _04745_, _04744_);
  or (_04747_, _04746_, _04743_);
  and (_04748_, _04296_, _04460_);
  and (_04749_, _04274_, _04466_);
  or (_04750_, _04749_, _04748_);
  and (_04751_, _04271_, _00583_);
  and (_04752_, _04262_, _04478_);
  or (_04753_, _04752_, _04751_);
  or (_04754_, _04753_, _04750_);
  and (_04755_, _04279_, _04445_);
  and (_04756_, _04231_, _04472_);
  and (_04757_, _04282_, _04455_);
  and (_04758_, _04285_, _04462_);
  or (_04759_, _04758_, _04757_);
  or (_04760_, _04759_, _04756_);
  or (_04761_, _04760_, _04755_);
  and (_04762_, _04293_, _04443_);
  and (_04763_, _04267_, _04457_);
  or (_04764_, _04763_, _04762_);
  or (_04765_, _04764_, _04761_);
  or (_04766_, _04765_, _04754_);
  and (_04767_, _04257_, _04452_);
  and (_04768_, _04254_, _04468_);
  or (_04769_, _04768_, _04767_);
  or (_04770_, _04769_, _04766_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _04770_, _04747_);
  and (_04771_, _04235_, _04486_);
  and (_04772_, _04244_, _04484_);
  or (_04773_, _04772_, _04771_);
  and (_04774_, _04239_, _04515_);
  and (_04775_, _04248_, _04495_);
  or (_04776_, _04775_, _04774_);
  or (_04777_, _04776_, _04773_);
  and (_04778_, _04296_, _04505_);
  and (_04779_, _04274_, _04511_);
  or (_04780_, _04779_, _04778_);
  and (_04781_, _04262_, _04523_);
  and (_04782_, _04267_, _04502_);
  or (_04783_, _04782_, _04781_);
  or (_04784_, _04783_, _04780_);
  and (_04785_, _04279_, _04491_);
  and (_04786_, _04231_, _04517_);
  and (_04787_, _04282_, _04500_);
  and (_04788_, _04285_, _04507_);
  or (_04789_, _04788_, _04787_);
  or (_04790_, _04789_, _04786_);
  or (_04791_, _04790_, _04785_);
  and (_04792_, _04271_, _00591_);
  and (_04793_, _04293_, _04489_);
  or (_04794_, _04793_, _04792_);
  or (_04795_, _04794_, _04791_);
  or (_04796_, _04795_, _04784_);
  and (_04797_, _04257_, _04497_);
  and (_04798_, _04254_, _04513_);
  or (_04799_, _04798_, _04797_);
  or (_04800_, _04799_, _04796_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _04800_, _04777_);
  and (_04801_, _04244_, _04534_);
  and (_04802_, _04235_, _04529_);
  or (_04803_, _04802_, _04801_);
  and (_04804_, _04239_, _04561_);
  and (_04805_, _04248_, _04540_);
  or (_04806_, _04805_, _04804_);
  or (_04807_, _04806_, _04803_);
  and (_04808_, _04271_, _00597_);
  and (_04809_, _04267_, _04548_);
  or (_04810_, _04809_, _04808_);
  and (_04811_, _04293_, _04536_);
  and (_04812_, _04274_, _04557_);
  or (_04813_, _04812_, _04811_);
  or (_04814_, _04813_, _04810_);
  and (_04815_, _04279_, _04531_);
  and (_04816_, _04282_, _04545_);
  and (_04817_, _04285_, _04553_);
  and (_04818_, _04231_, _04563_);
  or (_04819_, _04818_, _04817_);
  or (_04820_, _04819_, _04816_);
  or (_04821_, _04820_, _04815_);
  and (_04822_, _04262_, _04551_);
  and (_04823_, _04296_, _04569_);
  or (_04824_, _04823_, _04822_);
  or (_04825_, _04824_, _04821_);
  or (_04826_, _04825_, _04814_);
  and (_04827_, _04257_, _04542_);
  and (_04828_, _04254_, _04559_);
  or (_04829_, _04828_, _04827_);
  or (_04830_, _04829_, _04826_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _04830_, _04807_);
  and (_04831_, _04235_, _04575_);
  and (_04832_, _04239_, _04604_);
  or (_04833_, _04832_, _04831_);
  and (_04834_, _04244_, _04580_);
  and (_04835_, _04248_, _04586_);
  or (_04836_, _04835_, _04834_);
  or (_04837_, _04836_, _04833_);
  and (_04838_, _04296_, _04614_);
  and (_04839_, _04274_, _04602_);
  or (_04840_, _04839_, _04838_);
  and (_04841_, _04262_, _04596_);
  and (_04842_, _04267_, _04593_);
  or (_04843_, _04842_, _04841_);
  or (_04844_, _04843_, _04840_);
  and (_04845_, _04279_, _04577_);
  and (_04846_, _04231_, _04606_);
  and (_04847_, _04282_, _04591_);
  and (_04848_, _04285_, _04598_);
  or (_04849_, _04848_, _04847_);
  or (_04850_, _04849_, _04846_);
  or (_04851_, _04850_, _04845_);
  and (_04852_, _04271_, _00602_);
  and (_04853_, _04293_, _04582_);
  or (_04854_, _04853_, _04852_);
  or (_04855_, _04854_, _04851_);
  or (_04856_, _04855_, _04844_);
  and (_04857_, _04257_, _04588_);
  and (_04858_, _04254_, _04608_);
  or (_04859_, _04858_, _04857_);
  or (_04860_, _04859_, _04856_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _04860_, _04837_);
  and (_04861_, _04244_, _04620_);
  and (_04862_, _04235_, _04622_);
  or (_04863_, _04862_, _04861_);
  and (_04864_, _04239_, _04652_);
  and (_04865_, _04248_, _04631_);
  or (_04866_, _04865_, _04864_);
  or (_04867_, _04866_, _04863_);
  and (_04868_, _04296_, _04641_);
  and (_04869_, _04274_, _04648_);
  or (_04870_, _04869_, _04868_);
  and (_04871_, _04271_, _00607_);
  and (_04872_, _04293_, _04625_);
  or (_04873_, _04872_, _04871_);
  or (_04874_, _04873_, _04870_);
  and (_04875_, _04279_, _04627_);
  and (_04876_, _04285_, _04643_);
  and (_04877_, _04282_, _04636_);
  and (_04878_, _04231_, _04654_);
  or (_04879_, _04878_, _04877_);
  or (_04880_, _04879_, _04876_);
  or (_04881_, _04880_, _04875_);
  and (_04882_, _04262_, _04660_);
  and (_04883_, _04267_, _04638_);
  or (_04884_, _04883_, _04882_);
  or (_04885_, _04884_, _04881_);
  or (_04886_, _04885_, _04874_);
  and (_04887_, _04257_, _04633_);
  and (_04888_, _04254_, _04650_);
  or (_04889_, _04888_, _04887_);
  or (_04890_, _04889_, _04886_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _04890_, _04867_);
  and (_04891_, _04235_, _04668_);
  and (_04892_, _04239_, _04697_);
  or (_04893_, _04892_, _04891_);
  and (_04894_, _04244_, _04666_);
  and (_04895_, _04248_, _04677_);
  or (_04896_, _04895_, _04894_);
  or (_04897_, _04896_, _04893_);
  and (_04898_, _04296_, _04687_);
  and (_04899_, _04274_, _04693_);
  or (_04900_, _04899_, _04898_);
  and (_04901_, _04262_, _04705_);
  and (_04902_, _04267_, _04684_);
  or (_04903_, _04902_, _04901_);
  or (_04904_, _04903_, _04900_);
  and (_04905_, _04279_, _04673_);
  and (_04906_, _04231_, _04699_);
  and (_04907_, _04282_, _04682_);
  and (_04908_, _04285_, _04689_);
  or (_04909_, _04908_, _04907_);
  or (_04910_, _04909_, _04906_);
  or (_04911_, _04910_, _04905_);
  and (_04912_, _04271_, _00612_);
  and (_04913_, _04293_, _04671_);
  or (_04914_, _04913_, _04912_);
  or (_04915_, _04914_, _04911_);
  or (_04916_, _04915_, _04904_);
  and (_04917_, _04257_, _04679_);
  and (_04918_, _04254_, _04695_);
  or (_04919_, _04918_, _04917_);
  or (_04920_, _04919_, _04916_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _04920_, _04897_);
  and (_04921_, _04235_, _04393_);
  and (_04922_, _04239_, _04409_);
  or (_04923_, _04922_, _04921_);
  and (_04924_, _04244_, _04424_);
  and (_04925_, _04248_, _04406_);
  or (_04926_, _04925_, _04924_);
  or (_04927_, _04926_, _04923_);
  and (_04928_, _04254_, _04426_);
  and (_04929_, _04257_, _04422_);
  or (_04930_, _04929_, _04928_);
  and (_04931_, _04274_, _04400_);
  and (_04932_, _04296_, _04420_);
  or (_04933_, _04932_, _04931_);
  and (_04934_, _04262_, _04398_);
  and (_04935_, _04267_, _04414_);
  or (_04936_, _04935_, _04934_);
  or (_04937_, _04936_, _04933_);
  and (_04938_, _04279_, _04404_);
  and (_04939_, _04231_, _04416_);
  and (_04940_, _04285_, _00575_);
  and (_04941_, _04282_, _04411_);
  or (_04942_, _04941_, _04940_);
  or (_04943_, _04942_, _04939_);
  or (_04944_, _04943_, _04938_);
  and (_04945_, _04271_, _04432_);
  and (_04946_, _04293_, _04395_);
  or (_04947_, _04946_, _04945_);
  or (_04948_, _04947_, _04944_);
  or (_04949_, _04948_, _04937_);
  or (_04950_, _04949_, _04930_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _04950_, _04927_);
  and (_04951_, _04239_, _04455_);
  and (_04952_, _04244_, _04470_);
  or (_04953_, _04952_, _04951_);
  and (_04954_, _04235_, _04438_);
  and (_04955_, _04248_, _04452_);
  or (_04956_, _04955_, _04954_);
  or (_04957_, _04956_, _04953_);
  and (_04958_, _04254_, _04472_);
  and (_04959_, _04257_, _04468_);
  or (_04960_, _04959_, _04958_);
  and (_04961_, _04262_, _04443_);
  and (_04962_, _04271_, _04478_);
  or (_04963_, _04962_, _04961_);
  and (_04964_, _04274_, _04445_);
  and (_04965_, _04296_, _04466_);
  or (_04966_, _04965_, _04964_);
  or (_04967_, _04966_, _04963_);
  and (_04968_, _04279_, _04450_);
  and (_04969_, _04285_, _00583_);
  and (_04970_, _04282_, _04457_);
  and (_04971_, _04231_, _04462_);
  or (_04972_, _04971_, _04970_);
  or (_04973_, _04972_, _04969_);
  or (_04974_, _04973_, _04968_);
  and (_04975_, _04293_, _04440_);
  and (_04976_, _04267_, _04460_);
  or (_04977_, _04976_, _04975_);
  or (_04978_, _04977_, _04974_);
  or (_04979_, _04978_, _04967_);
  or (_04980_, _04979_, _04960_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _04980_, _04957_);
  and (_04981_, _04244_, _04515_);
  and (_04982_, _04239_, _04500_);
  or (_04983_, _04982_, _04981_);
  and (_04984_, _04235_, _04484_);
  and (_04985_, _04248_, _04497_);
  or (_04986_, _04985_, _04984_);
  or (_04987_, _04986_, _04983_);
  and (_04988_, _04254_, _04517_);
  and (_04989_, _04257_, _04513_);
  or (_04990_, _04989_, _04988_);
  and (_04991_, _04267_, _04505_);
  and (_04992_, _04274_, _04491_);
  or (_04993_, _04992_, _04991_);
  and (_04994_, _04293_, _04486_);
  and (_04995_, _04296_, _04511_);
  or (_04996_, _04995_, _04994_);
  or (_04997_, _04996_, _04993_);
  and (_04998_, _04271_, _04523_);
  and (_04999_, _04262_, _04489_);
  or (_05000_, _04999_, _04998_);
  and (_05001_, _04279_, _04495_);
  and (_05002_, _04231_, _04507_);
  and (_05003_, _04285_, _00591_);
  and (_05004_, _04282_, _04502_);
  or (_05005_, _05004_, _05003_);
  or (_05006_, _05005_, _05002_);
  or (_05007_, _05006_, _05001_);
  or (_05008_, _05007_, _05000_);
  or (_05009_, _05008_, _04997_);
  or (_05010_, _05009_, _04990_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _05010_, _04987_);
  and (_05011_, _04239_, _04545_);
  and (_05012_, _04244_, _04561_);
  or (_05013_, _05012_, _05011_);
  and (_05014_, _04235_, _04534_);
  and (_05015_, _04248_, _04542_);
  or (_05016_, _05015_, _05014_);
  or (_05017_, _05016_, _05013_);
  and (_05018_, _04254_, _04563_);
  and (_05019_, _04257_, _04559_);
  or (_05020_, _05019_, _05018_);
  and (_05021_, _04262_, _04536_);
  and (_05022_, _04271_, _04551_);
  or (_05023_, _05022_, _05021_);
  and (_05024_, _04274_, _04531_);
  and (_05025_, _04296_, _04557_);
  or (_05026_, _05025_, _05024_);
  or (_05027_, _05026_, _05023_);
  and (_05028_, _04279_, _04540_);
  and (_05029_, _04285_, _00597_);
  and (_05030_, _04282_, _04548_);
  and (_05031_, _04231_, _04553_);
  or (_05032_, _05031_, _05030_);
  or (_05033_, _05032_, _05029_);
  or (_05034_, _05033_, _05028_);
  and (_05035_, _04293_, _04529_);
  and (_05036_, _04267_, _04569_);
  or (_05037_, _05036_, _05035_);
  or (_05038_, _05037_, _05034_);
  or (_05039_, _05038_, _05027_);
  or (_05040_, _05039_, _05020_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _05040_, _05017_);
  and (_05041_, _04235_, _04580_);
  and (_05042_, _04239_, _04591_);
  or (_05043_, _05042_, _05041_);
  and (_05044_, _04244_, _04604_);
  and (_05045_, _04248_, _04588_);
  or (_05046_, _05045_, _05044_);
  or (_05047_, _05046_, _05043_);
  and (_05048_, _04254_, _04606_);
  and (_05049_, _04257_, _04608_);
  or (_05050_, _05049_, _05048_);
  and (_05051_, _04274_, _04577_);
  and (_05052_, _04296_, _04602_);
  or (_05053_, _05052_, _05051_);
  and (_05054_, _04262_, _04582_);
  and (_05055_, _04267_, _04614_);
  or (_05056_, _05055_, _05054_);
  or (_05057_, _05056_, _05053_);
  and (_05058_, _04279_, _04586_);
  and (_05059_, _04231_, _04598_);
  and (_05060_, _04285_, _00602_);
  and (_05061_, _04282_, _04593_);
  or (_05062_, _05061_, _05060_);
  or (_05063_, _05062_, _05059_);
  or (_05064_, _05063_, _05058_);
  and (_05065_, _04271_, _04596_);
  and (_05066_, _04293_, _04575_);
  or (_05067_, _05066_, _05065_);
  or (_05068_, _05067_, _05064_);
  or (_05069_, _05068_, _05057_);
  or (_05070_, _05069_, _05050_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _05070_, _05047_);
  and (_05071_, _04235_, _04620_);
  and (_05072_, _04244_, _04652_);
  or (_05073_, _05072_, _05071_);
  and (_05074_, _04239_, _04636_);
  and (_05075_, _04248_, _04633_);
  or (_05076_, _05075_, _05074_);
  or (_05077_, _05076_, _05073_);
  and (_05078_, _04254_, _04654_);
  and (_05079_, _04257_, _04650_);
  or (_05080_, _05079_, _05078_);
  and (_05081_, _04274_, _04627_);
  and (_05082_, _04296_, _04648_);
  or (_05083_, _05082_, _05081_);
  and (_05084_, _04262_, _04625_);
  and (_05086_, _04267_, _04641_);
  or (_05088_, _05086_, _05084_);
  or (_05090_, _05088_, _05083_);
  and (_05092_, _04279_, _04631_);
  and (_05094_, _04231_, _04643_);
  and (_05096_, _04285_, _00607_);
  and (_05098_, _04282_, _04638_);
  or (_05099_, _05098_, _05096_);
  or (_05100_, _05099_, _05094_);
  or (_05101_, _05100_, _05092_);
  and (_05102_, _04271_, _04660_);
  and (_05103_, _04293_, _04622_);
  or (_05104_, _05103_, _05102_);
  or (_05106_, _05104_, _05101_);
  or (_05107_, _05106_, _05090_);
  or (_05109_, _05107_, _05080_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _05109_, _05077_);
  and (_05110_, _04235_, _04666_);
  and (_05112_, _04244_, _04697_);
  or (_05113_, _05112_, _05110_);
  and (_05114_, _04239_, _04682_);
  and (_05116_, _04248_, _04679_);
  or (_05117_, _05116_, _05114_);
  or (_05118_, _05117_, _05113_);
  and (_05120_, _04254_, _04699_);
  and (_05121_, _04257_, _04695_);
  or (_05122_, _05121_, _05120_);
  and (_05124_, _04274_, _04673_);
  and (_05125_, _04296_, _04693_);
  or (_05126_, _05125_, _05124_);
  and (_05128_, _04262_, _04671_);
  and (_05129_, _04267_, _04687_);
  or (_05130_, _05129_, _05128_);
  or (_05132_, _05130_, _05126_);
  and (_05133_, _04279_, _04677_);
  and (_05134_, _04231_, _04689_);
  and (_05136_, _04285_, _00612_);
  and (_05137_, _04282_, _04684_);
  or (_05138_, _05137_, _05136_);
  or (_05139_, _05138_, _05134_);
  or (_05140_, _05139_, _05133_);
  and (_05141_, _04271_, _04705_);
  and (_05142_, _04293_, _04668_);
  or (_05143_, _05142_, _05141_);
  or (_05144_, _05143_, _05140_);
  or (_05145_, _05144_, _05132_);
  or (_05146_, _05145_, _05122_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _05146_, _05118_);
  and (_05147_, _04244_, _04409_);
  and (_05148_, _04235_, _04424_);
  or (_05149_, _05148_, _05147_);
  and (_05150_, _04239_, _04411_);
  and (_05151_, _04248_, _04422_);
  or (_05152_, _05151_, _05150_);
  or (_05153_, _05152_, _05149_);
  and (_05154_, _04271_, _04398_);
  and (_05155_, _04274_, _04404_);
  or (_05157_, _05155_, _05154_);
  and (_05158_, _04293_, _04393_);
  and (_05160_, _04267_, _04420_);
  or (_05161_, _05160_, _05158_);
  or (_05162_, _05161_, _05157_);
  and (_05164_, _04279_, _04406_);
  and (_05165_, _04231_, _00575_);
  and (_05166_, _04285_, _04432_);
  and (_05168_, _04282_, _04414_);
  or (_05169_, _05168_, _05166_);
  or (_05170_, _05169_, _05165_);
  or (_05172_, _05170_, _05164_);
  and (_05173_, _04262_, _04395_);
  and (_05174_, _04296_, _04400_);
  or (_05176_, _05174_, _05173_);
  or (_05177_, _05176_, _05172_);
  or (_05178_, _05177_, _05162_);
  and (_05180_, _04254_, _04416_);
  and (_05181_, _04257_, _04426_);
  or (_05182_, _05181_, _05180_);
  or (_05184_, _05182_, _05178_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _05184_, _05153_);
  and (_05185_, _04231_, _00583_);
  and (_05187_, _04248_, _04468_);
  and (_05188_, _04254_, _04462_);
  or (_05189_, _05188_, _05187_);
  and (_05190_, _04257_, _04472_);
  and (_05191_, _04267_, _04466_);
  and (_05192_, _04296_, _04445_);
  or (_05193_, _05192_, _05191_);
  and (_05194_, _04274_, _04450_);
  and (_05195_, _04279_, _04452_);
  or (_05196_, _05195_, _05194_);
  or (_05197_, _05196_, _05193_);
  or (_05198_, _05197_, _05190_);
  or (_05199_, _05198_, _05189_);
  and (_05200_, _04271_, _04443_);
  and (_05201_, _04285_, _04478_);
  or (_05202_, _05201_, _05200_);
  and (_05203_, _04293_, _04438_);
  and (_05204_, _04262_, _04440_);
  or (_05205_, _05204_, _05203_);
  or (_05206_, _05205_, _05202_);
  and (_05207_, _04235_, _04470_);
  and (_05209_, _04244_, _04455_);
  or (_05210_, _05209_, _05207_);
  and (_05212_, _04239_, _04457_);
  and (_05213_, _04282_, _04460_);
  or (_05214_, _05213_, _05212_);
  or (_05216_, _05214_, _05210_);
  or (_05217_, _05216_, _05206_);
  or (_05218_, _05217_, _05199_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _05218_, _05185_);
  and (_05220_, _04244_, _04500_);
  and (_05221_, _04235_, _04515_);
  or (_05223_, _05221_, _05220_);
  and (_05224_, _04239_, _04502_);
  and (_05225_, _04248_, _04513_);
  or (_05227_, _05225_, _05224_);
  or (_05228_, _05227_, _05223_);
  and (_05229_, _04267_, _04511_);
  and (_05231_, _04274_, _04495_);
  or (_05232_, _05231_, _05229_);
  and (_05233_, _04293_, _04484_);
  and (_05235_, _04296_, _04491_);
  or (_05236_, _05235_, _05233_);
  or (_05237_, _05236_, _05232_);
  and (_05239_, _04279_, _04497_);
  and (_05240_, _04231_, _00591_);
  and (_05241_, _04285_, _04523_);
  and (_05242_, _04282_, _04505_);
  or (_05243_, _05242_, _05241_);
  or (_05244_, _05243_, _05240_);
  or (_05245_, _05244_, _05239_);
  and (_05246_, _04271_, _04489_);
  and (_05247_, _04262_, _04486_);
  or (_05248_, _05247_, _05246_);
  or (_05249_, _05248_, _05245_);
  or (_05250_, _05249_, _05237_);
  and (_05251_, _04254_, _04507_);
  and (_05252_, _04257_, _04517_);
  or (_05253_, _05252_, _05251_);
  or (_05254_, _05253_, _05250_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _05254_, _05228_);
  and (_05255_, _04244_, _04545_);
  and (_05256_, _04235_, _04561_);
  or (_05257_, _05256_, _05255_);
  and (_05258_, _04239_, _04548_);
  and (_05260_, _04248_, _04559_);
  or (_05261_, _05260_, _05258_);
  or (_05263_, _05261_, _05257_);
  and (_05264_, _04271_, _04536_);
  and (_05265_, _04274_, _04540_);
  or (_05267_, _05265_, _05264_);
  and (_05268_, _04293_, _04534_);
  and (_05269_, _04267_, _04557_);
  or (_05271_, _05269_, _05268_);
  or (_05272_, _05271_, _05267_);
  and (_05273_, _04279_, _04542_);
  and (_05275_, _04231_, _00597_);
  and (_05276_, _04285_, _04551_);
  and (_05277_, _04282_, _04569_);
  or (_05279_, _05277_, _05276_);
  or (_05280_, _05279_, _05275_);
  or (_05281_, _05280_, _05273_);
  and (_05283_, _04262_, _04529_);
  and (_05284_, _04296_, _04531_);
  or (_05285_, _05284_, _05283_);
  or (_05287_, _05285_, _05281_);
  or (_05288_, _05287_, _05272_);
  and (_05289_, _04254_, _04553_);
  and (_05291_, _04257_, _04563_);
  or (_05292_, _05291_, _05289_);
  or (_05293_, _05292_, _05288_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _05293_, _05263_);
  and (_05294_, _04231_, _00602_);
  and (_05295_, _04248_, _04608_);
  and (_05296_, _04254_, _04598_);
  or (_05297_, _05296_, _05295_);
  and (_05298_, _04257_, _04606_);
  and (_05299_, _04267_, _04602_);
  and (_05300_, _04296_, _04577_);
  or (_05301_, _05300_, _05299_);
  and (_05302_, _04279_, _04588_);
  and (_05303_, _04274_, _04586_);
  or (_05304_, _05303_, _05302_);
  or (_05305_, _05304_, _05301_);
  or (_05306_, _05305_, _05298_);
  or (_05307_, _05306_, _05297_);
  and (_05308_, _04262_, _04575_);
  and (_05309_, _04293_, _04580_);
  or (_05310_, _05309_, _05308_);
  and (_05312_, _04271_, _04582_);
  and (_05313_, _04285_, _04596_);
  or (_05315_, _05313_, _05312_);
  or (_05316_, _05315_, _05310_);
  and (_05317_, _04235_, _04604_);
  and (_05319_, _04244_, _04591_);
  or (_05320_, _05319_, _05317_);
  and (_05321_, _04239_, _04593_);
  and (_05323_, _04282_, _04614_);
  or (_05324_, _05323_, _05321_);
  or (_05325_, _05324_, _05320_);
  or (_05327_, _05325_, _05316_);
  or (_05328_, _05327_, _05307_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _05328_, _05294_);
  and (_05330_, _04235_, _04652_);
  and (_05331_, _04244_, _04636_);
  or (_05332_, _05331_, _05330_);
  and (_05334_, _04239_, _04638_);
  and (_05335_, _04248_, _04650_);
  or (_05336_, _05335_, _05334_);
  or (_05338_, _05336_, _05332_);
  and (_05339_, _04254_, _04643_);
  and (_05340_, _04257_, _04654_);
  or (_05342_, _05340_, _05339_);
  and (_05343_, _04271_, _04625_);
  and (_05344_, _04296_, _04627_);
  or (_05345_, _05344_, _05343_);
  and (_05346_, _04267_, _04648_);
  and (_05347_, _04274_, _04631_);
  or (_05348_, _05347_, _05346_);
  or (_05349_, _05348_, _05345_);
  and (_05350_, _04262_, _04622_);
  and (_05351_, _04293_, _04620_);
  or (_05352_, _05351_, _05350_);
  and (_05353_, _04279_, _04633_);
  and (_05354_, _04282_, _04641_);
  and (_05355_, _04231_, _00607_);
  and (_05356_, _04285_, _04660_);
  or (_05357_, _05356_, _05355_);
  or (_05358_, _05357_, _05354_);
  or (_05359_, _05358_, _05353_);
  or (_05360_, _05359_, _05352_);
  or (_05361_, _05360_, _05349_);
  or (_05362_, _05361_, _05342_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _05362_, _05338_);
  and (_05364_, _04244_, _04682_);
  and (_05366_, _04235_, _04697_);
  or (_05367_, _05366_, _05364_);
  and (_05368_, _04239_, _04684_);
  and (_05370_, _04248_, _04695_);
  or (_05371_, _05370_, _05368_);
  or (_05372_, _05371_, _05367_);
  and (_05374_, _04271_, _04671_);
  and (_05375_, _04274_, _04677_);
  or (_05376_, _05375_, _05374_);
  and (_05378_, _04293_, _04666_);
  and (_05379_, _04267_, _04693_);
  or (_05380_, _05379_, _05378_);
  or (_05382_, _05380_, _05376_);
  and (_05383_, _04279_, _04679_);
  and (_05384_, _04231_, _00612_);
  and (_05386_, _04285_, _04705_);
  and (_05387_, _04282_, _04687_);
  or (_05388_, _05387_, _05386_);
  or (_05390_, _05388_, _05384_);
  or (_05391_, _05390_, _05383_);
  and (_05392_, _04262_, _04668_);
  and (_05394_, _04296_, _04673_);
  or (_05395_, _05394_, _05392_);
  or (_05396_, _05395_, _05391_);
  or (_05397_, _05396_, _05382_);
  and (_05398_, _04254_, _04689_);
  and (_05399_, _04257_, _04699_);
  or (_05400_, _05399_, _05398_);
  or (_05401_, _05400_, _05397_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _05401_, _05372_);
  nand (_05402_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_05403_, \oc8051_golden_model_1.PC [3]);
  or (_05404_, \oc8051_golden_model_1.PC [2], _05403_);
  or (_05405_, _05404_, _05402_);
  or (_05406_, _05405_, _00429_);
  not (_05407_, \oc8051_golden_model_1.PC [1]);
  or (_05408_, _05407_, \oc8051_golden_model_1.PC [0]);
  or (_05409_, _05408_, _05404_);
  or (_05410_, _05409_, _00388_);
  and (_05411_, _05410_, _05406_);
  not (_05412_, \oc8051_golden_model_1.PC [2]);
  or (_05413_, _05412_, \oc8051_golden_model_1.PC [3]);
  or (_05415_, _05413_, _05402_);
  or (_05416_, _05415_, _00265_);
  or (_05418_, _05413_, _05408_);
  or (_05419_, _05418_, _00224_);
  and (_05420_, _05419_, _05416_);
  and (_05422_, _05420_, _05411_);
  and (_05423_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  and (_05424_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  and (_05426_, _05424_, _05423_);
  nand (_05427_, _05426_, _00612_);
  nand (_05428_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_05430_, _05428_, _05408_);
  or (_05431_, _05430_, _00558_);
  and (_05432_, _05431_, _05427_);
  or (_05434_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_05435_, _05434_, _05402_);
  or (_05436_, _05435_, _00070_);
  or (_05438_, _05434_, _05408_);
  or (_05439_, _05438_, _00029_);
  and (_05440_, _05439_, _05436_);
  and (_05442_, _05440_, _05432_);
  and (_05443_, _05442_, _05422_);
  not (_05444_, \oc8051_golden_model_1.PC [0]);
  or (_05446_, \oc8051_golden_model_1.PC [1], _05444_);
  or (_05447_, _05446_, _05428_);
  or (_05448_, _05447_, _00511_);
  or (_05449_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_05450_, _05449_, _05428_);
  or (_05451_, _05450_, _00470_);
  and (_05452_, _05451_, _05448_);
  or (_05453_, _05434_, _05449_);
  or (_05454_, _05453_, _43974_);
  or (_05455_, _05434_, _05446_);
  or (_05456_, _05455_, _44015_);
  and (_05457_, _05456_, _05454_);
  and (_05458_, _05457_, _05452_);
  or (_05459_, _05446_, _05404_);
  or (_05460_, _05459_, _00347_);
  or (_05461_, _05449_, _05404_);
  or (_05462_, _05461_, _00306_);
  and (_05463_, _05462_, _05460_);
  or (_05464_, _05446_, _05413_);
  or (_05465_, _05464_, _00178_);
  or (_05466_, _05449_, _05413_);
  or (_05468_, _05466_, _00111_);
  and (_05469_, _05468_, _05465_);
  and (_05471_, _05469_, _05463_);
  and (_05472_, _05471_, _05458_);
  and (_05473_, _05472_, _05443_);
  or (_05475_, _05405_, _00394_);
  or (_05476_, _05409_, _00353_);
  and (_05477_, _05476_, _05475_);
  or (_05479_, _05415_, _00230_);
  or (_05480_, _05418_, _00189_);
  and (_05481_, _05480_, _05479_);
  and (_05483_, _05481_, _05477_);
  nand (_05484_, _05426_, _00567_);
  or (_05485_, _05430_, _00517_);
  and (_05487_, _05485_, _05484_);
  or (_05488_, _05435_, _00035_);
  or (_05489_, _05438_, _44021_);
  and (_05491_, _05489_, _05488_);
  and (_05492_, _05491_, _05487_);
  and (_05493_, _05492_, _05483_);
  or (_05495_, _05447_, _00476_);
  or (_05496_, _05450_, _00435_);
  and (_05497_, _05496_, _05495_);
  or (_05499_, _05453_, _43939_);
  or (_05500_, _05455_, _43980_);
  and (_05501_, _05500_, _05499_);
  and (_05502_, _05501_, _05497_);
  or (_05503_, _05459_, _00312_);
  or (_05504_, _05461_, _00271_);
  and (_05505_, _05504_, _05503_);
  or (_05506_, _05464_, _00117_);
  or (_05507_, _05466_, _00076_);
  and (_05508_, _05507_, _05506_);
  and (_05509_, _05508_, _05505_);
  and (_05510_, _05509_, _05502_);
  and (_05511_, _05510_, _05493_);
  and (_05512_, _05511_, _05473_);
  or (_05513_, _05405_, _00419_);
  or (_05514_, _05409_, _00378_);
  and (_05515_, _05514_, _05513_);
  or (_05516_, _05415_, _00255_);
  or (_05517_, _05418_, _00214_);
  and (_05518_, _05517_, _05516_);
  and (_05519_, _05518_, _05515_);
  nand (_05521_, _05426_, _00602_);
  or (_05522_, _05430_, _00542_);
  and (_05524_, _05522_, _05521_);
  or (_05525_, _05435_, _00060_);
  or (_05526_, _05438_, _00019_);
  and (_05528_, _05526_, _05525_);
  and (_05529_, _05528_, _05524_);
  and (_05530_, _05529_, _05519_);
  or (_05532_, _05447_, _00501_);
  or (_05533_, _05450_, _00460_);
  and (_05534_, _05533_, _05532_);
  or (_05536_, _05453_, _43964_);
  or (_05537_, _05455_, _44005_);
  and (_05538_, _05537_, _05536_);
  and (_05540_, _05538_, _05534_);
  or (_05541_, _05459_, _00337_);
  or (_05542_, _05461_, _00296_);
  and (_05544_, _05542_, _05541_);
  or (_05545_, _05464_, _00156_);
  or (_05546_, _05466_, _00101_);
  and (_05548_, _05546_, _05545_);
  and (_05549_, _05548_, _05544_);
  and (_05550_, _05549_, _05540_);
  and (_05552_, _05550_, _05530_);
  or (_05553_, _05405_, _00424_);
  or (_05554_, _05409_, _00383_);
  and (_05555_, _05554_, _05553_);
  or (_05556_, _05415_, _00260_);
  or (_05557_, _05418_, _00219_);
  and (_05558_, _05557_, _05556_);
  and (_05559_, _05558_, _05555_);
  nand (_05560_, _05426_, _00607_);
  or (_05561_, _05430_, _00550_);
  and (_05562_, _05561_, _05560_);
  or (_05563_, _05435_, _00065_);
  or (_05564_, _05438_, _00024_);
  and (_05565_, _05564_, _05563_);
  and (_05566_, _05565_, _05562_);
  and (_05567_, _05566_, _05559_);
  or (_05568_, _05447_, _00506_);
  or (_05569_, _05450_, _00465_);
  and (_05570_, _05569_, _05568_);
  or (_05571_, _05453_, _43969_);
  or (_05572_, _05455_, _44010_);
  and (_05574_, _05572_, _05571_);
  and (_05575_, _05574_, _05570_);
  or (_05577_, _05459_, _00342_);
  or (_05578_, _05461_, _00301_);
  and (_05579_, _05578_, _05577_);
  or (_05581_, _05464_, _00167_);
  or (_05582_, _05466_, _00106_);
  and (_05583_, _05582_, _05581_);
  and (_05585_, _05583_, _05579_);
  and (_05586_, _05585_, _05575_);
  nand (_05587_, _05586_, _05567_);
  or (_05589_, _05587_, _05552_);
  not (_05590_, _05589_);
  and (_05591_, _05590_, _05512_);
  or (_05593_, _05405_, _00409_);
  or (_05594_, _05409_, _00368_);
  and (_05595_, _05594_, _05593_);
  or (_05597_, _05415_, _00245_);
  or (_05598_, _05418_, _00204_);
  and (_05599_, _05598_, _05597_);
  and (_05601_, _05599_, _05595_);
  nand (_05602_, _05426_, _00591_);
  or (_05603_, _05430_, _00532_);
  and (_05605_, _05603_, _05602_);
  or (_05606_, _05435_, _00050_);
  or (_05607_, _05438_, _00009_);
  and (_05608_, _05607_, _05606_);
  and (_05609_, _05608_, _05605_);
  and (_05610_, _05609_, _05601_);
  or (_05611_, _05447_, _00491_);
  or (_05612_, _05450_, _00450_);
  and (_05613_, _05612_, _05611_);
  or (_05614_, _05453_, _43954_);
  or (_05615_, _05455_, _43995_);
  and (_05616_, _05615_, _05614_);
  and (_05617_, _05616_, _05613_);
  or (_05618_, _05459_, _00327_);
  or (_05619_, _05461_, _00286_);
  and (_05620_, _05619_, _05618_);
  or (_05621_, _05464_, _00134_);
  or (_05622_, _05466_, _00091_);
  and (_05623_, _05622_, _05621_);
  and (_05624_, _05623_, _05620_);
  and (_05625_, _05624_, _05617_);
  nand (_05627_, _05625_, _05610_);
  or (_05628_, _05405_, _00414_);
  or (_05630_, _05409_, _00373_);
  and (_05631_, _05630_, _05628_);
  or (_05632_, _05415_, _00250_);
  or (_05634_, _05418_, _00209_);
  and (_05635_, _05634_, _05632_);
  and (_05636_, _05635_, _05631_);
  nand (_05638_, _05426_, _00597_);
  or (_05639_, _05430_, _00537_);
  and (_05640_, _05639_, _05638_);
  or (_05642_, _05435_, _00055_);
  or (_05643_, _05438_, _00014_);
  and (_05644_, _05643_, _05642_);
  and (_05646_, _05644_, _05640_);
  and (_05647_, _05646_, _05636_);
  or (_05648_, _05447_, _00496_);
  or (_05650_, _05450_, _00455_);
  and (_05651_, _05650_, _05648_);
  or (_05652_, _05453_, _43959_);
  or (_05654_, _05455_, _44000_);
  and (_05655_, _05654_, _05652_);
  and (_05656_, _05655_, _05651_);
  or (_05658_, _05459_, _00332_);
  or (_05659_, _05461_, _00291_);
  and (_05660_, _05659_, _05658_);
  or (_05661_, _05464_, _00145_);
  or (_05662_, _05466_, _00096_);
  and (_05663_, _05662_, _05661_);
  and (_05664_, _05663_, _05660_);
  and (_05665_, _05664_, _05656_);
  nand (_05666_, _05665_, _05647_);
  or (_05667_, _05666_, _05627_);
  not (_05668_, _05667_);
  or (_05669_, _05405_, _00399_);
  or (_05670_, _05409_, _00358_);
  and (_05671_, _05670_, _05669_);
  or (_05672_, _05415_, _00235_);
  or (_05673_, _05418_, _00194_);
  and (_05674_, _05673_, _05672_);
  and (_05675_, _05674_, _05671_);
  nand (_05676_, _05426_, _00575_);
  or (_05677_, _05430_, _00522_);
  and (_05678_, _05677_, _05676_);
  or (_05680_, _05435_, _00040_);
  or (_05681_, _05438_, _44026_);
  and (_05683_, _05681_, _05680_);
  and (_05684_, _05683_, _05678_);
  and (_05685_, _05684_, _05675_);
  or (_05687_, _05447_, _00481_);
  or (_05688_, _05450_, _00440_);
  and (_05689_, _05688_, _05687_);
  or (_05691_, _05453_, _43944_);
  or (_05692_, _05455_, _43985_);
  and (_05693_, _05692_, _05691_);
  and (_05695_, _05693_, _05689_);
  or (_05696_, _05459_, _00317_);
  or (_05697_, _05461_, _00276_);
  and (_05699_, _05697_, _05696_);
  or (_05700_, _05464_, _00122_);
  or (_05701_, _05466_, _00081_);
  and (_05703_, _05701_, _05700_);
  and (_05704_, _05703_, _05699_);
  and (_05705_, _05704_, _05695_);
  and (_05707_, _05705_, _05685_);
  or (_05708_, _05405_, _00404_);
  or (_05709_, _05409_, _00363_);
  and (_05711_, _05709_, _05708_);
  or (_05712_, _05415_, _00240_);
  or (_05713_, _05418_, _00199_);
  and (_05714_, _05713_, _05712_);
  and (_05715_, _05714_, _05711_);
  nand (_05716_, _05426_, _00583_);
  or (_05717_, _05430_, _00527_);
  and (_05718_, _05717_, _05716_);
  or (_05719_, _05435_, _00045_);
  or (_05720_, _05438_, _00004_);
  and (_05721_, _05720_, _05719_);
  and (_05722_, _05721_, _05718_);
  and (_05723_, _05722_, _05715_);
  or (_05724_, _05447_, _00486_);
  or (_05725_, _05450_, _00445_);
  and (_05726_, _05725_, _05724_);
  or (_05727_, _05453_, _43949_);
  or (_05728_, _05455_, _43990_);
  and (_05729_, _05728_, _05727_);
  and (_05730_, _05729_, _05726_);
  or (_05731_, _05459_, _00322_);
  or (_05733_, _05461_, _00281_);
  and (_05734_, _05733_, _05731_);
  or (_05736_, _05464_, _00127_);
  or (_05737_, _05466_, _00086_);
  and (_05738_, _05737_, _05736_);
  and (_05740_, _05738_, _05734_);
  and (_05741_, _05740_, _05730_);
  nand (_05742_, _05741_, _05723_);
  not (_05744_, _05742_);
  and (_05745_, _05744_, _05707_);
  and (_05746_, _05745_, _05668_);
  and (_05748_, _05746_, _05591_);
  not (_05749_, _05748_);
  or (_05750_, _05742_, _05707_);
  or (_05752_, _05750_, _05667_);
  and (_05753_, _05586_, _05567_);
  or (_05754_, _05753_, _05552_);
  nand (_05756_, _05472_, _05443_);
  or (_05757_, _05511_, _05756_);
  or (_05758_, _05757_, _05754_);
  or (_05760_, _05758_, _05752_);
  or (_05761_, _05511_, _05473_);
  or (_05762_, _05761_, _05589_);
  or (_05764_, _05762_, _05752_);
  and (_05765_, _05764_, _05760_);
  nand (_05766_, _05550_, _05530_);
  or (_05767_, _05587_, _05766_);
  or (_05768_, _05767_, _05761_);
  or (_05769_, _05768_, _05752_);
  or (_05770_, _05753_, _05766_);
  or (_05771_, _05770_, _05761_);
  or (_05772_, _05771_, _05752_);
  and (_05773_, _05772_, _05769_);
  or (_05774_, _05770_, _05757_);
  or (_05775_, _05774_, _05752_);
  or (_05776_, _05761_, _05754_);
  or (_05777_, _05776_, _05752_);
  and (_05778_, _05777_, _05775_);
  and (_05779_, _05778_, _05773_);
  and (_05780_, _05779_, _05765_);
  nor (_05781_, _05767_, _05757_);
  not (_05782_, _05750_);
  not (_05783_, _05666_);
  and (_05784_, _05783_, _05627_);
  and (_05786_, _05784_, _05782_);
  and (_05787_, _05786_, _05781_);
  not (_05789_, _05752_);
  nor (_05790_, _05757_, _05589_);
  and (_05791_, _05790_, _05789_);
  nor (_05793_, _05791_, _05787_);
  and (_05794_, _05793_, _05780_);
  or (_05795_, _05794_, \oc8051_golden_model_1.PC [0]);
  not (_05797_, _05781_);
  or (_05798_, _05744_, _05707_);
  or (_05799_, _05798_, _05667_);
  nor (_05801_, _05799_, _05797_);
  not (_05802_, _05801_);
  not (_05803_, _05790_);
  or (_05805_, _05799_, _05803_);
  and (_05806_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_05807_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_05809_, _05807_, _05806_);
  or (_05810_, _05809_, _05805_);
  and (_05811_, _05805_, \oc8051_golden_model_1.PC [0]);
  nand (_05813_, _05811_, _05780_);
  nand (_05814_, _05813_, _05810_);
  nand (_05815_, _05814_, _05793_);
  and (_05817_, _05815_, _05802_);
  nand (_05818_, _05817_, _05795_);
  not (_05819_, _05767_);
  and (_05820_, _05819_, _05512_);
  and (_05821_, _05820_, _05789_);
  not (_05822_, _05821_);
  and (_05823_, _05789_, _05591_);
  not (_05824_, _05512_);
  nor (_05825_, _05770_, _05824_);
  and (_05826_, _05825_, _05789_);
  nor (_05827_, _05826_, _05823_);
  and (_05828_, _05827_, _05822_);
  and (_05829_, _05781_, _05789_);
  not (_05830_, _05829_);
  and (_05831_, _05511_, _05756_);
  not (_05832_, _05831_);
  or (_05833_, _05832_, _05770_);
  or (_05834_, _05833_, _05752_);
  or (_05835_, _05832_, _05754_);
  or (_05836_, _05835_, _05752_);
  and (_05837_, _05836_, _05834_);
  and (_05839_, _05837_, _05830_);
  and (_05840_, _05831_, _05819_);
  and (_05842_, _05840_, _05789_);
  not (_05843_, _05842_);
  or (_05844_, _05754_, _05824_);
  or (_05846_, _05844_, _05752_);
  or (_05847_, _05832_, _05589_);
  or (_05848_, _05847_, _05752_);
  and (_05850_, _05848_, _05846_);
  and (_05851_, _05850_, _05843_);
  and (_05852_, _05851_, _05839_);
  and (_05854_, _05852_, _05828_);
  not (_05855_, \oc8051_golden_model_1.ACC [0]);
  and (_05856_, _05855_, \oc8051_golden_model_1.PC [0]);
  and (_05858_, \oc8051_golden_model_1.ACC [0], _05444_);
  or (_05859_, _05858_, _05802_);
  or (_05860_, _05859_, _05856_);
  and (_05862_, _05860_, _05854_);
  nand (_05863_, _05862_, _05818_);
  nor (_05864_, _05854_, \oc8051_golden_model_1.PC [0]);
  not (_05866_, _05864_);
  and (_05867_, _05866_, _05863_);
  or (_05868_, _05794_, \oc8051_golden_model_1.PC [1]);
  not (_05870_, _05805_);
  and (_05871_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_05872_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_05873_, _05872_, _05871_);
  and (_05874_, _05873_, _05806_);
  nor (_05875_, _05873_, _05806_);
  nor (_05876_, _05875_, _05874_);
  and (_05877_, _05876_, _05870_);
  and (_05878_, _05446_, _05408_);
  not (_05879_, _05878_);
  and (_05880_, _05879_, _05805_);
  and (_05881_, _05880_, _05780_);
  or (_05882_, _05881_, _05877_);
  and (_05883_, _05854_, _05793_);
  nand (_05884_, _05883_, _05882_);
  nand (_05885_, _05884_, _05868_);
  nand (_05886_, _05885_, _05802_);
  not (_05887_, \oc8051_golden_model_1.ACC [1]);
  nor (_05888_, _05878_, _05887_);
  and (_05889_, _05878_, _05887_);
  nor (_05890_, _05889_, _05888_);
  and (_05892_, _05890_, _05858_);
  nor (_05893_, _05890_, _05858_);
  nor (_05895_, _05893_, _05892_);
  and (_05896_, _05895_, _05801_);
  nor (_05897_, _05854_, \oc8051_golden_model_1.PC [1]);
  nor (_05899_, _05897_, _05896_);
  and (_05900_, _05899_, _05886_);
  or (_05901_, _05900_, _05867_);
  nor (_05903_, _05892_, _05888_);
  and (_05904_, _05423_, \oc8051_golden_model_1.PC [2]);
  and (_05905_, _05402_, _05412_);
  nor (_05907_, _05905_, _05904_);
  and (_05908_, _05907_, \oc8051_golden_model_1.ACC [2]);
  nor (_05909_, _05907_, \oc8051_golden_model_1.ACC [2]);
  nor (_05911_, _05909_, _05908_);
  not (_05912_, _05911_);
  and (_05913_, _05912_, _05903_);
  nor (_05915_, _05912_, _05903_);
  nor (_05916_, _05915_, _05913_);
  and (_05917_, _05916_, _05801_);
  and (_05919_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_05920_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_05921_, _05920_, _05919_);
  not (_05923_, _05921_);
  or (_05924_, _05923_, _05780_);
  nand (_05925_, _05907_, _05780_);
  nand (_05926_, _05925_, _05924_);
  nand (_05927_, _05926_, _05805_);
  nor (_05928_, _05874_, _05871_);
  and (_05929_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_05930_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_05931_, _05930_, _05929_);
  not (_05932_, _05931_);
  nor (_05933_, _05932_, _05928_);
  and (_05934_, _05932_, _05928_);
  nor (_05935_, _05934_, _05933_);
  not (_05936_, _05935_);
  or (_05937_, _05936_, _05805_);
  and (_05938_, _05937_, _05793_);
  nand (_05939_, _05938_, _05927_);
  or (_05940_, _05921_, _05793_);
  and (_05941_, _05940_, _05802_);
  and (_05942_, _05941_, _05939_);
  or (_05943_, _05942_, _05917_);
  nand (_05944_, _05943_, _05854_);
  nor (_05945_, _05923_, _05854_);
  not (_05946_, _05945_);
  and (_05947_, _05946_, _05944_);
  nor (_05948_, _05915_, _05908_);
  not (_05949_, _05415_);
  nor (_05950_, _05904_, _05403_);
  nor (_05951_, _05950_, _05949_);
  nor (_05952_, _05951_, \oc8051_golden_model_1.ACC [3]);
  and (_05953_, _05951_, \oc8051_golden_model_1.ACC [3]);
  nor (_05954_, _05953_, _05952_);
  and (_05955_, _05954_, _05948_);
  nor (_05956_, _05954_, _05948_);
  nor (_05957_, _05956_, _05955_);
  and (_05958_, _05957_, _05801_);
  and (_05959_, _05805_, _05951_);
  nand (_05960_, _05959_, _05780_);
  nor (_05961_, _05933_, _05929_);
  and (_05962_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_05963_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_05964_, _05963_, _05962_);
  not (_05965_, _05964_);
  nor (_05966_, _05965_, _05961_);
  and (_05967_, _05965_, _05961_);
  nor (_05968_, _05967_, _05966_);
  or (_05969_, _05968_, _05805_);
  nand (_05970_, _05969_, _05960_);
  nand (_05971_, _05970_, _05793_);
  and (_05972_, _05424_, \oc8051_golden_model_1.PC [1]);
  nor (_05973_, _05919_, \oc8051_golden_model_1.PC [3]);
  nor (_05974_, _05973_, _05972_);
  or (_05975_, _05974_, _05794_);
  and (_05976_, _05975_, _05971_);
  nand (_05977_, _05976_, _05802_);
  nand (_05978_, _05977_, _05854_);
  nor (_05979_, _05978_, _05958_);
  nor (_05980_, _05974_, _05854_);
  or (_05981_, _05980_, _05979_);
  or (_05982_, _05981_, _05947_);
  or (_05983_, _05982_, _05901_);
  or (_05984_, _05983_, _00517_);
  nand (_05985_, _05866_, _05863_);
  nand (_05986_, _05899_, _05886_);
  or (_05987_, _05986_, _05985_);
  or (_05988_, _05987_, _05982_);
  or (_05989_, _05988_, _00476_);
  and (_05990_, _05989_, _05984_);
  or (_05991_, _05900_, _05985_);
  nor (_05992_, _05980_, _05979_);
  or (_05993_, _05992_, _05947_);
  or (_05994_, _05993_, _05991_);
  or (_05995_, _05994_, _00230_);
  nand (_05996_, _05946_, _05944_);
  or (_05997_, _05992_, _05996_);
  or (_05998_, _05997_, _05991_);
  or (_05999_, _05998_, _00035_);
  and (_06000_, _05999_, _05995_);
  and (_06001_, _06000_, _05990_);
  or (_06002_, _05997_, _05901_);
  or (_06003_, _06002_, _44021_);
  or (_06004_, _05997_, _05987_);
  or (_06005_, _06004_, _43980_);
  and (_06006_, _06005_, _06003_);
  or (_06007_, _05993_, _05901_);
  or (_06008_, _06007_, _00189_);
  or (_06009_, _05986_, _05867_);
  or (_06010_, _06009_, _05993_);
  or (_06011_, _06010_, _00076_);
  and (_06012_, _06011_, _06008_);
  and (_06013_, _06012_, _06006_);
  and (_06014_, _06013_, _06001_);
  or (_06015_, _05981_, _05996_);
  or (_06016_, _06015_, _05901_);
  or (_06017_, _06016_, _00353_);
  or (_06018_, _06015_, _06009_);
  or (_06019_, _06018_, _00271_);
  and (_06020_, _06019_, _06017_);
  nor (_06021_, _05991_, _05982_);
  nand (_06022_, _06021_, _00567_);
  or (_06023_, _06009_, _05982_);
  or (_06024_, _06023_, _00435_);
  and (_06025_, _06024_, _06022_);
  and (_06026_, _06025_, _06020_);
  or (_06027_, _05993_, _05987_);
  or (_06028_, _06027_, _00117_);
  or (_06029_, _06009_, _05997_);
  or (_06030_, _06029_, _43939_);
  and (_06031_, _06030_, _06028_);
  or (_06032_, _06015_, _05991_);
  or (_06033_, _06032_, _00394_);
  or (_06034_, _06015_, _05987_);
  or (_06035_, _06034_, _00312_);
  and (_06036_, _06035_, _06033_);
  and (_06037_, _06036_, _06031_);
  and (_06038_, _06037_, _06026_);
  nand (_06039_, _06038_, _06014_);
  nand (_06040_, _06021_, _00597_);
  or (_06041_, _05998_, _00055_);
  and (_06042_, _06041_, _06040_);
  or (_06043_, _05983_, _00537_);
  or (_06044_, _06034_, _00332_);
  and (_06045_, _06044_, _06043_);
  and (_06046_, _06045_, _06042_);
  or (_06047_, _06032_, _00414_);
  or (_06048_, _05994_, _00250_);
  and (_06049_, _06048_, _06047_);
  or (_06050_, _06007_, _00209_);
  or (_06051_, _06004_, _44000_);
  and (_06052_, _06051_, _06050_);
  and (_06053_, _06052_, _06049_);
  and (_06054_, _06053_, _06046_);
  or (_06055_, _05988_, _00496_);
  or (_06056_, _06023_, _00455_);
  and (_06057_, _06056_, _06055_);
  or (_06058_, _06018_, _00291_);
  or (_06059_, _06027_, _00145_);
  and (_06060_, _06059_, _06058_);
  and (_06061_, _06060_, _06057_);
  or (_06062_, _06016_, _00373_);
  or (_06063_, _06002_, _00014_);
  and (_06064_, _06063_, _06062_);
  or (_06065_, _06010_, _00096_);
  or (_06066_, _06029_, _43959_);
  and (_06067_, _06066_, _06065_);
  and (_06068_, _06067_, _06064_);
  and (_06069_, _06068_, _06061_);
  and (_06070_, _06069_, _06054_);
  or (_06071_, _06070_, _06039_);
  nor (_06072_, _06071_, _05749_);
  nor (_06073_, _06039_, _05749_);
  not (_06074_, _06073_);
  nor (_06075_, _05846_, \oc8051_golden_model_1.SP [0]);
  not (_06076_, _05836_);
  or (_06077_, _06007_, _00194_);
  or (_06078_, _06027_, _00122_);
  and (_06079_, _06078_, _06077_);
  or (_06080_, _05998_, _00040_);
  or (_06081_, _06002_, _44026_);
  and (_06082_, _06081_, _06080_);
  and (_06083_, _06082_, _06079_);
  or (_06084_, _06034_, _00317_);
  or (_06085_, _06018_, _00276_);
  and (_06086_, _06085_, _06084_);
  or (_06087_, _05988_, _00481_);
  or (_06088_, _06023_, _00440_);
  and (_06089_, _06088_, _06087_);
  and (_06090_, _06089_, _06086_);
  and (_06091_, _06090_, _06083_);
  or (_06092_, _06029_, _43944_);
  or (_06093_, _06004_, _43985_);
  and (_06094_, _06093_, _06092_);
  or (_06095_, _05994_, _00235_);
  or (_06096_, _06010_, _00081_);
  and (_06097_, _06096_, _06095_);
  and (_06098_, _06097_, _06094_);
  nand (_06099_, _06021_, _00575_);
  or (_06100_, _05983_, _00522_);
  and (_06101_, _06100_, _06099_);
  or (_06102_, _06032_, _00399_);
  or (_06103_, _06016_, _00358_);
  and (_06104_, _06103_, _06102_);
  and (_06105_, _06104_, _06101_);
  and (_06106_, _06105_, _06098_);
  and (_06107_, _06106_, _06091_);
  not (_06108_, _06107_);
  not (_06109_, _05835_);
  and (_06110_, _06109_, _05786_);
  not (_06111_, _06110_);
  nor (_06112_, _06111_, _06039_);
  and (_06113_, _06112_, _06108_);
  not (_06114_, _05787_);
  and (_06115_, _05784_, _05742_);
  and (_06116_, _06115_, _05781_);
  not (_06117_, _06116_);
  nor (_06118_, _05783_, _05627_);
  and (_06119_, _06118_, _05744_);
  and (_06120_, _06119_, _05781_);
  not (_06121_, _06120_);
  and (_06122_, _05666_, _05627_);
  and (_06123_, _06122_, _05782_);
  and (_06124_, _06122_, _05742_);
  or (_06125_, _06124_, _06123_);
  and (_06126_, _06125_, _05781_);
  and (_06127_, _06122_, _05745_);
  and (_06128_, _06118_, _05742_);
  nor (_06129_, _06128_, _06127_);
  nor (_06130_, _06129_, _05797_);
  nor (_06131_, _06130_, _06126_);
  and (_06132_, _06131_, _06121_);
  and (_06133_, _06132_, _06117_);
  and (_06134_, _06133_, _06114_);
  nor (_06135_, _06134_, _06039_);
  and (_06136_, _06135_, _06107_);
  and (_06137_, _05742_, _05707_);
  and (_06138_, _06137_, _05668_);
  and (_06139_, _06138_, _05790_);
  not (_06140_, _06139_);
  nor (_06141_, _06140_, _06071_);
  not (_06142_, \oc8051_golden_model_1.SP [0]);
  nor (_06143_, _05760_, _06142_);
  not (_06144_, _05758_);
  and (_06145_, _06138_, _06144_);
  not (_06146_, _06145_);
  nor (_06147_, _06146_, _06071_);
  nor (_06148_, _06146_, _06039_);
  not (_06149_, _06148_);
  not (_06150_, _05768_);
  and (_06151_, _06150_, _05746_);
  and (_06152_, _06138_, _06150_);
  not (_06153_, _06152_);
  nor (_06154_, _06153_, _06071_);
  not (_06155_, _05762_);
  and (_06156_, _06138_, _06155_);
  not (_06157_, _06156_);
  or (_06158_, _06157_, _06071_);
  nor (_06159_, _06157_, _06039_);
  and (_06160_, _05786_, _06155_);
  not (_06161_, _06160_);
  nor (_06162_, _06161_, _06039_);
  and (_06163_, _06162_, _06108_);
  not (_06164_, _05777_);
  and (_06165_, _05825_, _05746_);
  not (_06166_, _06165_);
  and (_06167_, _06138_, _05825_);
  not (_06168_, _06167_);
  and (_06169_, _05825_, _05786_);
  and (_06170_, _06169_, _06070_);
  not (_06171_, _06169_);
  not (_06172_, _06039_);
  and (_06173_, _06021_, _00612_);
  nor (_06174_, _06027_, _00178_);
  nor (_06175_, _06174_, _06173_);
  nor (_06176_, _05983_, _00558_);
  nor (_06177_, _06018_, _00306_);
  nor (_06178_, _06177_, _06176_);
  and (_06179_, _06178_, _06175_);
  nor (_06180_, _06004_, _44015_);
  nor (_06181_, _06002_, _00029_);
  nor (_06182_, _06181_, _06180_);
  nor (_06183_, _06032_, _00429_);
  nor (_06184_, _05998_, _00070_);
  nor (_06185_, _06184_, _06183_);
  and (_06186_, _06185_, _06182_);
  and (_06187_, _06186_, _06179_);
  nor (_06188_, _05988_, _00511_);
  nor (_06189_, _06023_, _00470_);
  nor (_06190_, _06189_, _06188_);
  nor (_06191_, _06034_, _00347_);
  nor (_06192_, _05994_, _00265_);
  nor (_06193_, _06192_, _06191_);
  and (_06194_, _06193_, _06190_);
  nor (_06195_, _06016_, _00388_);
  nor (_06196_, _06007_, _00224_);
  nor (_06197_, _06196_, _06195_);
  nor (_06198_, _06010_, _00111_);
  nor (_06199_, _06029_, _43974_);
  nor (_06200_, _06199_, _06198_);
  and (_06201_, _06200_, _06197_);
  and (_06202_, _06201_, _06194_);
  and (_06203_, _06202_, _06187_);
  and (_06204_, _06203_, _06172_);
  and (_06205_, _06070_, _06039_);
  or (_06206_, _06205_, _06204_);
  not (_06207_, _06206_);
  and (_06208_, _06138_, _06109_);
  and (_06209_, _06138_, _05781_);
  nor (_06210_, _06209_, _06208_);
  nor (_06211_, _06210_, _06207_);
  and (_06212_, _06144_, _05746_);
  nor (_06213_, _06145_, _06212_);
  or (_06214_, _06213_, _06206_);
  and (_06215_, _06206_, _06156_);
  not (_06216_, \oc8051_golden_model_1.SP [3]);
  and (_06217_, _06155_, _05746_);
  and (_06218_, _06217_, _06216_);
  or (_06219_, _06218_, _06215_);
  and (_06220_, _05786_, _06150_);
  nor (_06221_, _06217_, _06156_);
  not (_06222_, _05771_);
  and (_06223_, _05786_, _06222_);
  nor (_06224_, _06223_, _06160_);
  nand (_06225_, _06224_, \oc8051_golden_model_1.PSW [3]);
  and (_06226_, _06225_, _06221_);
  or (_06227_, _06226_, _06220_);
  not (_06228_, _06070_);
  not (_06229_, _06220_);
  nand (_06230_, _06224_, _06229_);
  nand (_06231_, _06230_, _06228_);
  and (_06232_, _06231_, _06227_);
  or (_06233_, _06232_, _06152_);
  or (_06234_, _06233_, _06219_);
  or (_06235_, _06206_, _06153_);
  and (_06236_, _05786_, _06144_);
  nor (_06237_, _06236_, _06151_);
  and (_06238_, _06237_, _06235_);
  and (_06239_, _06238_, _06234_);
  not (_06240_, _06213_);
  nor (_06241_, _06237_, _06228_);
  or (_06242_, _06241_, _06240_);
  or (_06243_, _06242_, _06239_);
  and (_06244_, _06243_, _06214_);
  not (_06245_, _05774_);
  and (_06246_, _06125_, _06245_);
  not (_06247_, _06246_);
  and (_06248_, _06127_, _06245_);
  and (_06249_, _06118_, _06245_);
  nor (_06250_, _06249_, _06248_);
  and (_06251_, _06250_, _06247_);
  not (_06252_, _06251_);
  or (_06253_, _06252_, _06244_);
  and (_06254_, _06245_, _05746_);
  and (_06255_, _06138_, _06245_);
  nor (_06256_, _06255_, _06254_);
  or (_06257_, _06251_, _06070_);
  and (_06258_, _06257_, _06256_);
  and (_06259_, _06258_, _06253_);
  and (_06260_, _05790_, _05786_);
  not (_06261_, _06256_);
  and (_06262_, _06261_, _06206_);
  or (_06263_, _06262_, _06260_);
  or (_06264_, _06263_, _06259_);
  not (_06265_, _06260_);
  or (_06266_, _06265_, _06070_);
  and (_06267_, _06266_, _06140_);
  and (_06268_, _06267_, _06264_);
  and (_06269_, _06206_, _06139_);
  or (_06270_, _06269_, _05787_);
  or (_06271_, _06270_, _06268_);
  and (_06272_, _06123_, _06144_);
  and (_06273_, _06118_, _05745_);
  and (_06274_, _06273_, _06144_);
  nor (_06275_, _06274_, _06272_);
  not (_06276_, _05707_);
  and (_06277_, _06124_, _06276_);
  and (_06278_, _06277_, _06144_);
  nor (_06279_, _06278_, _06160_);
  and (_06280_, _06279_, _06275_);
  and (_06281_, _06137_, _05784_);
  and (_06282_, _06281_, _06144_);
  not (_06283_, _05798_);
  and (_06284_, _06283_, _05784_);
  and (_06285_, _06284_, _06144_);
  nor (_06286_, _06285_, _06282_);
  and (_06287_, _06286_, _06280_);
  and (_06288_, _06118_, _05782_);
  and (_06289_, _06288_, _06144_);
  nor (_06290_, _06129_, _05758_);
  nor (_06291_, _06290_, _06289_);
  and (_06292_, _06291_, _06287_);
  and (_06293_, _05790_, _05746_);
  and (_06294_, _05784_, _05745_);
  and (_06295_, _06294_, _06144_);
  nor (_06296_, _06295_, _06293_);
  nor (_06297_, _05833_, _05799_);
  nor (_06298_, _06297_, _06110_);
  and (_06299_, _06298_, _06296_);
  not (_06300_, _05844_);
  and (_06301_, _06300_, _05746_);
  not (_06302_, _05799_);
  and (_06303_, _05840_, _06302_);
  nor (_06304_, _06303_, _06301_);
  and (_06305_, _06138_, _05820_);
  nor (_06306_, _05847_, _05799_);
  nor (_06307_, _06306_, _06305_);
  and (_06308_, _06307_, _06304_);
  and (_06309_, _06308_, _06299_);
  and (_06310_, _06138_, _05591_);
  nor (_06311_, _06310_, _05748_);
  and (_06312_, _06311_, _06166_);
  and (_06313_, _06122_, _06137_);
  and (_06314_, _06313_, _06144_);
  nor (_06315_, _06314_, _06236_);
  and (_06316_, _06315_, _06312_);
  and (_06317_, _06316_, _06309_);
  and (_06318_, _06317_, _06292_);
  nor (_06319_, _06318_, _05923_);
  and (_06320_, _06318_, _05907_);
  nor (_06321_, _06320_, _06319_);
  not (_06322_, _05974_);
  nor (_06323_, _06318_, _06322_);
  not (_06324_, _05951_);
  and (_06325_, _06318_, _06324_);
  nor (_06326_, _06325_, _06323_);
  nor (_06327_, _06326_, _06321_);
  nor (_06328_, _06318_, _05444_);
  and (_06329_, _06318_, _05444_);
  nor (_06330_, _06329_, _06328_);
  not (_06331_, _06330_);
  nor (_06332_, _06329_, _05407_);
  and (_06333_, _06329_, _05407_);
  nor (_06334_, _06333_, _06332_);
  and (_06335_, _06334_, _06331_);
  and (_06336_, _06335_, _06327_);
  and (_06337_, _06336_, _00597_);
  nor (_06338_, _06334_, _06330_);
  and (_06339_, _06326_, _06321_);
  and (_06340_, _06339_, _06338_);
  and (_06341_, _06340_, _04563_);
  nor (_06342_, _06341_, _06337_);
  not (_06343_, _06321_);
  nor (_06344_, _06326_, _06343_);
  and (_06345_, _06344_, _06335_);
  and (_06346_, _06345_, _04534_);
  nor (_06347_, _06334_, _06331_);
  and (_06348_, _06339_, _06347_);
  and (_06349_, _06348_, _04553_);
  nor (_06350_, _06349_, _06346_);
  and (_06351_, _06350_, _06342_);
  and (_06352_, _06344_, _06338_);
  and (_06353_, _06352_, _04545_);
  and (_06354_, _06334_, _06330_);
  and (_06355_, _06339_, _06354_);
  and (_06356_, _06355_, _04559_);
  nor (_06357_, _06356_, _06353_);
  and (_06358_, _06326_, _06343_);
  and (_06359_, _06358_, _06335_);
  and (_06360_, _06359_, _04569_);
  and (_06361_, _06358_, _06347_);
  and (_06362_, _06361_, _04540_);
  nor (_06363_, _06362_, _06360_);
  and (_06364_, _06363_, _06357_);
  and (_06365_, _06364_, _06351_);
  and (_06366_, _06358_, _06338_);
  and (_06367_, _06366_, _04531_);
  and (_06368_, _06339_, _06335_);
  and (_06369_, _06368_, _04542_);
  nor (_06370_, _06369_, _06367_);
  and (_06371_, _06338_, _06327_);
  and (_06372_, _06371_, _04536_);
  and (_06373_, _06344_, _06354_);
  and (_06374_, _06373_, _04561_);
  nor (_06375_, _06374_, _06372_);
  and (_06376_, _06375_, _06370_);
  and (_06377_, _06354_, _06327_);
  and (_06378_, _06377_, _04551_);
  and (_06379_, _06347_, _06344_);
  and (_06380_, _06379_, _04548_);
  nor (_06381_, _06380_, _06378_);
  and (_06382_, _06347_, _06327_);
  and (_06383_, _06382_, _04529_);
  and (_06384_, _06358_, _06354_);
  and (_06385_, _06384_, _04557_);
  nor (_06386_, _06385_, _06383_);
  and (_06387_, _06386_, _06381_);
  and (_06388_, _06387_, _06376_);
  and (_06389_, _06388_, _06365_);
  or (_06390_, _06389_, _06114_);
  and (_06391_, _06390_, _06210_);
  and (_06392_, _06391_, _06271_);
  or (_06393_, _06392_, _06211_);
  and (_06394_, _05840_, _05786_);
  not (_06395_, _06394_);
  and (_06396_, _06138_, _05840_);
  nor (_06397_, _06396_, _06303_);
  and (_06398_, _06397_, _06395_);
  not (_06399_, _05833_);
  and (_06400_, _06399_, _05786_);
  not (_06401_, _06400_);
  and (_06402_, _06138_, _06399_);
  nor (_06403_, _06402_, _06297_);
  and (_06404_, _06403_, _06401_);
  and (_06405_, _06404_, _06398_);
  and (_06406_, _06300_, _05786_);
  not (_06407_, _06406_);
  not (_06408_, _05847_);
  and (_06409_, _06408_, _05786_);
  not (_06410_, _06409_);
  and (_06411_, _06138_, _06408_);
  nor (_06412_, _06411_, _06306_);
  and (_06413_, _06412_, _06410_);
  and (_06414_, _06413_, _06407_);
  and (_06415_, _06414_, _06405_);
  and (_06416_, _06415_, _06393_);
  and (_06417_, _06138_, _06300_);
  nor (_06418_, _06415_, _06228_);
  or (_06419_, _06418_, _06417_);
  or (_06420_, _06419_, _06416_);
  not (_06421_, _06301_);
  nand (_06422_, _06417_, \oc8051_golden_model_1.SP [3]);
  and (_06423_, _06422_, _06421_);
  and (_06424_, _06423_, _06420_);
  and (_06425_, _06301_, _06206_);
  or (_06426_, _06425_, _06424_);
  and (_06427_, _06426_, _06171_);
  nor (_06428_, _06427_, _06170_);
  and (_06429_, _06428_, _06168_);
  and (_06430_, _06167_, \oc8051_golden_model_1.SP [3]);
  or (_06431_, _06430_, _06429_);
  and (_06432_, _06431_, _06166_);
  and (_06433_, _05786_, _05591_);
  nor (_06434_, _06206_, _06166_);
  or (_06435_, _06434_, _06433_);
  or (_06436_, _06435_, _06432_);
  nand (_06437_, _06433_, _06070_);
  and (_06438_, _06437_, _06436_);
  nor (_06439_, _06438_, _05748_);
  and (_06440_, _05820_, _05786_);
  and (_06441_, _06206_, _05748_);
  or (_06442_, _06441_, _06440_);
  nor (_06443_, _06442_, _06439_);
  not (_06444_, _06440_);
  nor (_06445_, _06444_, _06070_);
  nor (_06446_, _06445_, _06443_);
  and (_06447_, _06021_, _00607_);
  nor (_06448_, _06004_, _44010_);
  nor (_06449_, _06448_, _06447_);
  nor (_06450_, _06016_, _00383_);
  nor (_06451_, _06029_, _43969_);
  nor (_06452_, _06451_, _06450_);
  and (_06453_, _06452_, _06449_);
  nor (_06454_, _06018_, _00301_);
  nor (_06455_, _06002_, _00024_);
  nor (_06456_, _06455_, _06454_);
  nor (_06457_, _05994_, _00260_);
  nor (_06458_, _06010_, _00106_);
  nor (_06459_, _06458_, _06457_);
  and (_06460_, _06459_, _06456_);
  and (_06461_, _06460_, _06453_);
  nor (_06462_, _06027_, _00167_);
  nor (_06463_, _05998_, _00065_);
  nor (_06464_, _06463_, _06462_);
  nor (_06465_, _05983_, _00550_);
  nor (_06466_, _06032_, _00424_);
  nor (_06467_, _06466_, _06465_);
  and (_06468_, _06467_, _06464_);
  nor (_06469_, _06023_, _00465_);
  nor (_06470_, _06034_, _00342_);
  nor (_06471_, _06470_, _06469_);
  nor (_06472_, _05988_, _00506_);
  nor (_06473_, _06007_, _00219_);
  nor (_06474_, _06473_, _06472_);
  and (_06475_, _06474_, _06471_);
  and (_06476_, _06475_, _06468_);
  and (_06477_, _06476_, _06461_);
  nor (_06478_, _06477_, _06039_);
  not (_06479_, _06478_);
  nor (_06480_, _06165_, _06152_);
  and (_06481_, _06480_, _06421_);
  and (_06482_, _06256_, _06213_);
  nor (_06483_, _06139_, _05748_);
  and (_06484_, _06483_, _06210_);
  and (_06485_, _06484_, _06482_);
  and (_06486_, _06485_, _06481_);
  nor (_06487_, _06486_, _06479_);
  not (_06488_, _06487_);
  and (_06489_, _06478_, _06156_);
  not (_06490_, _06489_);
  and (_06491_, _06359_, _04505_);
  and (_06492_, _06368_, _04497_);
  nor (_06493_, _06492_, _06491_);
  and (_06494_, _06382_, _04486_);
  and (_06495_, _06352_, _04500_);
  nor (_06496_, _06495_, _06494_);
  and (_06497_, _06496_, _06493_);
  and (_06498_, _06384_, _04511_);
  and (_06499_, _06361_, _04495_);
  nor (_06500_, _06499_, _06498_);
  and (_06501_, _06366_, _04491_);
  and (_06502_, _06348_, _04507_);
  nor (_06503_, _06502_, _06501_);
  and (_06504_, _06503_, _06500_);
  and (_06505_, _06504_, _06497_);
  and (_06506_, _06336_, _00591_);
  and (_06507_, _06377_, _04523_);
  nor (_06508_, _06507_, _06506_);
  and (_06509_, _06371_, _04489_);
  and (_06510_, _06345_, _04484_);
  nor (_06511_, _06510_, _06509_);
  and (_06512_, _06511_, _06508_);
  and (_06513_, _06355_, _04513_);
  and (_06514_, _06340_, _04517_);
  nor (_06515_, _06514_, _06513_);
  and (_06516_, _06373_, _04515_);
  and (_06517_, _06379_, _04502_);
  nor (_06518_, _06517_, _06516_);
  and (_06519_, _06518_, _06515_);
  and (_06520_, _06519_, _06512_);
  and (_06521_, _06520_, _06505_);
  nor (_06522_, _06521_, _06114_);
  and (_06523_, _06124_, _06300_);
  and (_06524_, _06124_, _05840_);
  nor (_06525_, _06524_, _06523_);
  and (_06526_, _06124_, _05781_);
  not (_06527_, _06526_);
  and (_06528_, _06527_, _06525_);
  and (_06529_, _06124_, _06150_);
  and (_06530_, _06124_, _05591_);
  nor (_06531_, _06530_, _06529_);
  and (_06532_, _06167_, \oc8051_golden_model_1.SP [2]);
  and (_06533_, _06122_, _05744_);
  and (_06534_, _06533_, _05825_);
  nor (_06535_, _06534_, _06532_);
  and (_06536_, _06127_, _05790_);
  not (_06537_, _06536_);
  and (_06538_, _06533_, _06150_);
  and (_06539_, _06122_, _05820_);
  nor (_06540_, _06539_, _06538_);
  and (_06541_, _06540_, _06537_);
  and (_06542_, _06541_, _06535_);
  and (_06543_, _06542_, _06531_);
  and (_06544_, _06543_, _06528_);
  and (_06545_, _06124_, _06222_);
  and (_06546_, _06124_, _06155_);
  nor (_06547_, _06546_, _06545_);
  and (_06548_, _06124_, _05790_);
  and (_06549_, _06124_, _06144_);
  nor (_06550_, _06549_, _06548_);
  and (_06551_, _06550_, _06547_);
  and (_06552_, _06124_, _05825_);
  not (_06553_, _06552_);
  and (_06554_, _06533_, _06408_);
  and (_06555_, _06533_, _05840_);
  nor (_06556_, _06555_, _06554_);
  and (_06557_, _06124_, _06408_);
  and (_06558_, _06125_, _06399_);
  nor (_06559_, _06558_, _06557_);
  and (_06560_, _06559_, _06556_);
  and (_06561_, _06560_, _06553_);
  and (_06562_, _06127_, _05591_);
  and (_06563_, _06123_, _05591_);
  nor (_06564_, _06563_, _06562_);
  not (_06565_, _06564_);
  not (_06566_, \oc8051_golden_model_1.SP [2]);
  nor (_06567_, _06217_, _06417_);
  nor (_06568_, _06567_, _06566_);
  nor (_06569_, _06568_, _06565_);
  and (_06570_, _06569_, _06561_);
  and (_06571_, _06127_, _05781_);
  and (_06572_, _06127_, _06222_);
  nor (_06573_, _06572_, _06571_);
  and (_06574_, _06127_, _06399_);
  or (_06575_, _05790_, _05781_);
  and (_06576_, _06575_, _06123_);
  nor (_06577_, _06576_, _06574_);
  and (_06578_, _06577_, _06573_);
  and (_06579_, _06127_, _06144_);
  nor (_06580_, _06272_, _06579_);
  and (_06581_, _06123_, _06222_);
  not (_06582_, _06581_);
  and (_06583_, _06533_, _06300_);
  and (_06584_, _06533_, _06155_);
  nor (_06585_, _06584_, _06583_);
  and (_06586_, _06585_, _06582_);
  and (_06587_, _06586_, _06580_);
  and (_06588_, _06587_, _06578_);
  and (_06589_, _06588_, _06570_);
  and (_06590_, _06589_, _06551_);
  and (_06591_, _06590_, _06544_);
  not (_06592_, _06591_);
  nor (_06593_, _06592_, _06522_);
  not (_06594_, _06593_);
  nor (_06595_, _06023_, _00450_);
  nor (_06596_, _05994_, _00245_);
  nor (_06597_, _06596_, _06595_);
  nor (_06598_, _06007_, _00204_);
  nor (_06599_, _06029_, _43954_);
  nor (_06600_, _06599_, _06598_);
  and (_06601_, _06600_, _06597_);
  nor (_06602_, _06032_, _00409_);
  nor (_06603_, _05998_, _00050_);
  nor (_06604_, _06603_, _06602_);
  nor (_06605_, _06016_, _00368_);
  nor (_06606_, _06018_, _00286_);
  nor (_06607_, _06606_, _06605_);
  and (_06608_, _06607_, _06604_);
  and (_06609_, _06608_, _06601_);
  nor (_06610_, _06027_, _00134_);
  nor (_06611_, _06010_, _00091_);
  nor (_06612_, _06611_, _06610_);
  and (_06613_, _06021_, _00591_);
  nor (_06614_, _06004_, _43995_);
  nor (_06615_, _06614_, _06613_);
  and (_06616_, _06615_, _06612_);
  nor (_06617_, _05983_, _00532_);
  nor (_06618_, _06002_, _00009_);
  nor (_06619_, _06618_, _06617_);
  nor (_06620_, _05988_, _00491_);
  nor (_06621_, _06034_, _00327_);
  nor (_06622_, _06621_, _06620_);
  and (_06623_, _06622_, _06619_);
  and (_06624_, _06623_, _06616_);
  and (_06625_, _06624_, _06609_);
  not (_06626_, _06625_);
  nand (_06627_, _06265_, _06237_);
  nor (_06628_, _06627_, _06230_);
  nand (_06629_, _06628_, _06251_);
  nor (_06630_, _06440_, _06433_);
  and (_06631_, _06630_, _06171_);
  nand (_06632_, _06631_, _06415_);
  or (_06633_, _06632_, _06629_);
  and (_06634_, _06633_, _06626_);
  nor (_06635_, _06634_, _06594_);
  and (_06636_, _06635_, _06490_);
  and (_06637_, _06636_, _06488_);
  not (_06638_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_06639_, _06444_, _06107_);
  not (_06640_, _06639_);
  nor (_06641_, _06265_, _06107_);
  nor (_06642_, _06256_, _06071_);
  not (_06643_, _06236_);
  nor (_06644_, _06643_, _06107_);
  or (_06645_, _06229_, _06107_);
  nor (_06646_, _06224_, _06107_);
  and (_06647_, _06281_, _06155_);
  nand (_06648_, _05707_, _05666_);
  nor (_06649_, _06648_, _05762_);
  nor (_06650_, _06649_, _06647_);
  not (_06651_, _05776_);
  and (_06652_, _06281_, _06651_);
  and (_06653_, _06313_, _06222_);
  nor (_06654_, _06653_, _06652_);
  nor (_06655_, _06572_, _06160_);
  and (_06656_, _06655_, _06654_);
  nor (_06657_, _06281_, _05786_);
  or (_06658_, _06657_, _05771_);
  nand (_06659_, _06118_, _05707_);
  nor (_06660_, _06659_, _05771_);
  not (_06661_, _06660_);
  and (_06662_, _06661_, _06658_);
  and (_06663_, _06662_, _06656_);
  and (_06665_, _06663_, _06650_);
  or (_06666_, _06665_, _06646_);
  nand (_06667_, _06666_, _06157_);
  nand (_06668_, _06158_, _06667_);
  and (_06669_, _06217_, _06142_);
  nor (_06670_, _06669_, _06220_);
  not (_06671_, _06670_);
  and (_06672_, _06122_, _05707_);
  not (_06673_, _06672_);
  not (_06674_, _06281_);
  and (_06675_, _06659_, _06674_);
  and (_06676_, _06675_, _06673_);
  nor (_06677_, _06676_, _05768_);
  nor (_06678_, _06677_, _06671_);
  nand (_06679_, _06678_, _06668_);
  nand (_06680_, _06679_, _06645_);
  and (_06681_, _06680_, _06153_);
  or (_06682_, _06154_, _06681_);
  and (_06683_, _06151_, _06107_);
  and (_06684_, _06118_, _06137_);
  and (_06685_, _06684_, _06144_);
  nor (_06686_, _06274_, _06685_);
  and (_06687_, _06115_, _06144_);
  and (_06688_, _06687_, _05707_);
  nor (_06689_, _06688_, _06579_);
  and (_06690_, _06689_, _06686_);
  and (_06691_, _06690_, _06315_);
  not (_06692_, _06691_);
  nor (_06693_, _06692_, _06683_);
  and (_06694_, _06693_, _06682_);
  or (_06695_, _06694_, _06644_);
  nand (_06696_, _06695_, _06213_);
  nor (_06697_, _06213_, _06071_);
  nor (_06698_, _06697_, _06252_);
  nand (_06699_, _06698_, _06696_);
  and (_06700_, _06252_, _06107_);
  and (_06701_, _06115_, _06245_);
  and (_06702_, _06701_, _05707_);
  nor (_06703_, _06702_, _06261_);
  not (_06704_, _06703_);
  nor (_06705_, _06704_, _06700_);
  and (_06706_, _06705_, _06699_);
  or (_06707_, _06706_, _06642_);
  nor (_06708_, _06536_, _06260_);
  and (_06709_, _06281_, _05790_);
  not (_06710_, _06709_);
  and (_06711_, _06137_, _05666_);
  nor (_06712_, _06273_, _06711_);
  or (_06713_, _06712_, _05803_);
  and (_06714_, _06713_, _06710_);
  and (_06715_, _06714_, _06708_);
  and (_06716_, _06715_, _06707_);
  or (_06717_, _06716_, _06641_);
  and (_06718_, _06717_, _06140_);
  or (_06719_, _06718_, _06141_);
  nor (_06720_, _06684_, _06127_);
  or (_06721_, _06720_, _05797_);
  not (_06722_, _06313_);
  nor (_06723_, _06281_, _06273_);
  and (_06724_, _06723_, _06722_);
  or (_06725_, _06724_, _05797_);
  and (_06726_, _06725_, _06721_);
  and (_06727_, _06726_, _06719_);
  and (_06728_, _06336_, _00575_);
  and (_06729_, _06345_, _04393_);
  nor (_06730_, _06729_, _06728_);
  and (_06731_, _06384_, _04420_);
  and (_06732_, _06348_, _04416_);
  nor (_06733_, _06732_, _06731_);
  and (_06734_, _06733_, _06730_);
  and (_06735_, _06373_, _04424_);
  and (_06736_, _06352_, _04409_);
  nor (_06737_, _06736_, _06735_);
  and (_06738_, _06371_, _04398_);
  and (_06739_, _06382_, _04395_);
  nor (_06740_, _06739_, _06738_);
  and (_06741_, _06740_, _06737_);
  and (_06742_, _06741_, _06734_);
  and (_06743_, _06361_, _04404_);
  and (_06744_, _06368_, _04406_);
  nor (_06745_, _06744_, _06743_);
  and (_06746_, _06359_, _04414_);
  and (_06747_, _06366_, _04400_);
  nor (_06748_, _06747_, _06746_);
  and (_06749_, _06748_, _06745_);
  and (_06750_, _06355_, _04422_);
  and (_06751_, _06340_, _04426_);
  nor (_06752_, _06751_, _06750_);
  and (_06753_, _06377_, _04432_);
  and (_06754_, _06379_, _04411_);
  nor (_06755_, _06754_, _06753_);
  and (_06756_, _06755_, _06752_);
  and (_06757_, _06756_, _06749_);
  and (_06758_, _06757_, _06742_);
  and (_06759_, _06758_, _05787_);
  nor (_06760_, _06759_, _06209_);
  and (_06761_, _06760_, _06727_);
  not (_06762_, _06209_);
  nor (_06763_, _06762_, _06071_);
  or (_06764_, _06763_, _06761_);
  and (_06765_, _06281_, _06109_);
  nor (_06766_, _06765_, _06208_);
  and (_06767_, _06766_, _06764_);
  not (_06768_, _06208_);
  nor (_06769_, _06768_, _06071_);
  or (_06770_, _06769_, _06767_);
  and (_06771_, _06273_, _06399_);
  nor (_06772_, _06771_, _06574_);
  and (_06773_, _06281_, _06399_);
  and (_06774_, _06711_, _06399_);
  nor (_06775_, _06774_, _06773_);
  and (_06776_, _06775_, _06772_);
  and (_06777_, _06776_, _06770_);
  nor (_06778_, _06404_, _06108_);
  nor (_06779_, _06676_, _05847_);
  nor (_06780_, _06779_, _06778_);
  and (_06781_, _06780_, _06777_);
  nor (_06782_, _06413_, _06108_);
  not (_06783_, _05840_);
  nor (_06784_, _06676_, _06783_);
  nor (_06785_, _06784_, _06782_);
  and (_06786_, _06785_, _06781_);
  nor (_06787_, _06398_, _06108_);
  nor (_06788_, _06722_, _05844_);
  nor (_06789_, _06788_, _06406_);
  and (_06790_, _06273_, _06300_);
  not (_06791_, _06790_);
  and (_06792_, _06281_, _06300_);
  not (_06793_, _06792_);
  and (_06794_, _06127_, _06300_);
  and (_06795_, _06684_, _06300_);
  nor (_06796_, _06795_, _06794_);
  and (_06797_, _06796_, _06793_);
  and (_06798_, _06797_, _06791_);
  and (_06799_, _06798_, _06789_);
  not (_06800_, _06799_);
  nor (_06801_, _06800_, _06787_);
  and (_06802_, _06801_, _06786_);
  nor (_06803_, _06407_, _06107_);
  or (_06804_, _06803_, _06802_);
  and (_06805_, _06417_, _06142_);
  nor (_06806_, _06805_, _06301_);
  and (_06807_, _06806_, _06804_);
  nor (_06808_, _06421_, _06071_);
  or (_06809_, _06808_, _06807_);
  and (_06810_, _06127_, _05825_);
  not (_06811_, _05825_);
  and (_06812_, _06712_, _06657_);
  nor (_06813_, _06812_, _06811_);
  nor (_06814_, _06813_, _06810_);
  and (_06815_, _06814_, _06809_);
  nor (_06816_, _06171_, _06107_);
  or (_06817_, _06816_, _06815_);
  and (_06818_, _06167_, _06142_);
  nor (_06819_, _06818_, _06165_);
  and (_06820_, _06819_, _06817_);
  nor (_06821_, _06166_, _06071_);
  nor (_06822_, _06821_, _06820_);
  not (_06823_, _05591_);
  nor (_06824_, _06127_, _05786_);
  and (_06825_, _06824_, _06722_);
  and (_06826_, _06825_, _06675_);
  nor (_06827_, _06826_, _06823_);
  nor (_06828_, _06827_, _06822_);
  not (_06829_, _06433_);
  nor (_06830_, _06829_, _06107_);
  or (_06831_, _06830_, _06828_);
  and (_06832_, _06831_, _05749_);
  or (_06833_, _06832_, _06072_);
  and (_06834_, _06281_, _05820_);
  not (_06835_, _06834_);
  and (_06836_, _06273_, _05820_);
  nor (_06837_, _06836_, _06440_);
  and (_06838_, _06837_, _06835_);
  and (_06839_, _06684_, _05820_);
  and (_06840_, _06672_, _05820_);
  nor (_06841_, _06840_, _06839_);
  and (_06842_, _06841_, _06838_);
  nand (_06843_, _06842_, _06833_);
  nand (_06844_, _06843_, _06640_);
  or (_06845_, _06844_, _06638_);
  nor (_06846_, _06004_, _44005_);
  nor (_06847_, _06002_, _00019_);
  nor (_06848_, _06847_, _06846_);
  nor (_06849_, _05983_, _00542_);
  nor (_06850_, _06007_, _00214_);
  nor (_06851_, _06850_, _06849_);
  and (_06852_, _06851_, _06848_);
  nor (_06853_, _05998_, _00060_);
  nor (_06854_, _06010_, _00101_);
  nor (_06855_, _06854_, _06853_);
  nor (_06856_, _06032_, _00419_);
  nor (_06857_, _06018_, _00296_);
  nor (_06858_, _06857_, _06856_);
  and (_06859_, _06858_, _06855_);
  and (_06860_, _06859_, _06852_);
  nor (_06861_, _06023_, _00460_);
  nor (_06862_, _06034_, _00337_);
  nor (_06863_, _06862_, _06861_);
  and (_06864_, _06021_, _00602_);
  nor (_06865_, _05988_, _00501_);
  nor (_06866_, _06865_, _06864_);
  and (_06867_, _06866_, _06863_);
  nor (_06868_, _06016_, _00378_);
  nor (_06869_, _06029_, _43964_);
  nor (_06870_, _06869_, _06868_);
  nor (_06871_, _05994_, _00255_);
  nor (_06872_, _06027_, _00156_);
  nor (_06873_, _06872_, _06871_);
  and (_06874_, _06873_, _06870_);
  and (_06875_, _06874_, _06867_);
  and (_06876_, _06875_, _06860_);
  nor (_06877_, _06876_, _06039_);
  and (_06878_, _06486_, _06157_);
  not (_06879_, _06878_);
  and (_06880_, _06879_, _06877_);
  not (_06881_, _06880_);
  and (_06882_, _06021_, _00583_);
  nor (_06883_, _05998_, _00045_);
  nor (_06884_, _06883_, _06882_);
  nor (_06885_, _05983_, _00527_);
  nor (_06886_, _06034_, _00322_);
  nor (_06887_, _06886_, _06885_);
  and (_06888_, _06887_, _06884_);
  nor (_06889_, _06027_, _00127_);
  nor (_06890_, _06007_, _00199_);
  nor (_06891_, _06890_, _06889_);
  nor (_06892_, _06032_, _00404_);
  nor (_06893_, _05994_, _00240_);
  nor (_06894_, _06893_, _06892_);
  and (_06895_, _06894_, _06891_);
  and (_06896_, _06895_, _06888_);
  nor (_06897_, _05988_, _00486_);
  nor (_06898_, _06023_, _00445_);
  nor (_06899_, _06898_, _06897_);
  nor (_06900_, _06018_, _00281_);
  nor (_06901_, _06002_, _00004_);
  nor (_06902_, _06901_, _06900_);
  and (_06903_, _06902_, _06899_);
  nor (_06904_, _06016_, _00363_);
  nor (_06905_, _06010_, _00086_);
  nor (_06906_, _06905_, _06904_);
  nor (_06907_, _06029_, _43949_);
  nor (_06908_, _06004_, _43990_);
  nor (_06909_, _06908_, _06907_);
  and (_06910_, _06909_, _06906_);
  and (_06911_, _06910_, _06903_);
  and (_06912_, _06911_, _06896_);
  not (_06913_, _06912_);
  and (_06914_, _06913_, _06633_);
  and (_06915_, _06359_, _04460_);
  and (_06916_, _06368_, _04452_);
  nor (_06917_, _06916_, _06915_);
  and (_06918_, _06373_, _04470_);
  and (_06919_, _06379_, _04457_);
  nor (_06920_, _06919_, _06918_);
  and (_06921_, _06920_, _06917_);
  and (_06922_, _06384_, _04466_);
  and (_06923_, _06366_, _04445_);
  nor (_06924_, _06923_, _06922_);
  and (_06925_, _06355_, _04468_);
  and (_06926_, _06340_, _04472_);
  nor (_06927_, _06926_, _06925_);
  and (_06928_, _06927_, _06924_);
  and (_06929_, _06928_, _06921_);
  and (_06930_, _06382_, _04440_);
  and (_06931_, _06345_, _04438_);
  nor (_06932_, _06931_, _06930_);
  and (_06933_, _06377_, _04478_);
  and (_06934_, _06352_, _04455_);
  nor (_06935_, _06934_, _06933_);
  and (_06936_, _06935_, _06932_);
  and (_06937_, _06361_, _04450_);
  and (_06938_, _06348_, _04462_);
  nor (_06939_, _06938_, _06937_);
  and (_06940_, _06336_, _00583_);
  and (_06941_, _06371_, _04443_);
  nor (_06942_, _06941_, _06940_);
  and (_06943_, _06942_, _06939_);
  and (_06944_, _06943_, _06936_);
  and (_06945_, _06944_, _06929_);
  nor (_06946_, _06945_, _06114_);
  and (_06947_, _06217_, \oc8051_golden_model_1.SP [1]);
  not (_06948_, _06128_);
  nor (_06949_, _05820_, _06150_);
  nor (_06950_, _06949_, _06948_);
  nor (_06951_, _06950_, _06947_);
  and (_06952_, _06684_, _05825_);
  and (_06953_, _06539_, _05742_);
  nor (_06954_, _06953_, _06952_);
  and (_06955_, _06954_, _06951_);
  and (_06956_, _06124_, _06399_);
  and (_06957_, _06118_, _06283_);
  and (_06958_, _06957_, _05825_);
  or (_06959_, _06958_, _06557_);
  nor (_06960_, _06959_, _06956_);
  and (_06961_, _06960_, _06553_);
  and (_06962_, _06961_, _06955_);
  and (_06963_, _06531_, _06528_);
  and (_06964_, _06963_, _06962_);
  and (_06965_, _06128_, _06408_);
  and (_06966_, _05771_, _05758_);
  and (_06967_, _05833_, _05797_);
  and (_06968_, _06967_, _06966_);
  nor (_06969_, _06968_, _06948_);
  nor (_06970_, _06969_, _06965_);
  and (_06971_, _06128_, _05790_);
  and (_06972_, _06128_, _05591_);
  nor (_06973_, _06972_, _06971_);
  and (_06974_, _06973_, _06970_);
  and (_06975_, _06128_, _05840_);
  and (_06976_, _06128_, _06300_);
  nor (_06977_, _06976_, _06975_);
  and (_06978_, _06128_, _06155_);
  not (_06979_, \oc8051_golden_model_1.SP [1]);
  nor (_06980_, _06417_, _06167_);
  nor (_06981_, _06980_, _06979_);
  nor (_06982_, _06981_, _06978_);
  and (_06983_, _06982_, _06977_);
  and (_06984_, _06983_, _06974_);
  and (_06985_, _06984_, _06551_);
  and (_06986_, _06985_, _06964_);
  not (_06987_, _06986_);
  nor (_06988_, _06987_, _06946_);
  not (_06989_, _06988_);
  nor (_06990_, _06989_, _06914_);
  and (_06991_, _06990_, _06881_);
  not (_06992_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_06993_, _06843_, _06640_);
  or (_06994_, _06993_, _06992_);
  and (_06995_, _06994_, _06991_);
  nand (_06996_, _06995_, _06845_);
  not (_06997_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_06998_, _06993_, _06997_);
  not (_06999_, _06991_);
  not (_07000_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_07001_, _06844_, _07000_);
  and (_07002_, _07001_, _06999_);
  nand (_07003_, _07002_, _06998_);
  nand (_07004_, _07003_, _06996_);
  nand (_07005_, _07004_, _06637_);
  not (_07006_, _06637_);
  not (_07007_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_07008_, _06993_, _07007_);
  not (_07009_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_07010_, _06844_, _07009_);
  and (_07011_, _07010_, _06999_);
  nand (_07012_, _07011_, _07008_);
  not (_07013_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_07014_, _06844_, _07013_);
  not (_07015_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_07016_, _06993_, _07015_);
  and (_07017_, _07016_, _06991_);
  nand (_07018_, _07017_, _07014_);
  nand (_07019_, _07018_, _07012_);
  nand (_07020_, _07019_, _07006_);
  nand (_07021_, _07020_, _07005_);
  nand (_07022_, _07021_, _06446_);
  not (_07023_, _06446_);
  nand (_07024_, _06844_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_07025_, _06993_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_07026_, _07025_, _06999_);
  nand (_07027_, _07026_, _07024_);
  nand (_07028_, _06993_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand (_07029_, _06844_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_07030_, _07029_, _06991_);
  nand (_07031_, _07030_, _07028_);
  nand (_07032_, _07031_, _07027_);
  nand (_07033_, _07032_, _06637_);
  not (_07034_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_07035_, _06993_, _07034_);
  nand (_07036_, _06993_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_07037_, _07036_, _06999_);
  nand (_07038_, _07037_, _07035_);
  not (_07039_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_07040_, _06844_, _07039_);
  not (_07041_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_07042_, _06993_, _07041_);
  and (_07043_, _07042_, _06991_);
  nand (_07044_, _07043_, _07040_);
  nand (_07045_, _07044_, _07038_);
  nand (_07046_, _07045_, _07006_);
  nand (_07047_, _07046_, _07033_);
  nand (_07048_, _07047_, _07023_);
  and (_07049_, _07048_, _07022_);
  and (_07050_, _07049_, _06164_);
  nor (_07051_, _06294_, _05789_);
  and (_07052_, _07051_, _06723_);
  nor (_07053_, _07052_, _05776_);
  not (_07054_, _07053_);
  nor (_07055_, _07054_, _07050_);
  and (_07056_, _06277_, _06222_);
  not (_07057_, _07056_);
  nor (_07058_, _07057_, _06039_);
  and (_07059_, _07058_, _06107_);
  nor (_07060_, _07059_, _07055_);
  and (_07061_, _06581_, \oc8051_golden_model_1.SP [0]);
  nor (_07062_, _07061_, _06649_);
  and (_07063_, _07062_, _07060_);
  and (_07064_, _06115_, _06155_);
  not (_07065_, _07064_);
  nor (_07066_, _07065_, _07049_);
  nor (_07067_, _07066_, _06162_);
  and (_07068_, _07067_, _07063_);
  nor (_07069_, _07068_, _06163_);
  nor (_07070_, _07069_, _06159_);
  not (_07071_, _07070_);
  and (_07072_, _07071_, _06158_);
  nor (_07073_, _05764_, _06142_);
  nor (_07074_, _07073_, _07072_);
  not (_07075_, _06217_);
  nor (_07076_, _07075_, _06039_);
  and (_07077_, _07076_, _06107_);
  nor (_07078_, _06648_, _05768_);
  nor (_07079_, _07078_, _07077_);
  and (_07080_, _07079_, _07074_);
  and (_07081_, _06115_, _06150_);
  not (_07082_, _07081_);
  nor (_07083_, _07082_, _07049_);
  not (_07084_, _07083_);
  and (_07085_, _07084_, _07080_);
  nor (_07086_, _06153_, _06039_);
  nor (_07087_, _06229_, _06039_);
  and (_07088_, _07087_, _06107_);
  nor (_07089_, _07088_, _07086_);
  and (_07090_, _07089_, _07085_);
  nor (_07091_, _07090_, _06154_);
  or (_07092_, _07091_, _06151_);
  nand (_07093_, _06151_, _06142_);
  nand (_07094_, _07093_, _07092_);
  and (_07095_, _07094_, _06149_);
  nor (_07096_, _07095_, _06147_);
  and (_07097_, _06313_, _06245_);
  or (_07098_, _06248_, _07097_);
  nor (_07099_, _06659_, _05774_);
  or (_07100_, _07099_, _07098_);
  or (_07101_, _07100_, _07096_);
  nor (_07102_, _07101_, _06143_);
  nor (_07103_, _06140_, _06039_);
  not (_07104_, _06701_);
  nor (_07105_, _07049_, _07104_);
  nor (_07106_, _07105_, _07103_);
  and (_07107_, _07106_, _07102_);
  nor (_07108_, _07107_, _06141_);
  nor (_07109_, _07108_, _05791_);
  and (_07110_, _05791_, _06142_);
  nor (_07111_, _07110_, _07109_);
  nor (_07112_, _06648_, _05835_);
  or (_07113_, _07112_, _07111_);
  nor (_07114_, _07113_, _06136_);
  and (_07115_, _06115_, _06109_);
  not (_07116_, _07115_);
  nor (_07117_, _07116_, _07049_);
  nor (_07118_, _07117_, _06112_);
  and (_07119_, _07118_, _07114_);
  nor (_07120_, _07119_, _06113_);
  nor (_07121_, _07120_, _06076_);
  nor (_07122_, _05836_, \oc8051_golden_model_1.SP [0]);
  nor (_07123_, _07122_, _07121_);
  not (_07124_, _05848_);
  not (_07125_, _06402_);
  nor (_07126_, _07125_, _06039_);
  not (_07127_, _06297_);
  nor (_07128_, _07127_, _06039_);
  nor (_07129_, _07128_, _07126_);
  not (_07130_, _06411_);
  nor (_07131_, _07130_, _06039_);
  not (_07132_, _06306_);
  nor (_07133_, _07132_, _06039_);
  nor (_07134_, _07133_, _07131_);
  and (_07135_, _07134_, _07129_);
  nor (_07136_, _07135_, _06108_);
  nor (_07137_, _07136_, _07124_);
  not (_07138_, _07137_);
  nor (_07139_, _07138_, _07123_);
  nor (_07140_, _05848_, \oc8051_golden_model_1.SP [0]);
  nor (_07141_, _07140_, _07139_);
  not (_07142_, _05846_);
  nor (_07143_, _06397_, _06039_);
  and (_07144_, _07143_, _06107_);
  nor (_07145_, _07144_, _07142_);
  not (_07146_, _07145_);
  nor (_07147_, _07146_, _07141_);
  nor (_07148_, _07147_, _06075_);
  not (_07149_, _06648_);
  and (_07150_, _07149_, _05591_);
  nor (_07151_, _07150_, _07148_);
  nor (_07152_, _06829_, _06039_);
  and (_07153_, _06115_, _05591_);
  not (_07154_, _07153_);
  nor (_07155_, _07154_, _07049_);
  nor (_07156_, _07155_, _07152_);
  and (_07157_, _07156_, _07151_);
  and (_07158_, _07152_, _06108_);
  nor (_07159_, _07158_, _07157_);
  nor (_07160_, _06310_, _05823_);
  nor (_07161_, _07160_, _06142_);
  nor (_07162_, _07161_, _07159_);
  and (_07163_, _07162_, _06074_);
  nor (_07164_, _07163_, _06072_);
  and (_07165_, _07149_, _05820_);
  nor (_07166_, _07165_, _07164_);
  nor (_07167_, _06444_, _06039_);
  and (_07168_, _06115_, _05820_);
  not (_07169_, _07168_);
  nor (_07170_, _07169_, _07049_);
  nor (_07171_, _07170_, _07167_);
  and (_07172_, _07171_, _07166_);
  and (_07173_, _07167_, _06108_);
  nor (_07174_, _07173_, _07172_);
  and (_07175_, _07167_, _06913_);
  and (_07176_, _06877_, _05748_);
  and (_07177_, _06979_, \oc8051_golden_model_1.SP [0]);
  and (_07178_, \oc8051_golden_model_1.SP [1], _06142_);
  nor (_07179_, _07178_, _07177_);
  nor (_07180_, _07179_, _05846_);
  and (_07181_, _06913_, _06112_);
  and (_07182_, _06135_, _06912_);
  and (_07183_, _06273_, _06109_);
  and (_07184_, _06127_, _06109_);
  nor (_07185_, _07184_, _07183_);
  not (_07186_, _07185_);
  nor (_07187_, _07186_, _07182_);
  and (_07188_, _06877_, _06139_);
  not (_07189_, _07179_);
  and (_07190_, _07189_, _06151_);
  not (_07191_, _06151_);
  and (_07192_, _06115_, _06651_);
  not (_07193_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_07194_, _06844_, _07193_);
  not (_07195_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_07196_, _06993_, _07195_);
  and (_07197_, _07196_, _06991_);
  nand (_07198_, _07197_, _07194_);
  not (_07199_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_07200_, _06993_, _07199_);
  not (_07201_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_07202_, _06844_, _07201_);
  and (_07203_, _07202_, _06999_);
  nand (_07204_, _07203_, _07200_);
  nand (_07205_, _07204_, _07198_);
  nand (_07206_, _07205_, _06637_);
  not (_07207_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_07208_, _06993_, _07207_);
  not (_07209_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_07210_, _06844_, _07209_);
  and (_07211_, _07210_, _06999_);
  nand (_07212_, _07211_, _07208_);
  not (_07213_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_07214_, _06844_, _07213_);
  not (_07215_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_07216_, _06993_, _07215_);
  and (_07217_, _07216_, _06991_);
  nand (_07218_, _07217_, _07214_);
  nand (_07219_, _07218_, _07212_);
  nand (_07220_, _07219_, _07006_);
  nand (_07221_, _07220_, _07206_);
  nand (_07222_, _07221_, _06446_);
  not (_07223_, \oc8051_golden_model_1.IRAM[11] [1]);
  or (_07224_, _06993_, _07223_);
  not (_07225_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_07226_, _06844_, _07225_);
  and (_07227_, _07226_, _06999_);
  nand (_07228_, _07227_, _07224_);
  not (_07229_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_07230_, _06844_, _07229_);
  not (_07231_, \oc8051_golden_model_1.IRAM[9] [1]);
  or (_07232_, _06993_, _07231_);
  and (_07233_, _07232_, _06991_);
  nand (_07234_, _07233_, _07230_);
  nand (_07235_, _07234_, _07228_);
  nand (_07236_, _07235_, _06637_);
  not (_07237_, \oc8051_golden_model_1.IRAM[15] [1]);
  or (_07238_, _06993_, _07237_);
  nand (_07239_, _06993_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_07240_, _07239_, _06999_);
  nand (_07241_, _07240_, _07238_);
  not (_07242_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_07243_, _06844_, _07242_);
  not (_07244_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_07245_, _06993_, _07244_);
  and (_07246_, _07245_, _06991_);
  nand (_07247_, _07246_, _07243_);
  nand (_07248_, _07247_, _07241_);
  nand (_07249_, _07248_, _07006_);
  nand (_07250_, _07249_, _07236_);
  nand (_07251_, _07250_, _07023_);
  nand (_07252_, _07251_, _07222_);
  and (_07253_, _07252_, _06164_);
  or (_07254_, _07253_, _07192_);
  and (_07255_, _07058_, _06912_);
  nor (_07256_, _07255_, _07254_);
  and (_07257_, _07179_, _06581_);
  not (_07258_, _07257_);
  and (_07259_, _06119_, _06155_);
  nor (_07260_, _07259_, _06584_);
  and (_07261_, _07260_, _07258_);
  and (_07262_, _07261_, _07256_);
  and (_07263_, _07252_, _07064_);
  nor (_07264_, _07263_, _06162_);
  and (_07265_, _07264_, _07262_);
  and (_07266_, _06913_, _06162_);
  nor (_07267_, _07266_, _07265_);
  and (_07268_, _06876_, _06159_);
  nor (_07269_, _07268_, _07267_);
  or (_07270_, _07189_, _05764_);
  nand (_07271_, _07270_, _07269_);
  and (_07272_, _07076_, _06912_);
  and (_07273_, _06119_, _06150_);
  nor (_07274_, _07273_, _06538_);
  not (_07275_, _07274_);
  nor (_07276_, _07275_, _07272_);
  not (_07277_, _07276_);
  nor (_07278_, _07277_, _07271_);
  and (_07279_, _07252_, _07081_);
  nor (_07280_, _07279_, _07087_);
  and (_07281_, _07280_, _07278_);
  and (_07282_, _07087_, _06913_);
  nor (_07283_, _07282_, _07281_);
  and (_07284_, _06876_, _07086_);
  nor (_07285_, _07284_, _07283_);
  and (_07286_, _07285_, _07191_);
  nor (_07287_, _07286_, _07190_);
  and (_07288_, _06148_, _06876_);
  or (_07289_, _07288_, _07287_);
  nor (_07290_, _07189_, _05760_);
  and (_07291_, _05744_, _05666_);
  and (_07292_, _07291_, _06245_);
  or (_07293_, _07292_, _07290_);
  nor (_07294_, _07293_, _07289_);
  and (_07295_, _07252_, _06701_);
  nor (_07296_, _07295_, _07103_);
  and (_07297_, _07296_, _07294_);
  nor (_07298_, _07297_, _07188_);
  nor (_07299_, _07298_, _05791_);
  and (_07300_, _07189_, _05791_);
  nor (_07301_, _07300_, _07299_);
  or (_07302_, _06288_, _06123_);
  and (_07303_, _07302_, _06109_);
  nor (_07304_, _07303_, _07301_);
  and (_07305_, _07304_, _07187_);
  and (_07306_, _07251_, _07222_);
  nor (_07307_, _07306_, _07116_);
  nor (_07308_, _07307_, _06112_);
  and (_07309_, _07308_, _07305_);
  nor (_07310_, _07309_, _07181_);
  nor (_07311_, _07310_, _06076_);
  nor (_07312_, _07179_, _05836_);
  nor (_07313_, _07312_, _07311_);
  nor (_07314_, _07135_, _06913_);
  nor (_07315_, _07314_, _07124_);
  not (_07316_, _07315_);
  nor (_07317_, _07316_, _07313_);
  nor (_07318_, _07179_, _05848_);
  nor (_07319_, _07318_, _07317_);
  and (_07320_, _07143_, _06912_);
  nor (_07321_, _07320_, _07142_);
  not (_07322_, _07321_);
  nor (_07323_, _07322_, _07319_);
  nor (_07324_, _07323_, _07180_);
  and (_07325_, _06119_, _05591_);
  not (_07326_, _07325_);
  and (_07327_, _07326_, _06564_);
  not (_07328_, _07327_);
  nor (_07329_, _07328_, _07324_);
  and (_07330_, _07252_, _07153_);
  nor (_07331_, _07330_, _07152_);
  and (_07332_, _07331_, _07329_);
  and (_07333_, _07152_, _06913_);
  nor (_07334_, _07333_, _07332_);
  nor (_07335_, _07189_, _07160_);
  nor (_07336_, _07335_, _06073_);
  not (_07337_, _07336_);
  nor (_07338_, _07337_, _07334_);
  nor (_07339_, _07338_, _07176_);
  and (_07340_, _07291_, _05820_);
  nor (_07341_, _07340_, _07339_);
  and (_07342_, _07252_, _07168_);
  nor (_07343_, _07342_, _07167_);
  and (_07344_, _07343_, _07341_);
  nor (_07345_, _07344_, _07175_);
  not (_07346_, _00000_);
  nor (_07347_, _07076_, _06159_);
  nor (_07348_, _07058_, _06162_);
  and (_07349_, _07348_, _07347_);
  not (_07350_, _06112_);
  and (_07351_, _06125_, _06109_);
  not (_07352_, _07351_);
  nor (_07353_, _06972_, _06562_);
  and (_07354_, _07353_, _06531_);
  and (_07355_, _07354_, _07352_);
  nor (_07356_, _06563_, _06248_);
  not (_07357_, _06950_);
  and (_07358_, _07357_, _06540_);
  and (_07359_, _07358_, _07356_);
  and (_07360_, _05836_, _05764_);
  and (_07361_, _07360_, _06582_);
  and (_07362_, _07160_, _05850_);
  and (_07363_, _07362_, _07361_);
  and (_07364_, _07363_, _07359_);
  nor (_07365_, _06119_, _06115_);
  nor (_07366_, _07365_, _05768_);
  and (_07367_, _06249_, _05742_);
  nor (_07368_, _07367_, _07366_);
  not (_07369_, _05745_);
  and (_07370_, _06118_, _06109_);
  and (_07371_, _07370_, _07369_);
  nor (_07372_, _07365_, _05776_);
  nor (_07373_, _07372_, _07371_);
  and (_07374_, _07373_, _07368_);
  and (_07375_, _07374_, _06247_);
  and (_07376_, _07375_, _07364_);
  and (_07377_, _06122_, _06155_);
  not (_07378_, _07377_);
  and (_07379_, _06294_, _06651_);
  and (_07380_, _05786_, _06651_);
  nor (_07381_, _07380_, _07379_);
  nand (_07382_, _07381_, _05777_);
  nor (_07383_, _07382_, _07186_);
  and (_07384_, _07383_, _07378_);
  nor (_07385_, _06701_, _06151_);
  nor (_07386_, _07115_, _07064_);
  and (_07387_, _07386_, _07385_);
  not (_07388_, _05760_);
  nor (_07389_, _05791_, _07388_);
  nor (_07390_, _07168_, _07153_);
  and (_07391_, _07390_, _07389_);
  and (_07392_, _07391_, _07387_);
  not (_07393_, _06978_);
  and (_07394_, _06119_, _05820_);
  nor (_07395_, _07394_, _07259_);
  and (_07396_, _06119_, _06245_);
  nor (_07397_, _07396_, _07325_);
  and (_07398_, _07397_, _07395_);
  and (_07399_, _07398_, _07393_);
  and (_07400_, _07399_, _07392_);
  and (_07401_, _07400_, _07384_);
  and (_07402_, _07401_, _07376_);
  and (_07403_, _07402_, _07355_);
  and (_07404_, _07403_, _07350_);
  nor (_07405_, _07087_, _07086_);
  and (_07406_, _07405_, _07404_);
  and (_07407_, _07406_, _07349_);
  not (_07408_, _06135_);
  nor (_07409_, _07167_, _06073_);
  and (_07410_, _07409_, _07408_);
  nor (_07411_, _06148_, _07103_);
  nor (_07412_, _07152_, _07143_);
  and (_07413_, _07412_, _07411_);
  and (_07414_, _07413_, _07410_);
  and (_07415_, _07414_, _07135_);
  and (_07416_, _07415_, _07407_);
  nor (_07417_, _07416_, _07346_);
  not (_07418_, _07417_);
  nor (_07419_, _07418_, _07345_);
  not (_07420_, _07419_);
  nor (_07421_, _07420_, _07174_);
  not (_07422_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_07423_, _06844_, _07422_);
  not (_07424_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_07425_, _06993_, _07424_);
  and (_07426_, _07425_, _06991_);
  nand (_07427_, _07426_, _07423_);
  not (_07428_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_07429_, _06993_, _07428_);
  not (_07430_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_07431_, _06844_, _07430_);
  and (_07432_, _07431_, _06999_);
  nand (_07433_, _07432_, _07429_);
  nand (_07434_, _07433_, _07427_);
  nand (_07435_, _07434_, _06637_);
  not (_07436_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_07437_, _06993_, _07436_);
  not (_07438_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_07439_, _06844_, _07438_);
  and (_07440_, _07439_, _06999_);
  nand (_07441_, _07440_, _07437_);
  not (_07442_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_07443_, _06844_, _07442_);
  not (_07444_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_07445_, _06993_, _07444_);
  and (_07446_, _07445_, _06991_);
  nand (_07447_, _07446_, _07443_);
  nand (_07448_, _07447_, _07441_);
  nand (_07449_, _07448_, _07006_);
  nand (_07450_, _07449_, _07435_);
  nand (_07451_, _07450_, _06446_);
  nand (_07452_, _06844_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_07453_, _06993_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_07454_, _07453_, _06999_);
  nand (_07455_, _07454_, _07452_);
  nand (_07456_, _06993_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_07457_, _06844_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_07458_, _07457_, _06991_);
  nand (_07459_, _07458_, _07456_);
  nand (_07460_, _07459_, _07455_);
  nand (_07461_, _07460_, _06637_);
  nand (_07462_, _06844_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_07463_, _06993_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_07464_, _07463_, _06999_);
  nand (_07465_, _07464_, _07462_);
  nand (_07466_, _06993_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_07467_, _06844_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_07468_, _07467_, _06991_);
  nand (_07469_, _07468_, _07466_);
  nand (_07470_, _07469_, _07465_);
  nand (_07471_, _07470_, _07006_);
  nand (_07472_, _07471_, _07461_);
  nand (_07473_, _07472_, _07023_);
  nand (_07474_, _07473_, _07451_);
  and (_07475_, _07474_, _07168_);
  and (_07476_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_07477_, _07476_, \oc8051_golden_model_1.SP [2]);
  nor (_07478_, _07477_, \oc8051_golden_model_1.SP [3]);
  and (_07479_, _07477_, \oc8051_golden_model_1.SP [3]);
  nor (_07480_, _07479_, _07478_);
  and (_07481_, _07480_, _05791_);
  not (_07482_, _06203_);
  and (_07483_, _07103_, _07482_);
  and (_07484_, _07480_, _07388_);
  not (_07485_, _05764_);
  and (_07486_, _06203_, _06159_);
  and (_07487_, _07480_, _06581_);
  and (_07488_, _07474_, _06164_);
  nor (_07489_, _06164_, \oc8051_golden_model_1.PSW [3]);
  nor (_07490_, _07489_, _07058_);
  not (_07491_, _07490_);
  nor (_07492_, _07491_, _07488_);
  and (_07493_, _07058_, _06228_);
  nor (_07494_, _07493_, _07492_);
  nor (_07495_, _07494_, _06581_);
  or (_07496_, _07495_, _07064_);
  nor (_07497_, _07496_, _07487_);
  and (_07498_, _07474_, _07064_);
  nor (_07499_, _07498_, _06162_);
  not (_07500_, _07499_);
  nor (_07501_, _07500_, _07497_);
  nor (_07502_, _06161_, _06071_);
  or (_07503_, _07502_, _06159_);
  nor (_07504_, _07503_, _07501_);
  nor (_07505_, _07504_, _07486_);
  nor (_07506_, _07505_, _07485_);
  nor (_07507_, _07480_, _05764_);
  nor (_07508_, _07507_, _07076_);
  not (_07509_, _07508_);
  nor (_07510_, _07509_, _07506_);
  and (_07511_, _07076_, _06228_);
  nor (_07512_, _07511_, _07081_);
  not (_07513_, _07512_);
  nor (_07514_, _07513_, _07510_);
  and (_07515_, _07474_, _07081_);
  nor (_07516_, _07515_, _07087_);
  not (_07517_, _07516_);
  nor (_07518_, _07517_, _07514_);
  and (_07519_, _07087_, _06228_);
  or (_07520_, _07519_, _07086_);
  nor (_07521_, _07520_, _07518_);
  and (_07522_, _06203_, _07086_);
  nor (_07523_, _07522_, _07521_);
  and (_07524_, _07523_, _07191_);
  and (_07525_, _07480_, _06151_);
  nor (_07526_, _07525_, _07524_);
  nor (_07527_, _07526_, _06148_);
  nor (_07528_, _06149_, _06206_);
  or (_07529_, _07528_, _07527_);
  and (_07530_, _07529_, _05760_);
  or (_07531_, _07530_, _06701_);
  nor (_07532_, _07531_, _07484_);
  and (_07533_, _07474_, _06701_);
  nor (_07534_, _07533_, _07103_);
  not (_07535_, _07534_);
  nor (_07536_, _07535_, _07532_);
  nor (_07537_, _07536_, _07483_);
  nor (_07538_, _07537_, _05791_);
  or (_07539_, _07538_, _06135_);
  nor (_07540_, _07539_, _07481_);
  and (_07541_, _06135_, _06070_);
  or (_07542_, _07541_, _07540_);
  and (_07543_, _07542_, _07116_);
  and (_07544_, _07473_, _07451_);
  nor (_07545_, _07544_, _07116_);
  nor (_07546_, _07545_, _06112_);
  not (_07547_, _07546_);
  nor (_07548_, _07547_, _07543_);
  nor (_07549_, _06111_, _06071_);
  nor (_07550_, _07549_, _07548_);
  nor (_07551_, _07550_, _06076_);
  and (_07552_, _07480_, _06076_);
  not (_07553_, _07552_);
  and (_07554_, _07553_, _07135_);
  not (_07555_, _07554_);
  nor (_07556_, _07555_, _07551_);
  nor (_07557_, _07135_, _06228_);
  nor (_07558_, _07557_, _07124_);
  not (_07559_, _07558_);
  nor (_07560_, _07559_, _07556_);
  and (_07561_, _07480_, _07124_);
  nor (_07562_, _07561_, _07143_);
  not (_07563_, _07562_);
  nor (_07564_, _07563_, _07560_);
  and (_07565_, _07143_, _06070_);
  nor (_07566_, _07565_, _07142_);
  not (_07567_, _07566_);
  nor (_07568_, _07567_, _07564_);
  and (_07569_, _07480_, _07142_);
  nor (_07570_, _07569_, _07153_);
  not (_07571_, _07570_);
  nor (_07572_, _07571_, _07568_);
  and (_07573_, _07474_, _07153_);
  nor (_07574_, _07573_, _07152_);
  not (_07575_, _07574_);
  nor (_07576_, _07575_, _07572_);
  not (_07577_, _07160_);
  and (_07578_, _07152_, _06228_);
  nor (_07579_, _07578_, _07577_);
  not (_07580_, _07579_);
  nor (_07581_, _07580_, _07576_);
  nor (_07582_, _07480_, _07160_);
  nor (_07583_, _07582_, _06073_);
  not (_07584_, _07583_);
  nor (_07585_, _07584_, _07581_);
  and (_07586_, _06073_, _07482_);
  nor (_07587_, _07586_, _07168_);
  not (_07588_, _07587_);
  nor (_07589_, _07588_, _07585_);
  or (_07590_, _07589_, _07167_);
  nor (_07591_, _07590_, _07475_);
  and (_07592_, _07167_, _06228_);
  nor (_07593_, _07592_, _07591_);
  and (_07594_, _06478_, _05748_);
  nor (_07595_, _07476_, \oc8051_golden_model_1.SP [2]);
  nor (_07596_, _07595_, _07477_);
  not (_07597_, _07596_);
  nor (_07598_, _07597_, _05846_);
  and (_07599_, _06626_, _06112_);
  and (_07600_, _06478_, _06139_);
  and (_07601_, _07596_, _06151_);
  and (_07602_, _06626_, _06162_);
  not (_07603_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_07604_, _06844_, _07603_);
  not (_07605_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_07606_, _06993_, _07605_);
  and (_07607_, _07606_, _06991_);
  nand (_07608_, _07607_, _07604_);
  not (_07609_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_07610_, _06993_, _07609_);
  not (_07611_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_07612_, _06844_, _07611_);
  and (_07613_, _07612_, _06999_);
  nand (_07614_, _07613_, _07610_);
  nand (_07615_, _07614_, _07608_);
  nand (_07616_, _07615_, _06637_);
  not (_07617_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_07618_, _06993_, _07617_);
  not (_07619_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_07620_, _06844_, _07619_);
  and (_07621_, _07620_, _06999_);
  nand (_07622_, _07621_, _07618_);
  not (_07623_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_07624_, _06844_, _07623_);
  not (_07625_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_07626_, _06993_, _07625_);
  and (_07627_, _07626_, _06991_);
  nand (_07628_, _07627_, _07624_);
  nand (_07629_, _07628_, _07622_);
  nand (_07630_, _07629_, _07006_);
  nand (_07631_, _07630_, _07616_);
  nand (_07632_, _07631_, _06446_);
  not (_07633_, \oc8051_golden_model_1.IRAM[11] [2]);
  or (_07634_, _06993_, _07633_);
  not (_07635_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_07636_, _06844_, _07635_);
  and (_07637_, _07636_, _06999_);
  nand (_07638_, _07637_, _07634_);
  nand (_07639_, _06993_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_07640_, _06844_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_07641_, _07640_, _06991_);
  nand (_07642_, _07641_, _07639_);
  nand (_07643_, _07642_, _07638_);
  nand (_07644_, _07643_, _06637_);
  nand (_07645_, _06844_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_07646_, _06993_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_07647_, _07646_, _06999_);
  nand (_07648_, _07647_, _07645_);
  nand (_07649_, _06993_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_07650_, _06844_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_07651_, _07650_, _06991_);
  nand (_07652_, _07651_, _07649_);
  nand (_07653_, _07652_, _07648_);
  nand (_07654_, _07653_, _07006_);
  nand (_07655_, _07654_, _07644_);
  nand (_07656_, _07655_, _07023_);
  nand (_07657_, _07656_, _07632_);
  or (_07658_, _07657_, _05752_);
  and (_07659_, _07658_, _07382_);
  and (_07660_, _07058_, _06625_);
  nor (_07661_, _07660_, _07659_);
  and (_07662_, _07597_, _06581_);
  not (_07663_, _07662_);
  and (_07664_, _06273_, _06155_);
  and (_07665_, _06288_, _06155_);
  or (_07666_, _07665_, _06978_);
  nor (_07667_, _07666_, _07664_);
  and (_07668_, _07667_, _07663_);
  and (_07669_, _07668_, _07661_);
  and (_07670_, _07657_, _07064_);
  nor (_07671_, _07670_, _06162_);
  and (_07672_, _07671_, _07669_);
  nor (_07673_, _07672_, _07602_);
  nor (_07674_, _07673_, _06159_);
  nor (_07675_, _07674_, _06489_);
  nor (_07676_, _07596_, _05764_);
  nor (_07677_, _07676_, _07675_);
  and (_07678_, _06118_, _06150_);
  and (_07679_, _07076_, _06625_);
  nor (_07680_, _07679_, _07678_);
  and (_07681_, _07680_, _07677_);
  and (_07682_, _07657_, _07081_);
  nor (_07683_, _07682_, _07087_);
  and (_07684_, _07683_, _07681_);
  and (_07685_, _07087_, _06626_);
  nor (_07686_, _07685_, _07684_);
  and (_07687_, _06477_, _07086_);
  nor (_07688_, _07687_, _07686_);
  and (_07689_, _07688_, _07191_);
  nor (_07690_, _07689_, _07601_);
  and (_07691_, _06148_, _06477_);
  or (_07692_, _07691_, _07690_);
  nor (_07693_, _07596_, _05760_);
  nor (_07694_, _07693_, _06249_);
  not (_07695_, _07694_);
  nor (_07696_, _07695_, _07692_);
  and (_07697_, _07657_, _06701_);
  nor (_07698_, _07697_, _07103_);
  and (_07699_, _07698_, _07696_);
  nor (_07700_, _07699_, _07600_);
  nor (_07701_, _07700_, _05791_);
  and (_07702_, _07596_, _05791_);
  nor (_07703_, _07702_, _07701_);
  and (_07704_, _06135_, _06625_);
  nor (_07705_, _07704_, _07370_);
  not (_07706_, _07705_);
  nor (_07707_, _07706_, _07703_);
  and (_07708_, _07656_, _07632_);
  nor (_07709_, _07708_, _07116_);
  nor (_07710_, _07709_, _06112_);
  and (_07711_, _07710_, _07707_);
  nor (_07712_, _07711_, _07599_);
  nor (_07713_, _07712_, _06076_);
  nor (_07714_, _07597_, _05836_);
  nor (_07715_, _07714_, _07713_);
  nor (_07716_, _07135_, _06626_);
  nor (_07717_, _07716_, _07124_);
  not (_07718_, _07717_);
  nor (_07719_, _07718_, _07715_);
  nor (_07720_, _07597_, _05848_);
  nor (_07721_, _07720_, _07719_);
  and (_07722_, _07143_, _06625_);
  nor (_07723_, _07722_, _07142_);
  not (_07724_, _07723_);
  nor (_07725_, _07724_, _07721_);
  nor (_07726_, _07725_, _07598_);
  nor (_07727_, _07325_, _06972_);
  not (_07728_, _07727_);
  nor (_07729_, _07728_, _07726_);
  and (_07730_, _07657_, _07153_);
  nor (_07731_, _07730_, _07152_);
  and (_07732_, _07731_, _07729_);
  and (_07733_, _07152_, _06626_);
  nor (_07734_, _07733_, _07732_);
  nor (_07735_, _07596_, _07160_);
  nor (_07736_, _07735_, _06073_);
  not (_07737_, _07736_);
  nor (_07738_, _07737_, _07734_);
  nor (_07739_, _07738_, _07594_);
  and (_07740_, _06118_, _05820_);
  nor (_07741_, _07740_, _07739_);
  and (_07742_, _07657_, _07168_);
  nor (_07743_, _07742_, _07167_);
  and (_07744_, _07743_, _07741_);
  and (_07745_, _07167_, _06626_);
  nor (_07746_, _07745_, _07744_);
  nor (_07747_, _07746_, _07418_);
  not (_07748_, _07747_);
  nor (_07749_, _07748_, _07593_);
  and (_07750_, _07749_, _07421_);
  or (_07751_, _07750_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_07752_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_07753_, _07752_, _06142_);
  nor (_07754_, _07596_, _07178_);
  nor (_07755_, _07754_, _07753_);
  and (_07756_, _07752_, \oc8051_golden_model_1.SP [3]);
  and (_07757_, _07756_, _06142_);
  nor (_07758_, _07753_, _07480_);
  nor (_07759_, _07758_, _07757_);
  and (_07760_, _07389_, _07360_);
  and (_07761_, _07160_, _06582_);
  and (_07762_, _07761_, _05850_);
  and (_07763_, _07762_, _07760_);
  nor (_07764_, _07763_, _07346_);
  and (_07765_, _07764_, _07759_);
  and (_07766_, _07765_, _07755_);
  and (_07767_, _07766_, _07177_);
  not (_07768_, _07767_);
  and (_07769_, _07768_, _07751_);
  not (_07770_, _07750_);
  and (_07771_, _06912_, _06107_);
  and (_07772_, _07771_, _06625_);
  and (_07773_, _07772_, _06228_);
  and (_07774_, _06203_, _06039_);
  not (_07775_, _06876_);
  and (_07776_, _07775_, _06477_);
  and (_07777_, _07776_, _07774_);
  and (_07778_, _07777_, _07773_);
  and (_07779_, _07778_, \oc8051_golden_model_1.SCON [7]);
  and (_07780_, _06912_, _06108_);
  and (_07781_, _07780_, _06625_);
  and (_07782_, _07781_, _06228_);
  and (_07783_, _07782_, _07777_);
  and (_07784_, _07783_, \oc8051_golden_model_1.SBUF [7]);
  or (_07785_, _07784_, _07779_);
  and (_07786_, _07774_, _06477_);
  and (_07787_, _07786_, _06876_);
  and (_07788_, _07787_, _07773_);
  and (_07789_, _07788_, \oc8051_golden_model_1.TCON [7]);
  nand (_07790_, _07772_, _06070_);
  nor (_07791_, _06203_, _06172_);
  and (_07792_, _07791_, _07776_);
  not (_07793_, _07792_);
  nor (_07794_, _07793_, _07790_);
  and (_07795_, _07794_, \oc8051_golden_model_1.PSW [7]);
  or (_07796_, _07795_, _07789_);
  or (_07797_, _07796_, _07785_);
  not (_07798_, _07787_);
  nand (_07799_, _06625_, _06228_);
  nor (_07800_, _06912_, _06108_);
  not (_07801_, _07800_);
  or (_07802_, _07801_, _07799_);
  nor (_07803_, _07802_, _07798_);
  and (_07804_, _07803_, \oc8051_golden_model_1.TL0 [7]);
  not (_07805_, _06477_);
  and (_07806_, _06876_, _07805_);
  and (_07807_, _07806_, _07791_);
  not (_07808_, _07807_);
  nor (_07809_, _07808_, _07790_);
  and (_07810_, _07809_, \oc8051_golden_model_1.ACC [7]);
  or (_07811_, _07810_, _07804_);
  and (_07812_, _07787_, _07782_);
  and (_07813_, _07812_, \oc8051_golden_model_1.TMOD [7]);
  not (_07814_, _07780_);
  or (_07815_, _06625_, _06070_);
  or (_07816_, _07815_, _07814_);
  nor (_07817_, _07816_, _07798_);
  and (_07818_, _07817_, \oc8051_golden_model_1.TH1 [7]);
  or (_07819_, _07818_, _07813_);
  or (_07820_, _07819_, _07811_);
  not (_07821_, _07771_);
  or (_07822_, _07815_, _07821_);
  nor (_07823_, _07822_, _07798_);
  and (_07824_, _07823_, \oc8051_golden_model_1.TH0 [7]);
  and (_07825_, _07806_, _07774_);
  and (_07826_, _07825_, _07773_);
  and (_07827_, _07826_, \oc8051_golden_model_1.IE [7]);
  nor (_07828_, _06876_, _06477_);
  and (_07829_, _07828_, _07774_);
  and (_07830_, _07829_, _07773_);
  and (_07831_, _07830_, \oc8051_golden_model_1.IP [7]);
  or (_07832_, _07831_, _07827_);
  or (_07833_, _07832_, _07824_);
  nor (_07834_, _06912_, _06107_);
  not (_07835_, _07834_);
  or (_07836_, _07835_, _07799_);
  nor (_07837_, _07836_, _07798_);
  and (_07838_, _07837_, \oc8051_golden_model_1.TL1 [7]);
  and (_07839_, _07828_, _07791_);
  not (_07840_, _07839_);
  nor (_07841_, _07840_, _07790_);
  and (_07842_, _07841_, \oc8051_golden_model_1.B [7]);
  or (_07843_, _07842_, _07838_);
  or (_07844_, _07843_, _07833_);
  or (_07845_, _07844_, _07820_);
  or (_07846_, _07845_, _07797_);
  and (_07847_, _07787_, _06070_);
  and (_07848_, _07800_, _06625_);
  and (_07849_, _07848_, _07847_);
  and (_07850_, _07849_, \oc8051_golden_model_1.DPL [7]);
  and (_07851_, _07834_, _06625_);
  and (_07852_, _07851_, _07847_);
  and (_07853_, _07852_, \oc8051_golden_model_1.DPH [7]);
  or (_07854_, _07853_, _07850_);
  and (_07855_, _07834_, _06626_);
  and (_07856_, _07855_, _07847_);
  and (_07857_, _07856_, \oc8051_golden_model_1.PCON [7]);
  and (_07858_, _07847_, _07781_);
  and (_07859_, _07858_, \oc8051_golden_model_1.SP [7]);
  or (_07860_, _07859_, _07857_);
  or (_07861_, _07860_, _07854_);
  or (_07862_, _07861_, _07846_);
  not (_07863_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_07864_, _06844_, _07863_);
  not (_07865_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_07866_, _06993_, _07865_);
  and (_07867_, _07866_, _06991_);
  nand (_07868_, _07867_, _07864_);
  not (_07869_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_07870_, _06993_, _07869_);
  not (_07871_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_07872_, _06844_, _07871_);
  and (_07873_, _07872_, _06999_);
  nand (_07874_, _07873_, _07870_);
  nand (_07875_, _07874_, _07868_);
  nand (_07876_, _07875_, _06637_);
  not (_07877_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_07878_, _06993_, _07877_);
  not (_07879_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_07880_, _06844_, _07879_);
  and (_07881_, _07880_, _06999_);
  nand (_07882_, _07881_, _07878_);
  not (_07883_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_07884_, _06844_, _07883_);
  not (_07885_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_07886_, _06993_, _07885_);
  and (_07887_, _07886_, _06991_);
  nand (_07888_, _07887_, _07884_);
  nand (_07889_, _07888_, _07882_);
  nand (_07890_, _07889_, _07006_);
  nand (_07891_, _07890_, _07876_);
  nand (_07892_, _07891_, _06446_);
  not (_07893_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_07894_, _06993_, _07893_);
  not (_07895_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_07896_, _06844_, _07895_);
  and (_07897_, _07896_, _06999_);
  nand (_07898_, _07897_, _07894_);
  not (_07899_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_07900_, _06844_, _07899_);
  not (_07901_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_07902_, _06993_, _07901_);
  and (_07903_, _07902_, _06991_);
  nand (_07904_, _07903_, _07900_);
  nand (_07905_, _07904_, _07898_);
  nand (_07906_, _07905_, _06637_);
  not (_07907_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_07908_, _06993_, _07907_);
  not (_07909_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_07910_, _06844_, _07909_);
  and (_07911_, _07910_, _06999_);
  nand (_07912_, _07911_, _07908_);
  not (_07913_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_07914_, _06844_, _07913_);
  not (_07915_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_07916_, _06993_, _07915_);
  and (_07917_, _07916_, _06991_);
  nand (_07918_, _07917_, _07914_);
  nand (_07919_, _07918_, _07912_);
  nand (_07920_, _07919_, _07006_);
  nand (_07921_, _07920_, _07906_);
  nand (_07922_, _07921_, _07023_);
  and (_07923_, _07922_, _07892_);
  and (_07924_, _07923_, _06172_);
  nor (_07925_, _07924_, _07862_);
  not (_07926_, _07925_);
  and (_07927_, _07837_, \oc8051_golden_model_1.TL1 [6]);
  and (_07928_, _07817_, \oc8051_golden_model_1.TH1 [6]);
  or (_07929_, _07928_, _07927_);
  and (_07930_, _07788_, \oc8051_golden_model_1.TCON [6]);
  and (_07931_, _07812_, \oc8051_golden_model_1.TMOD [6]);
  or (_07932_, _07931_, _07930_);
  or (_07933_, _07932_, _07929_);
  and (_07934_, _07803_, \oc8051_golden_model_1.TL0 [6]);
  and (_07935_, _07778_, \oc8051_golden_model_1.SCON [6]);
  or (_07936_, _07935_, _07934_);
  and (_07937_, _07823_, \oc8051_golden_model_1.TH0 [6]);
  and (_07938_, _07794_, \oc8051_golden_model_1.PSW [6]);
  or (_07939_, _07938_, _07937_);
  or (_07940_, _07939_, _07936_);
  and (_07941_, _07841_, \oc8051_golden_model_1.B [6]);
  and (_07942_, _07826_, \oc8051_golden_model_1.IE [6]);
  and (_07943_, _07830_, \oc8051_golden_model_1.IP [6]);
  or (_07944_, _07943_, _07942_);
  or (_07945_, _07944_, _07941_);
  and (_07946_, _07783_, \oc8051_golden_model_1.SBUF [6]);
  and (_07947_, _07809_, \oc8051_golden_model_1.ACC [6]);
  or (_07948_, _07947_, _07946_);
  or (_07949_, _07948_, _07945_);
  or (_07950_, _07949_, _07940_);
  or (_07951_, _07950_, _07933_);
  and (_07952_, _07856_, \oc8051_golden_model_1.PCON [6]);
  and (_07953_, _07852_, \oc8051_golden_model_1.DPH [6]);
  or (_07954_, _07953_, _07952_);
  and (_07955_, _07849_, \oc8051_golden_model_1.DPL [6]);
  and (_07956_, _07858_, \oc8051_golden_model_1.SP [6]);
  or (_07957_, _07956_, _07955_);
  or (_07958_, _07957_, _07954_);
  or (_07959_, _07958_, _07951_);
  not (_07960_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_07961_, _06844_, _07960_);
  not (_07962_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_07963_, _06993_, _07962_);
  and (_07964_, _07963_, _06991_);
  nand (_07965_, _07964_, _07961_);
  not (_07966_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_07967_, _06993_, _07966_);
  not (_07968_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_07969_, _06844_, _07968_);
  and (_07970_, _07969_, _06999_);
  nand (_07971_, _07970_, _07967_);
  nand (_07972_, _07971_, _07965_);
  nand (_07973_, _07972_, _06637_);
  not (_07974_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_07975_, _06993_, _07974_);
  not (_07976_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_07977_, _06844_, _07976_);
  and (_07978_, _07977_, _06999_);
  nand (_07979_, _07978_, _07975_);
  not (_07980_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_07981_, _06844_, _07980_);
  not (_07982_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_07983_, _06993_, _07982_);
  and (_07984_, _07983_, _06991_);
  nand (_07985_, _07984_, _07981_);
  nand (_07986_, _07985_, _07979_);
  nand (_07987_, _07986_, _07006_);
  nand (_07988_, _07987_, _07973_);
  nand (_07989_, _07988_, _06446_);
  nand (_07990_, _06844_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_07991_, _06993_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_07992_, _07991_, _06999_);
  nand (_07993_, _07992_, _07990_);
  nand (_07994_, _06993_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_07995_, _06844_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_07996_, _07995_, _06991_);
  nand (_07997_, _07996_, _07994_);
  nand (_07998_, _07997_, _07993_);
  nand (_07999_, _07998_, _06637_);
  nand (_08000_, _06844_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_08001_, _06993_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_08002_, _08001_, _06999_);
  nand (_08003_, _08002_, _08000_);
  nand (_08004_, _06993_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_08005_, _06844_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_08006_, _08005_, _06991_);
  nand (_08007_, _08006_, _08004_);
  nand (_08008_, _08007_, _08003_);
  nand (_08009_, _08008_, _07006_);
  nand (_08010_, _08009_, _07999_);
  nand (_08011_, _08010_, _07023_);
  and (_08012_, _08011_, _07989_);
  and (_08013_, _08012_, _06172_);
  nor (_08014_, _08013_, _07959_);
  not (_08015_, _08014_);
  and (_08016_, _07788_, \oc8051_golden_model_1.TCON [5]);
  and (_08017_, _07812_, \oc8051_golden_model_1.TMOD [5]);
  or (_08018_, _08017_, _08016_);
  and (_08019_, _07778_, \oc8051_golden_model_1.SCON [5]);
  and (_08020_, _07794_, \oc8051_golden_model_1.PSW [5]);
  or (_08021_, _08020_, _08019_);
  or (_08022_, _08021_, _08018_);
  and (_08023_, _07817_, \oc8051_golden_model_1.TH1 [5]);
  and (_08024_, _07783_, \oc8051_golden_model_1.SBUF [5]);
  or (_08025_, _08024_, _08023_);
  and (_08026_, _07803_, \oc8051_golden_model_1.TL0 [5]);
  and (_08027_, _07837_, \oc8051_golden_model_1.TL1 [5]);
  or (_08028_, _08027_, _08026_);
  or (_08029_, _08028_, _08025_);
  and (_08030_, _07841_, \oc8051_golden_model_1.B [5]);
  and (_08031_, _07826_, \oc8051_golden_model_1.IE [5]);
  and (_08032_, _07830_, \oc8051_golden_model_1.IP [5]);
  or (_08033_, _08032_, _08031_);
  or (_08034_, _08033_, _08030_);
  and (_08035_, _07823_, \oc8051_golden_model_1.TH0 [5]);
  and (_08036_, _07809_, \oc8051_golden_model_1.ACC [5]);
  or (_08037_, _08036_, _08035_);
  or (_08038_, _08037_, _08034_);
  or (_08039_, _08038_, _08029_);
  or (_08040_, _08039_, _08022_);
  and (_08041_, _07849_, \oc8051_golden_model_1.DPL [5]);
  and (_08042_, _07852_, \oc8051_golden_model_1.DPH [5]);
  or (_08043_, _08042_, _08041_);
  and (_08044_, _07856_, \oc8051_golden_model_1.PCON [5]);
  and (_08045_, _07858_, \oc8051_golden_model_1.SP [5]);
  or (_08046_, _08045_, _08044_);
  or (_08047_, _08046_, _08043_);
  or (_08048_, _08047_, _08040_);
  not (_08049_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_08050_, _06844_, _08049_);
  not (_08051_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_08052_, _06993_, _08051_);
  and (_08053_, _08052_, _06991_);
  nand (_08054_, _08053_, _08050_);
  not (_08055_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_08056_, _06993_, _08055_);
  not (_08057_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_08058_, _06844_, _08057_);
  and (_08059_, _08058_, _06999_);
  nand (_08060_, _08059_, _08056_);
  nand (_08061_, _08060_, _08054_);
  nand (_08062_, _08061_, _06637_);
  not (_08063_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_08064_, _06993_, _08063_);
  not (_08065_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_08066_, _06844_, _08065_);
  and (_08067_, _08066_, _06999_);
  nand (_08068_, _08067_, _08064_);
  not (_08069_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_08070_, _06844_, _08069_);
  not (_08071_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_08072_, _06993_, _08071_);
  and (_08073_, _08072_, _06991_);
  nand (_08074_, _08073_, _08070_);
  nand (_08075_, _08074_, _08068_);
  nand (_08076_, _08075_, _07006_);
  nand (_08077_, _08076_, _08062_);
  nand (_08078_, _08077_, _06446_);
  nand (_08079_, _06844_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_08080_, _06993_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_08081_, _08080_, _06999_);
  nand (_08082_, _08081_, _08079_);
  nand (_08083_, _06993_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_08084_, _06844_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_08085_, _08084_, _06991_);
  nand (_08086_, _08085_, _08083_);
  nand (_08087_, _08086_, _08082_);
  nand (_08088_, _08087_, _06637_);
  nand (_08089_, _06844_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_08090_, _06993_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_08091_, _08090_, _06999_);
  nand (_08092_, _08091_, _08089_);
  nand (_08093_, _06993_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand (_08094_, _06844_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_08095_, _08094_, _06991_);
  nand (_08096_, _08095_, _08093_);
  nand (_08097_, _08096_, _08092_);
  nand (_08098_, _08097_, _07006_);
  nand (_08099_, _08098_, _08088_);
  nand (_08100_, _08099_, _07023_);
  and (_08101_, _08100_, _08078_);
  and (_08102_, _08101_, _06172_);
  nor (_08103_, _08102_, _08048_);
  not (_08104_, _08103_);
  and (_08105_, _07788_, \oc8051_golden_model_1.TCON [3]);
  and (_08106_, _07812_, \oc8051_golden_model_1.TMOD [3]);
  or (_08107_, _08106_, _08105_);
  and (_08108_, _07778_, \oc8051_golden_model_1.SCON [3]);
  and (_08109_, _07794_, \oc8051_golden_model_1.PSW [3]);
  or (_08110_, _08109_, _08108_);
  or (_08111_, _08110_, _08107_);
  and (_08112_, _07823_, \oc8051_golden_model_1.TH0 [3]);
  and (_08113_, _07837_, \oc8051_golden_model_1.TL1 [3]);
  or (_08114_, _08113_, _08112_);
  and (_08115_, _07803_, \oc8051_golden_model_1.TL0 [3]);
  and (_08116_, _07817_, \oc8051_golden_model_1.TH1 [3]);
  or (_08117_, _08116_, _08115_);
  or (_08118_, _08117_, _08114_);
  and (_08119_, _07841_, \oc8051_golden_model_1.B [3]);
  and (_08120_, _07826_, \oc8051_golden_model_1.IE [3]);
  and (_08121_, _07830_, \oc8051_golden_model_1.IP [3]);
  or (_08122_, _08121_, _08120_);
  or (_08123_, _08122_, _08119_);
  and (_08124_, _07783_, \oc8051_golden_model_1.SBUF [3]);
  and (_08125_, _07809_, \oc8051_golden_model_1.ACC [3]);
  or (_08126_, _08125_, _08124_);
  or (_08127_, _08126_, _08123_);
  or (_08128_, _08127_, _08118_);
  or (_08129_, _08128_, _08111_);
  and (_08130_, _07856_, \oc8051_golden_model_1.PCON [3]);
  and (_08131_, _07858_, \oc8051_golden_model_1.SP [3]);
  or (_08132_, _08131_, _08130_);
  and (_08133_, _07849_, \oc8051_golden_model_1.DPL [3]);
  and (_08134_, _07852_, \oc8051_golden_model_1.DPH [3]);
  or (_08135_, _08134_, _08133_);
  or (_08136_, _08135_, _08132_);
  or (_08137_, _08136_, _08129_);
  and (_08138_, _07544_, _06172_);
  nor (_08139_, _08138_, _08137_);
  not (_08140_, _08139_);
  and (_08141_, _07778_, \oc8051_golden_model_1.SCON [1]);
  and (_08142_, _07783_, \oc8051_golden_model_1.SBUF [1]);
  or (_08143_, _08142_, _08141_);
  and (_08144_, _07788_, \oc8051_golden_model_1.TCON [1]);
  and (_08145_, _07794_, \oc8051_golden_model_1.PSW [1]);
  or (_08146_, _08145_, _08144_);
  or (_08147_, _08146_, _08143_);
  and (_08148_, _07841_, \oc8051_golden_model_1.B [1]);
  and (_08149_, _07809_, \oc8051_golden_model_1.ACC [1]);
  or (_08150_, _08149_, _08148_);
  and (_08151_, _07823_, \oc8051_golden_model_1.TH0 [1]);
  and (_08152_, _07837_, \oc8051_golden_model_1.TL1 [1]);
  or (_08153_, _08152_, _08151_);
  or (_08154_, _08153_, _08150_);
  and (_08155_, _07817_, \oc8051_golden_model_1.TH1 [1]);
  and (_08156_, _07826_, \oc8051_golden_model_1.IE [1]);
  and (_08157_, _07830_, \oc8051_golden_model_1.IP [1]);
  or (_08158_, _08157_, _08156_);
  or (_08159_, _08158_, _08155_);
  and (_08160_, _07812_, \oc8051_golden_model_1.TMOD [1]);
  and (_08161_, _07803_, \oc8051_golden_model_1.TL0 [1]);
  or (_08162_, _08161_, _08160_);
  or (_08163_, _08162_, _08159_);
  or (_08164_, _08163_, _08154_);
  or (_08165_, _08164_, _08147_);
  and (_08166_, _07858_, \oc8051_golden_model_1.SP [1]);
  and (_08167_, _07852_, \oc8051_golden_model_1.DPH [1]);
  or (_08168_, _08167_, _08166_);
  and (_08169_, _07849_, \oc8051_golden_model_1.DPL [1]);
  and (_08170_, _07856_, \oc8051_golden_model_1.PCON [1]);
  or (_08171_, _08170_, _08169_);
  or (_08172_, _08171_, _08168_);
  or (_08173_, _08172_, _08165_);
  and (_08174_, _07306_, _06172_);
  nor (_08175_, _08174_, _08173_);
  not (_08176_, _08175_);
  and (_08177_, _07788_, \oc8051_golden_model_1.TCON [0]);
  and (_08178_, _07778_, \oc8051_golden_model_1.SCON [0]);
  or (_08179_, _08178_, _08177_);
  and (_08180_, _07783_, \oc8051_golden_model_1.SBUF [0]);
  and (_08181_, _07809_, \oc8051_golden_model_1.ACC [0]);
  or (_08182_, _08181_, _08180_);
  or (_08183_, _08182_, _08179_);
  and (_08184_, _07812_, \oc8051_golden_model_1.TMOD [0]);
  and (_08185_, _07803_, \oc8051_golden_model_1.TL0 [0]);
  or (_08186_, _08185_, _08184_);
  and (_08187_, _07823_, \oc8051_golden_model_1.TH0 [0]);
  and (_08188_, _07837_, \oc8051_golden_model_1.TL1 [0]);
  or (_08189_, _08188_, _08187_);
  or (_08190_, _08189_, _08186_);
  and (_08191_, _07794_, \oc8051_golden_model_1.PSW [0]);
  and (_08192_, _07826_, \oc8051_golden_model_1.IE [0]);
  and (_08193_, _07830_, \oc8051_golden_model_1.IP [0]);
  or (_08194_, _08193_, _08192_);
  or (_08195_, _08194_, _08191_);
  and (_08196_, _07817_, \oc8051_golden_model_1.TH1 [0]);
  and (_08197_, _07841_, \oc8051_golden_model_1.B [0]);
  or (_08198_, _08197_, _08196_);
  or (_08199_, _08198_, _08195_);
  or (_08200_, _08199_, _08190_);
  or (_08201_, _08200_, _08183_);
  and (_08202_, _07849_, \oc8051_golden_model_1.DPL [0]);
  and (_08203_, _07852_, \oc8051_golden_model_1.DPH [0]);
  or (_08204_, _08203_, _08202_);
  and (_08205_, _07856_, \oc8051_golden_model_1.PCON [0]);
  and (_08206_, _07858_, \oc8051_golden_model_1.SP [0]);
  or (_08207_, _08206_, _08205_);
  or (_08208_, _08207_, _08204_);
  or (_08209_, _08208_, _08201_);
  and (_08210_, _07049_, _06172_);
  or (_08211_, _08210_, _08209_);
  and (_08212_, _08211_, _08176_);
  and (_08213_, _07837_, \oc8051_golden_model_1.TL1 [2]);
  and (_08214_, _07817_, \oc8051_golden_model_1.TH1 [2]);
  or (_08215_, _08214_, _08213_);
  and (_08216_, _07788_, \oc8051_golden_model_1.TCON [2]);
  and (_08217_, _07812_, \oc8051_golden_model_1.TMOD [2]);
  or (_08218_, _08217_, _08216_);
  or (_08219_, _08218_, _08215_);
  and (_08220_, _07803_, \oc8051_golden_model_1.TL0 [2]);
  and (_08221_, _07809_, \oc8051_golden_model_1.ACC [2]);
  or (_08222_, _08221_, _08220_);
  and (_08223_, _07823_, \oc8051_golden_model_1.TH0 [2]);
  and (_08224_, _07841_, \oc8051_golden_model_1.B [2]);
  or (_08225_, _08224_, _08223_);
  or (_08226_, _08225_, _08222_);
  and (_08227_, _07783_, \oc8051_golden_model_1.SBUF [2]);
  and (_08228_, _07826_, \oc8051_golden_model_1.IE [2]);
  and (_08229_, _07830_, \oc8051_golden_model_1.IP [2]);
  or (_08230_, _08229_, _08228_);
  or (_08231_, _08230_, _08227_);
  and (_08232_, _07778_, \oc8051_golden_model_1.SCON [2]);
  and (_08233_, _07794_, \oc8051_golden_model_1.PSW [2]);
  or (_08234_, _08233_, _08232_);
  or (_08235_, _08234_, _08231_);
  or (_08236_, _08235_, _08226_);
  or (_08237_, _08236_, _08219_);
  and (_08238_, _07849_, \oc8051_golden_model_1.DPL [2]);
  and (_08239_, _07852_, \oc8051_golden_model_1.DPH [2]);
  or (_08240_, _08239_, _08238_);
  and (_08241_, _07856_, \oc8051_golden_model_1.PCON [2]);
  and (_08242_, _07858_, \oc8051_golden_model_1.SP [2]);
  or (_08243_, _08242_, _08241_);
  or (_08244_, _08243_, _08240_);
  or (_08245_, _08244_, _08237_);
  and (_08246_, _07708_, _06172_);
  nor (_08247_, _08246_, _08245_);
  not (_08248_, _08247_);
  and (_08249_, _08248_, _08212_);
  and (_08250_, _08249_, _08140_);
  and (_08251_, _07788_, \oc8051_golden_model_1.TCON [4]);
  and (_08252_, _07778_, \oc8051_golden_model_1.SCON [4]);
  or (_08253_, _08252_, _08251_);
  and (_08254_, _07794_, \oc8051_golden_model_1.PSW [4]);
  and (_08255_, _07809_, \oc8051_golden_model_1.ACC [4]);
  or (_08256_, _08255_, _08254_);
  or (_08257_, _08256_, _08253_);
  and (_08258_, _07812_, \oc8051_golden_model_1.TMOD [4]);
  and (_08259_, _07803_, \oc8051_golden_model_1.TL0 [4]);
  or (_08260_, _08259_, _08258_);
  and (_08261_, _07823_, \oc8051_golden_model_1.TH0 [4]);
  and (_08262_, _07837_, \oc8051_golden_model_1.TL1 [4]);
  or (_08263_, _08262_, _08261_);
  or (_08264_, _08263_, _08260_);
  and (_08265_, _07783_, \oc8051_golden_model_1.SBUF [4]);
  and (_08266_, _07826_, \oc8051_golden_model_1.IE [4]);
  and (_08267_, _07830_, \oc8051_golden_model_1.IP [4]);
  or (_08268_, _08267_, _08266_);
  or (_08269_, _08268_, _08265_);
  and (_08270_, _07817_, \oc8051_golden_model_1.TH1 [4]);
  and (_08271_, _07841_, \oc8051_golden_model_1.B [4]);
  or (_08272_, _08271_, _08270_);
  or (_08273_, _08272_, _08269_);
  or (_08274_, _08273_, _08264_);
  or (_08275_, _08274_, _08257_);
  and (_08276_, _07849_, \oc8051_golden_model_1.DPL [4]);
  and (_08277_, _07852_, \oc8051_golden_model_1.DPH [4]);
  or (_08278_, _08277_, _08276_);
  and (_08279_, _07856_, \oc8051_golden_model_1.PCON [4]);
  and (_08280_, _07858_, \oc8051_golden_model_1.SP [4]);
  or (_08281_, _08280_, _08279_);
  or (_08282_, _08281_, _08278_);
  or (_08283_, _08282_, _08275_);
  not (_08284_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_08285_, _06844_, _08284_);
  not (_08286_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_08287_, _06993_, _08286_);
  and (_08288_, _08287_, _06991_);
  nand (_08289_, _08288_, _08285_);
  not (_08290_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_08291_, _06993_, _08290_);
  not (_08292_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_08293_, _06844_, _08292_);
  and (_08294_, _08293_, _06999_);
  nand (_08295_, _08294_, _08291_);
  nand (_08296_, _08295_, _08289_);
  nand (_08297_, _08296_, _06637_);
  not (_08298_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_08299_, _06993_, _08298_);
  not (_08300_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_08301_, _06844_, _08300_);
  and (_08302_, _08301_, _06999_);
  nand (_08303_, _08302_, _08299_);
  not (_08304_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_08305_, _06844_, _08304_);
  not (_08306_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_08307_, _06993_, _08306_);
  and (_08308_, _08307_, _06991_);
  nand (_08309_, _08308_, _08305_);
  nand (_08310_, _08309_, _08303_);
  nand (_08311_, _08310_, _07006_);
  nand (_08312_, _08311_, _08297_);
  nand (_08313_, _08312_, _06446_);
  nand (_08314_, _06844_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_08315_, _06993_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_08316_, _08315_, _06999_);
  nand (_08317_, _08316_, _08314_);
  nand (_08318_, _06993_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_08319_, _06844_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_08320_, _08319_, _06991_);
  nand (_08321_, _08320_, _08318_);
  nand (_08322_, _08321_, _08317_);
  nand (_08323_, _08322_, _06637_);
  nand (_08324_, _06844_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_08325_, _06993_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_08326_, _08325_, _06999_);
  nand (_08327_, _08326_, _08324_);
  nand (_08328_, _06993_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand (_08329_, _06844_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_08330_, _08329_, _06991_);
  nand (_08331_, _08330_, _08328_);
  nand (_08332_, _08331_, _08327_);
  nand (_08333_, _08332_, _07006_);
  nand (_08334_, _08333_, _08323_);
  nand (_08335_, _08334_, _07023_);
  and (_08336_, _08335_, _08313_);
  and (_08337_, _08336_, _06172_);
  nor (_08338_, _08337_, _08283_);
  not (_08339_, _08338_);
  and (_08340_, _08339_, _08250_);
  and (_08341_, _08340_, _08104_);
  and (_08342_, _08341_, _08015_);
  nor (_08343_, _08342_, _07926_);
  and (_08344_, _08342_, _07926_);
  nor (_08345_, _08344_, _08343_);
  and (_08346_, _08345_, _07167_);
  nand (_08347_, _08011_, _07989_);
  nand (_08348_, _08100_, _08078_);
  nand (_08349_, _08335_, _08313_);
  and (_08350_, _08349_, _08348_);
  and (_08351_, _07657_, _07474_);
  nor (_08352_, _07306_, _07049_);
  and (_08353_, _08352_, _08351_);
  and (_08354_, _08353_, _08350_);
  and (_08355_, _08354_, _08347_);
  or (_08356_, _08355_, _07923_);
  nand (_08357_, _08355_, _07923_);
  and (_08358_, _08357_, _08356_);
  and (_08359_, _06125_, _05591_);
  not (_08360_, _08359_);
  and (_08361_, _08360_, _07353_);
  and (_08362_, _08361_, _07326_);
  or (_08363_, _08362_, _08358_);
  not (_08364_, _07131_);
  and (_08365_, _06366_, _04273_);
  and (_08366_, _06368_, _04246_);
  nor (_08367_, _08366_, _08365_);
  and (_08368_, _06377_, _04270_);
  and (_08369_, _06382_, _04292_);
  nor (_08370_, _08369_, _08368_);
  and (_08371_, _08370_, _08367_);
  and (_08372_, _06355_, _04256_);
  and (_08373_, _06340_, _04253_);
  nor (_08374_, _08373_, _08372_);
  and (_08375_, _06384_, _04295_);
  and (_08376_, _06361_, _04278_);
  nor (_08377_, _08376_, _08375_);
  and (_08378_, _08377_, _08374_);
  and (_08379_, _08378_, _08371_);
  and (_08380_, _06373_, _04242_);
  and (_08381_, _06379_, _04281_);
  nor (_08382_, _08381_, _08380_);
  and (_08383_, _06336_, _00567_);
  and (_08384_, _06371_, _04260_);
  nor (_08385_, _08384_, _08383_);
  and (_08386_, _08385_, _08382_);
  and (_08387_, _06359_, _04264_);
  and (_08388_, _06348_, _04287_);
  nor (_08389_, _08388_, _08387_);
  and (_08390_, _06345_, _04210_);
  and (_08391_, _06352_, _04237_);
  nor (_08392_, _08391_, _08390_);
  and (_08393_, _08392_, _08389_);
  and (_08394_, _08393_, _08386_);
  and (_08395_, _08394_, _08379_);
  nor (_08396_, _08395_, _07925_);
  and (_08397_, _08396_, _07133_);
  not (_08398_, _07086_);
  not (_08399_, _07855_);
  not (_08400_, _06071_);
  nor (_08401_, _06877_, _08400_);
  and (_08402_, _08401_, _06479_);
  and (_08403_, _08402_, _06206_);
  and (_08404_, _08403_, _07792_);
  nand (_08405_, _08404_, \oc8051_golden_model_1.PSW [7]);
  and (_08406_, _08402_, _06207_);
  and (_08407_, _08406_, _07787_);
  nand (_08408_, _08407_, \oc8051_golden_model_1.TCON [7]);
  and (_08409_, _08403_, _07807_);
  nand (_08410_, _08409_, \oc8051_golden_model_1.ACC [7]);
  and (_08411_, _08410_, _08408_);
  nand (_08412_, _08411_, _08405_);
  and (_08413_, _08406_, _07777_);
  nand (_08414_, _08413_, \oc8051_golden_model_1.SCON [7]);
  and (_08415_, _08406_, _07829_);
  nand (_08416_, _08415_, \oc8051_golden_model_1.IP [7]);
  nand (_08417_, _08416_, _08414_);
  and (_08418_, _08406_, _07825_);
  nand (_08419_, _08418_, \oc8051_golden_model_1.IE [7]);
  and (_08420_, _08403_, _07839_);
  nand (_08421_, _08420_, \oc8051_golden_model_1.B [7]);
  nand (_08422_, _08421_, _08419_);
  or (_08423_, _08422_, _08417_);
  or (_08424_, _08423_, _08412_);
  or (_08425_, _08424_, _07924_);
  and (_08426_, _08425_, _08399_);
  or (_08427_, _08426_, _08398_);
  not (_08428_, _06159_);
  not (_08429_, _06162_);
  not (_08430_, \oc8051_golden_model_1.ACC [7]);
  nor (_08431_, _06581_, _08430_);
  and (_08432_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_08433_, _08432_, \oc8051_golden_model_1.PC [6]);
  and (_08434_, _08433_, _05972_);
  and (_08435_, _08434_, \oc8051_golden_model_1.PC [7]);
  nor (_08436_, _08434_, \oc8051_golden_model_1.PC [7]);
  nor (_08437_, _08436_, _08435_);
  and (_08438_, _08437_, _06581_);
  or (_08439_, _08438_, _08431_);
  not (_08440_, _06129_);
  nor (_08441_, _08440_, _06125_);
  nor (_08442_, _08441_, _05762_);
  nor (_08443_, _08442_, _07259_);
  and (_08444_, _08443_, _08439_);
  not (_08445_, _08443_);
  and (_08446_, _08445_, _08358_);
  or (_08447_, _08446_, _08444_);
  and (_08448_, _08447_, _07065_);
  nor (_08449_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_08450_, _08449_, _06566_);
  nor (_08451_, _08450_, _06216_);
  nor (_08452_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_08453_, _08452_, _06216_);
  and (_08454_, _08453_, _06142_);
  nor (_08455_, _08454_, _08451_);
  nor (_08456_, _08455_, _06980_);
  not (_08457_, _08456_);
  or (_08458_, _07544_, _06701_);
  not (_08459_, _06980_);
  and (_08460_, _06701_, _06070_);
  nor (_08461_, _08460_, _08459_);
  nand (_08462_, _08461_, _08458_);
  and (_08463_, _08462_, _08457_);
  nor (_08464_, _08449_, _06566_);
  nor (_08465_, _08464_, _08450_);
  nor (_08466_, _08465_, _06980_);
  not (_08467_, _08466_);
  or (_08468_, _07708_, _06701_);
  and (_08469_, _06701_, _06625_);
  nor (_08470_, _08469_, _08459_);
  nand (_08471_, _08470_, _08468_);
  and (_08472_, _08471_, _08467_);
  or (_08473_, _07049_, _06701_);
  and (_08474_, _06701_, _06107_);
  nor (_08475_, _08474_, _08459_);
  nand (_08476_, _08475_, _08473_);
  nor (_08477_, _06980_, \oc8051_golden_model_1.SP [0]);
  not (_08478_, _08477_);
  nand (_08479_, _08478_, _08476_);
  or (_08480_, _08479_, _07863_);
  nor (_08481_, _07179_, _06980_);
  not (_08482_, _08481_);
  and (_08483_, _07306_, _07104_);
  nor (_08484_, _06912_, _07104_);
  or (_08485_, _08484_, _08459_);
  or (_08486_, _08485_, _08483_);
  nand (_08487_, _08486_, _08482_);
  and (_08488_, _08478_, _08476_);
  or (_08489_, _08488_, _07865_);
  and (_08490_, _08489_, _08487_);
  nand (_08491_, _08490_, _08480_);
  or (_08492_, _08479_, _07871_);
  and (_08493_, _08486_, _08482_);
  or (_08494_, _08488_, _07869_);
  and (_08495_, _08494_, _08493_);
  nand (_08496_, _08495_, _08492_);
  nand (_08497_, _08496_, _08491_);
  nand (_08498_, _08497_, _08472_);
  not (_08499_, _08472_);
  or (_08500_, _08479_, _07883_);
  or (_08501_, _08488_, _07885_);
  and (_08502_, _08501_, _08487_);
  nand (_08503_, _08502_, _08500_);
  or (_08504_, _08479_, _07879_);
  or (_08505_, _08488_, _07877_);
  and (_08506_, _08505_, _08493_);
  nand (_08507_, _08506_, _08504_);
  nand (_08508_, _08507_, _08503_);
  nand (_08509_, _08508_, _08499_);
  nand (_08510_, _08509_, _08498_);
  nand (_08511_, _08510_, _08463_);
  not (_08512_, _08463_);
  or (_08513_, _08479_, _07895_);
  or (_08514_, _08488_, _07893_);
  and (_08515_, _08514_, _08493_);
  nand (_08516_, _08515_, _08513_);
  or (_08517_, _08479_, _07899_);
  or (_08518_, _08488_, _07901_);
  and (_08519_, _08518_, _08487_);
  nand (_08520_, _08519_, _08517_);
  nand (_08521_, _08520_, _08516_);
  nand (_08522_, _08521_, _08472_);
  or (_08523_, _08479_, _07913_);
  or (_08524_, _08488_, _07915_);
  and (_08525_, _08524_, _08487_);
  nand (_08526_, _08525_, _08523_);
  or (_08527_, _08479_, _07909_);
  or (_08528_, _08488_, _07907_);
  and (_08529_, _08528_, _08493_);
  nand (_08530_, _08529_, _08527_);
  nand (_08531_, _08530_, _08526_);
  nand (_08532_, _08531_, _08499_);
  nand (_08533_, _08532_, _08522_);
  nand (_08534_, _08533_, _08512_);
  and (_08535_, _08534_, _08511_);
  and (_08536_, _08535_, _07064_);
  or (_08537_, _08536_, _08448_);
  and (_08538_, _08537_, _08429_);
  and (_08539_, _08338_, _08103_);
  not (_08540_, _08211_);
  and (_08541_, _08540_, _08175_);
  and (_08542_, _08247_, _08139_);
  and (_08543_, _08542_, _08541_);
  and (_08544_, _08543_, _08539_);
  and (_08545_, _08544_, _08014_);
  or (_08546_, _08545_, _07926_);
  nand (_08547_, _08545_, _07926_);
  and (_08548_, _08547_, _08546_);
  and (_08549_, _08548_, _06162_);
  or (_08550_, _08549_, _08538_);
  and (_08551_, _08550_, _08428_);
  or (_08552_, _08425_, _07855_);
  and (_08553_, _08552_, _06159_);
  or (_08554_, _08553_, _07485_);
  or (_08555_, _08554_, _08551_);
  nor (_08556_, _08437_, _05764_);
  nor (_08557_, _08556_, _07076_);
  and (_08558_, _08557_, _08555_);
  and (_08559_, _07923_, _07076_);
  or (_08560_, _08559_, _07086_);
  or (_08561_, _08560_, _08558_);
  and (_08562_, _08561_, _08427_);
  or (_08563_, _08562_, _06151_);
  nand (_08564_, _07925_, _06151_);
  and (_08565_, _08564_, _06149_);
  and (_08566_, _08565_, _08563_);
  and (_08567_, _08425_, _07855_);
  not (_08568_, _08567_);
  and (_08569_, _08568_, _08552_);
  and (_08570_, _08569_, _06148_);
  or (_08571_, _08570_, _08566_);
  and (_08572_, _08571_, _05760_);
  not (_08573_, _08437_);
  or (_08574_, _08573_, _05760_);
  nand (_08575_, _08574_, _06251_);
  or (_08576_, _08575_, _08572_);
  nand (_08577_, _07925_, _06252_);
  and (_08578_, _08577_, _08576_);
  or (_08579_, _08578_, _06701_);
  not (_08580_, _07103_);
  and (_08581_, _08535_, _06172_);
  or (_08582_, _07862_, _07104_);
  or (_08583_, _08582_, _08581_);
  and (_08584_, _08583_, _08580_);
  and (_08585_, _08584_, _08579_);
  and (_08586_, _07855_, \oc8051_golden_model_1.PSW [7]);
  or (_08587_, _08586_, _08426_);
  and (_08588_, _08587_, _07103_);
  or (_08589_, _08588_, _05791_);
  or (_08590_, _08589_, _08585_);
  nor (_08591_, _06132_, _06039_);
  and (_08592_, _08573_, _05791_);
  nor (_08593_, _08592_, _08591_);
  and (_08594_, _08593_, _08590_);
  nor (_08595_, _06117_, _06039_);
  and (_08596_, _07923_, _08591_);
  or (_08597_, _08596_, _08595_);
  or (_08598_, _08597_, _08594_);
  nor (_08599_, _06039_, _06114_);
  not (_08600_, _08599_);
  not (_08601_, _08595_);
  or (_08602_, _08535_, _08601_);
  and (_08603_, _08602_, _08600_);
  and (_08604_, _08603_, _08598_);
  and (_08605_, _08395_, _07923_);
  and (_08606_, _06945_, _06758_);
  not (_08607_, _08395_);
  and (_08608_, _06359_, _04687_);
  and (_08609_, _06368_, _04679_);
  nor (_08610_, _08609_, _08608_);
  and (_08611_, _06371_, _04671_);
  and (_08612_, _06382_, _04668_);
  nor (_08613_, _08612_, _08611_);
  and (_08614_, _08613_, _08610_);
  and (_08615_, _06384_, _04693_);
  and (_08616_, _06366_, _04673_);
  nor (_08617_, _08616_, _08615_);
  and (_08618_, _06355_, _04695_);
  and (_08619_, _06340_, _04699_);
  nor (_08620_, _08619_, _08618_);
  and (_08621_, _08620_, _08617_);
  and (_08622_, _08621_, _08614_);
  and (_08623_, _06345_, _04666_);
  and (_08624_, _06373_, _04697_);
  nor (_08625_, _08624_, _08623_);
  and (_08626_, _06336_, _00612_);
  and (_08627_, _06352_, _04682_);
  nor (_08628_, _08627_, _08626_);
  and (_08629_, _08628_, _08625_);
  and (_08630_, _06361_, _04677_);
  and (_08631_, _06348_, _04689_);
  nor (_08632_, _08631_, _08630_);
  and (_08633_, _06377_, _04705_);
  and (_08634_, _06379_, _04684_);
  nor (_08635_, _08634_, _08633_);
  and (_08636_, _08635_, _08632_);
  and (_08637_, _08636_, _08629_);
  and (_08638_, _08637_, _08622_);
  and (_08639_, _08638_, _08607_);
  and (_08640_, _06359_, _04614_);
  and (_08641_, _06368_, _04588_);
  nor (_08642_, _08641_, _08640_);
  and (_08643_, _06377_, _04596_);
  and (_08644_, _06352_, _04591_);
  nor (_08645_, _08644_, _08643_);
  and (_08646_, _08645_, _08642_);
  and (_08647_, _06355_, _04608_);
  and (_08648_, _06340_, _04606_);
  nor (_08649_, _08648_, _08647_);
  and (_08650_, _06384_, _04602_);
  and (_08651_, _06361_, _04586_);
  nor (_08652_, _08651_, _08650_);
  and (_08653_, _08652_, _08649_);
  and (_08654_, _08653_, _08646_);
  and (_08655_, _06382_, _04575_);
  and (_08656_, _06345_, _04580_);
  nor (_08657_, _08656_, _08655_);
  and (_08658_, _06336_, _00602_);
  and (_08659_, _06371_, _04582_);
  nor (_08660_, _08659_, _08658_);
  and (_08661_, _08660_, _08657_);
  and (_08662_, _06366_, _04577_);
  and (_08663_, _06348_, _04598_);
  nor (_08664_, _08663_, _08662_);
  and (_08665_, _06373_, _04604_);
  and (_08666_, _06379_, _04593_);
  nor (_08667_, _08666_, _08665_);
  and (_08668_, _08667_, _08664_);
  and (_08669_, _08668_, _08661_);
  and (_08670_, _08669_, _08654_);
  and (_08671_, _06359_, _04641_);
  and (_08672_, _06340_, _04654_);
  nor (_08673_, _08672_, _08671_);
  and (_08674_, _06379_, _04638_);
  and (_08675_, _06355_, _04650_);
  nor (_08676_, _08675_, _08674_);
  and (_08677_, _08676_, _08673_);
  and (_08678_, _06345_, _04620_);
  and (_08679_, _06348_, _04643_);
  nor (_08680_, _08679_, _08678_);
  and (_08681_, _06371_, _04625_);
  and (_08682_, _06382_, _04622_);
  nor (_08683_, _08682_, _08681_);
  and (_08684_, _08683_, _08680_);
  and (_08685_, _08684_, _08677_);
  and (_08686_, _06377_, _04660_);
  and (_08687_, _06368_, _04633_);
  nor (_08688_, _08687_, _08686_);
  and (_08689_, _06352_, _04636_);
  and (_08690_, _06384_, _04648_);
  nor (_08691_, _08690_, _08689_);
  and (_08692_, _08691_, _08688_);
  and (_08693_, _06373_, _04652_);
  and (_08694_, _06361_, _04631_);
  nor (_08695_, _08694_, _08693_);
  and (_08696_, _06336_, _00607_);
  and (_08697_, _06366_, _04627_);
  nor (_08698_, _08697_, _08696_);
  and (_08699_, _08698_, _08695_);
  and (_08700_, _08699_, _08692_);
  and (_08701_, _08700_, _08685_);
  and (_08702_, _08701_, _08670_);
  and (_08703_, _08702_, _08639_);
  nor (_08704_, _06521_, _06389_);
  and (_08705_, _08704_, _08703_);
  and (_08706_, _08705_, _08606_);
  and (_08707_, _08706_, \oc8051_golden_model_1.TH0 [7]);
  not (_08708_, _06758_);
  and (_08709_, _06945_, _08708_);
  and (_08710_, _08709_, _08705_);
  and (_08711_, _08710_, \oc8051_golden_model_1.TH1 [7]);
  not (_08712_, _06389_);
  and (_08713_, _06521_, _08712_);
  and (_08714_, _08713_, _08606_);
  not (_08715_, _08670_);
  and (_08716_, _08701_, _08715_);
  and (_08717_, _08716_, _08639_);
  and (_08718_, _08717_, _08714_);
  and (_08719_, _08718_, \oc8051_golden_model_1.SCON [7]);
  or (_08720_, _08719_, _08711_);
  or (_08721_, _08720_, _08707_);
  nor (_08722_, _06945_, _06758_);
  and (_08723_, _08722_, _08703_);
  and (_08724_, _08723_, _08713_);
  and (_08725_, _08724_, \oc8051_golden_model_1.TL1 [7]);
  and (_08726_, _08714_, _08703_);
  and (_08727_, _08726_, \oc8051_golden_model_1.TCON [7]);
  or (_08728_, _08727_, _08725_);
  or (_08729_, _08728_, _08721_);
  and (_08730_, _06521_, _06389_);
  and (_08731_, _08730_, _08606_);
  nor (_08732_, _08638_, _08395_);
  and (_08733_, _08732_, _08731_);
  and (_08734_, _08716_, _08733_);
  and (_08735_, _08734_, \oc8051_golden_model_1.PSW [7]);
  not (_08736_, _08701_);
  and (_08737_, _08736_, _08670_);
  and (_08738_, _08733_, _08737_);
  and (_08739_, _08738_, \oc8051_golden_model_1.ACC [7]);
  nor (_08740_, _08701_, _08670_);
  and (_08741_, _08733_, _08740_);
  and (_08742_, _08741_, \oc8051_golden_model_1.B [7]);
  or (_08743_, _08742_, _08739_);
  or (_08744_, _08743_, _08735_);
  and (_08745_, _08740_, _08639_);
  and (_08746_, _08745_, _08714_);
  and (_08747_, _08746_, \oc8051_golden_model_1.IP [7]);
  and (_08748_, _08737_, _08639_);
  and (_08749_, _08748_, _08714_);
  and (_08750_, _08749_, \oc8051_golden_model_1.IE [7]);
  and (_08751_, _08713_, _08709_);
  and (_08752_, _08751_, _08717_);
  and (_08753_, _08752_, \oc8051_golden_model_1.SBUF [7]);
  or (_08754_, _08753_, _08750_);
  or (_08755_, _08754_, _08747_);
  or (_08756_, _08755_, _08744_);
  and (_08757_, _08730_, _08703_);
  and (_08758_, _08757_, _08709_);
  and (_08759_, _08758_, \oc8051_golden_model_1.SP [7]);
  and (_08760_, _08730_, _08723_);
  and (_08761_, _08760_, \oc8051_golden_model_1.DPH [7]);
  or (_08762_, _08761_, _08759_);
  not (_08763_, _06945_);
  and (_08764_, _08763_, _06758_);
  and (_08765_, _08757_, _08764_);
  and (_08766_, _08765_, \oc8051_golden_model_1.DPL [7]);
  or (_08767_, _08766_, _08762_);
  not (_08768_, _06521_);
  and (_08769_, _08768_, _06389_);
  and (_08770_, _08769_, _08723_);
  and (_08771_, _08770_, \oc8051_golden_model_1.PCON [7]);
  and (_08772_, _08713_, _08703_);
  and (_08773_, _08772_, _08764_);
  and (_08774_, _08773_, \oc8051_golden_model_1.TL0 [7]);
  and (_08775_, _08751_, _08703_);
  and (_08776_, _08775_, \oc8051_golden_model_1.TMOD [7]);
  or (_08777_, _08776_, _08774_);
  or (_08778_, _08777_, _08771_);
  or (_08779_, _08778_, _08767_);
  or (_08780_, _08779_, _08756_);
  or (_08781_, _08780_, _08729_);
  or (_08782_, _08781_, _08605_);
  and (_08783_, _08782_, _08599_);
  not (_08784_, _07184_);
  nor (_08785_, _07115_, _07370_);
  and (_08786_, _08785_, _08784_);
  and (_08787_, _08786_, _07352_);
  not (_08788_, _08787_);
  or (_08789_, _08788_, _08783_);
  or (_08790_, _08789_, _08604_);
  nor (_08791_, _08787_, _06039_);
  nor (_08792_, _08791_, _06112_);
  and (_08793_, _08792_, _08790_);
  and (_08794_, _08607_, _06112_);
  or (_08795_, _08794_, _06076_);
  or (_08796_, _08795_, _08793_);
  nor (_08797_, _08437_, _05836_);
  nor (_08798_, _08797_, _07128_);
  and (_08799_, _08798_, _08796_);
  not (_08800_, _08396_);
  nand (_08801_, _08395_, _07925_);
  and (_08802_, _08801_, _08800_);
  nor (_08803_, _08802_, _07126_);
  nor (_08804_, _08803_, _07129_);
  or (_08805_, _08804_, _08799_);
  not (_08806_, _07133_);
  not (_08807_, _07126_);
  nor (_08808_, _07925_, _08430_);
  and (_08809_, _07925_, _08430_);
  nor (_08810_, _08809_, _08808_);
  or (_08811_, _08810_, _08807_);
  and (_08812_, _08811_, _08806_);
  and (_08813_, _08812_, _08805_);
  or (_08814_, _08813_, _08397_);
  and (_08815_, _08814_, _08364_);
  and (_08816_, _08808_, _07131_);
  or (_08817_, _08816_, _07124_);
  or (_08818_, _08817_, _08815_);
  not (_08819_, _06303_);
  nor (_08820_, _08819_, _06039_);
  nor (_08821_, _08437_, _05848_);
  nor (_08822_, _08821_, _08820_);
  and (_08823_, _08822_, _08818_);
  not (_08824_, _06396_);
  nor (_08825_, _08824_, _06039_);
  and (_08826_, _08801_, _08820_);
  or (_08827_, _08826_, _08825_);
  or (_08828_, _08827_, _08823_);
  nand (_08829_, _08809_, _08825_);
  and (_08830_, _08829_, _05846_);
  and (_08831_, _08830_, _08828_);
  or (_08832_, _08573_, _05846_);
  nand (_08833_, _08832_, _08362_);
  or (_08834_, _08833_, _08831_);
  and (_08835_, _08834_, _08363_);
  or (_08836_, _08835_, _07153_);
  not (_08837_, _07152_);
  nand (_08838_, _08534_, _08511_);
  or (_08839_, _08479_, _07960_);
  or (_08840_, _08488_, _07962_);
  and (_08841_, _08840_, _08487_);
  nand (_08842_, _08841_, _08839_);
  or (_08843_, _08479_, _07968_);
  or (_08844_, _08488_, _07966_);
  and (_08845_, _08844_, _08493_);
  nand (_08846_, _08845_, _08843_);
  nand (_08847_, _08846_, _08842_);
  nand (_08848_, _08847_, _08472_);
  or (_08849_, _08479_, _07980_);
  or (_08850_, _08488_, _07982_);
  and (_08851_, _08850_, _08487_);
  nand (_08852_, _08851_, _08849_);
  or (_08853_, _08479_, _07976_);
  or (_08854_, _08488_, _07974_);
  and (_08855_, _08854_, _08493_);
  nand (_08856_, _08855_, _08853_);
  nand (_08857_, _08856_, _08852_);
  nand (_08858_, _08857_, _08499_);
  and (_08859_, _08858_, _08463_);
  and (_08860_, _08859_, _08848_);
  or (_08861_, _08479_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_08862_, _08488_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_08863_, _08862_, _08861_);
  nand (_08864_, _08863_, _08493_);
  or (_08865_, _08479_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_08866_, _08488_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_08867_, _08866_, _08865_);
  nand (_08868_, _08867_, _08487_);
  nand (_08869_, _08868_, _08864_);
  nand (_08870_, _08869_, _08472_);
  or (_08871_, _08479_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_08872_, _08488_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_08873_, _08872_, _08871_);
  nand (_08874_, _08873_, _08493_);
  or (_08875_, _08479_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_08876_, _08488_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand (_08877_, _08876_, _08875_);
  nand (_08878_, _08877_, _08487_);
  nand (_08879_, _08878_, _08874_);
  nand (_08880_, _08879_, _08499_);
  and (_08881_, _08880_, _08512_);
  and (_08882_, _08881_, _08870_);
  nor (_08883_, _08882_, _08860_);
  or (_08884_, _08479_, _08049_);
  or (_08885_, _08488_, _08051_);
  and (_08886_, _08885_, _08487_);
  nand (_08887_, _08886_, _08884_);
  or (_08888_, _08479_, _08057_);
  or (_08889_, _08488_, _08055_);
  and (_08890_, _08889_, _08493_);
  nand (_08891_, _08890_, _08888_);
  nand (_08892_, _08891_, _08887_);
  nand (_08893_, _08892_, _08472_);
  or (_08894_, _08479_, _08069_);
  or (_08895_, _08488_, _08071_);
  and (_08896_, _08895_, _08487_);
  nand (_08897_, _08896_, _08894_);
  or (_08898_, _08479_, _08065_);
  or (_08899_, _08488_, _08063_);
  and (_08900_, _08899_, _08493_);
  nand (_08901_, _08900_, _08898_);
  nand (_08902_, _08901_, _08897_);
  nand (_08903_, _08902_, _08499_);
  and (_08904_, _08903_, _08463_);
  and (_08906_, _08904_, _08893_);
  or (_08907_, _08479_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_08908_, _08488_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_08909_, _08908_, _08907_);
  nand (_08910_, _08909_, _08493_);
  or (_08911_, _08479_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_08912_, _08488_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_08913_, _08912_, _08911_);
  nand (_08914_, _08913_, _08487_);
  nand (_08915_, _08914_, _08910_);
  nand (_08917_, _08915_, _08472_);
  or (_08918_, _08479_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_08919_, _08488_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_08920_, _08919_, _08918_);
  nand (_08921_, _08920_, _08493_);
  or (_08922_, _08479_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_08923_, _08488_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand (_08924_, _08923_, _08922_);
  nand (_08925_, _08924_, _08487_);
  nand (_08926_, _08925_, _08921_);
  nand (_08928_, _08926_, _08499_);
  and (_08929_, _08928_, _08512_);
  and (_08930_, _08929_, _08917_);
  nor (_08931_, _08930_, _08906_);
  or (_08932_, _08479_, _08284_);
  or (_08933_, _08488_, _08286_);
  and (_08934_, _08933_, _08487_);
  nand (_08935_, _08934_, _08932_);
  or (_08936_, _08479_, _08292_);
  or (_08937_, _08488_, _08290_);
  and (_08939_, _08937_, _08493_);
  nand (_08940_, _08939_, _08936_);
  nand (_08941_, _08940_, _08935_);
  nand (_08942_, _08941_, _08472_);
  or (_08943_, _08479_, _08304_);
  or (_08944_, _08488_, _08306_);
  and (_08945_, _08944_, _08487_);
  nand (_08946_, _08945_, _08943_);
  or (_08947_, _08479_, _08300_);
  or (_08948_, _08488_, _08298_);
  and (_08950_, _08948_, _08493_);
  nand (_08951_, _08950_, _08947_);
  nand (_08952_, _08951_, _08946_);
  nand (_08953_, _08952_, _08499_);
  and (_08954_, _08953_, _08463_);
  and (_08955_, _08954_, _08942_);
  or (_08956_, _08479_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_08957_, _08488_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_08958_, _08957_, _08956_);
  nand (_08959_, _08958_, _08493_);
  or (_08961_, _08479_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_08962_, _08488_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_08963_, _08962_, _08961_);
  nand (_08964_, _08963_, _08487_);
  nand (_08965_, _08964_, _08959_);
  nand (_08966_, _08965_, _08472_);
  or (_08967_, _08479_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_08968_, _08488_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_08969_, _08968_, _08967_);
  nand (_08970_, _08969_, _08493_);
  or (_08972_, _08479_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_08973_, _08488_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand (_08974_, _08973_, _08972_);
  nand (_08975_, _08974_, _08487_);
  nand (_08976_, _08975_, _08970_);
  nand (_08977_, _08976_, _08499_);
  and (_08978_, _08977_, _08512_);
  and (_08979_, _08978_, _08966_);
  nor (_08980_, _08979_, _08955_);
  or (_08981_, _08479_, _07422_);
  or (_08982_, _08488_, _07424_);
  and (_08983_, _08982_, _08487_);
  nand (_08984_, _08983_, _08981_);
  or (_08985_, _08479_, _07430_);
  or (_08986_, _08488_, _07428_);
  and (_08987_, _08986_, _08493_);
  nand (_08988_, _08987_, _08985_);
  nand (_08989_, _08988_, _08984_);
  nand (_08990_, _08989_, _08472_);
  or (_08991_, _08479_, _07442_);
  or (_08992_, _08488_, _07444_);
  and (_08993_, _08992_, _08487_);
  nand (_08994_, _08993_, _08991_);
  or (_08995_, _08479_, _07438_);
  or (_08996_, _08488_, _07436_);
  and (_08997_, _08996_, _08493_);
  nand (_08998_, _08997_, _08995_);
  nand (_08999_, _08998_, _08994_);
  nand (_09000_, _08999_, _08499_);
  and (_09001_, _09000_, _08463_);
  and (_09002_, _09001_, _08990_);
  or (_09003_, _08479_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_09004_, _08488_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_09005_, _09004_, _09003_);
  nand (_09006_, _09005_, _08493_);
  or (_09007_, _08479_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_09008_, _08488_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_09009_, _09008_, _09007_);
  nand (_09010_, _09009_, _08487_);
  nand (_09011_, _09010_, _09006_);
  nand (_09012_, _09011_, _08472_);
  or (_09013_, _08479_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_09014_, _08488_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_09015_, _09014_, _09013_);
  nand (_09016_, _09015_, _08493_);
  or (_09017_, _08479_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_09018_, _08488_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_09019_, _09018_, _09017_);
  nand (_09020_, _09019_, _08487_);
  nand (_09021_, _09020_, _09016_);
  nand (_09022_, _09021_, _08499_);
  and (_09023_, _09022_, _08512_);
  and (_09024_, _09023_, _09012_);
  nor (_09025_, _09024_, _09002_);
  or (_09026_, _08479_, _07603_);
  or (_09027_, _08488_, _07605_);
  and (_09028_, _09027_, _08487_);
  nand (_09029_, _09028_, _09026_);
  or (_09030_, _08479_, _07611_);
  or (_09031_, _08488_, _07609_);
  and (_09032_, _09031_, _08493_);
  nand (_09033_, _09032_, _09030_);
  nand (_09034_, _09033_, _09029_);
  nand (_09035_, _09034_, _08472_);
  or (_09036_, _08479_, _07623_);
  or (_09037_, _08488_, _07625_);
  and (_09038_, _09037_, _08487_);
  nand (_09039_, _09038_, _09036_);
  or (_09040_, _08479_, _07619_);
  or (_09041_, _08488_, _07617_);
  and (_09042_, _09041_, _08493_);
  nand (_09043_, _09042_, _09040_);
  nand (_09044_, _09043_, _09039_);
  nand (_09045_, _09044_, _08499_);
  and (_09046_, _09045_, _08463_);
  and (_09047_, _09046_, _09035_);
  or (_09048_, _08479_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_09049_, _08488_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_09050_, _09049_, _09048_);
  nand (_09051_, _09050_, _08493_);
  or (_09052_, _08479_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_09053_, _08488_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_09054_, _09053_, _09052_);
  nand (_09055_, _09054_, _08487_);
  nand (_09056_, _09055_, _09051_);
  nand (_09057_, _09056_, _08472_);
  or (_09058_, _08479_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_09059_, _08488_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_09060_, _09059_, _09058_);
  nand (_09061_, _09060_, _08493_);
  or (_09062_, _08479_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_09063_, _08488_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_09064_, _09063_, _09062_);
  nand (_09065_, _09064_, _08487_);
  nand (_09066_, _09065_, _09061_);
  nand (_09067_, _09066_, _08499_);
  and (_09068_, _09067_, _08512_);
  and (_09069_, _09068_, _09057_);
  nor (_09070_, _09069_, _09047_);
  or (_09071_, _08479_, _07193_);
  or (_09072_, _08488_, _07195_);
  and (_09073_, _09072_, _08487_);
  nand (_09074_, _09073_, _09071_);
  or (_09075_, _08479_, _07201_);
  or (_09076_, _08488_, _07199_);
  and (_09077_, _09076_, _08493_);
  nand (_09078_, _09077_, _09075_);
  nand (_09079_, _09078_, _09074_);
  nand (_09080_, _09079_, _08472_);
  or (_09081_, _08479_, _07213_);
  or (_09082_, _08488_, _07215_);
  and (_09083_, _09082_, _08487_);
  nand (_09084_, _09083_, _09081_);
  or (_09085_, _08479_, _07209_);
  or (_09086_, _08488_, _07207_);
  and (_09087_, _09086_, _08493_);
  nand (_09088_, _09087_, _09085_);
  nand (_09089_, _09088_, _09084_);
  nand (_09090_, _09089_, _08499_);
  and (_09091_, _09090_, _08463_);
  and (_09092_, _09091_, _09080_);
  or (_09093_, _08479_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_09094_, _08488_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_09095_, _09094_, _09093_);
  nand (_09096_, _09095_, _08493_);
  or (_09097_, _08479_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_09098_, _08488_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_09099_, _09098_, _09097_);
  nand (_09100_, _09099_, _08487_);
  nand (_09101_, _09100_, _09096_);
  nand (_09102_, _09101_, _08472_);
  or (_09103_, _08479_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_09104_, _08488_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_09105_, _09104_, _09103_);
  nand (_09106_, _09105_, _08493_);
  or (_09107_, _08479_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_09108_, _08488_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_09109_, _09108_, _09107_);
  nand (_09110_, _09109_, _08487_);
  nand (_09111_, _09110_, _09106_);
  nand (_09112_, _09111_, _08499_);
  and (_09113_, _09112_, _08512_);
  and (_09114_, _09113_, _09102_);
  or (_09115_, _09114_, _09092_);
  or (_09116_, _08479_, _06638_);
  or (_09117_, _08488_, _06992_);
  and (_09118_, _09117_, _08487_);
  nand (_09119_, _09118_, _09116_);
  or (_09120_, _08479_, _07000_);
  or (_09121_, _08488_, _06997_);
  and (_09122_, _09121_, _08493_);
  nand (_09123_, _09122_, _09120_);
  nand (_09124_, _09123_, _09119_);
  nand (_09125_, _09124_, _08472_);
  or (_09126_, _08479_, _07013_);
  or (_09127_, _08488_, _07015_);
  and (_09128_, _09127_, _08487_);
  nand (_09129_, _09128_, _09126_);
  or (_09130_, _08479_, _07009_);
  or (_09131_, _08488_, _07007_);
  and (_09132_, _09131_, _08493_);
  nand (_09133_, _09132_, _09130_);
  nand (_09134_, _09133_, _09129_);
  nand (_09135_, _09134_, _08499_);
  and (_09136_, _09135_, _08463_);
  and (_09137_, _09136_, _09125_);
  or (_09138_, _08479_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_09139_, _08488_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_09140_, _09139_, _09138_);
  nand (_09141_, _09140_, _08493_);
  or (_09142_, _08479_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_09143_, _08488_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_09144_, _09143_, _09142_);
  nand (_09145_, _09144_, _08487_);
  nand (_09146_, _09145_, _09141_);
  nand (_09147_, _09146_, _08472_);
  or (_09148_, _08479_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_09149_, _08488_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_09150_, _09149_, _09148_);
  nand (_09151_, _09150_, _08493_);
  or (_09152_, _08479_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_09153_, _08488_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand (_09154_, _09153_, _09152_);
  nand (_09155_, _09154_, _08487_);
  nand (_09156_, _09155_, _09151_);
  nand (_09157_, _09156_, _08499_);
  and (_09158_, _09157_, _08512_);
  and (_09159_, _09158_, _09147_);
  or (_09160_, _09159_, _09137_);
  nor (_09161_, _09160_, _09115_);
  and (_09162_, _09161_, _09070_);
  and (_09163_, _09162_, _09025_);
  and (_09164_, _09163_, _08980_);
  and (_09165_, _09164_, _08931_);
  and (_09166_, _09165_, _08883_);
  nor (_09167_, _09166_, _08838_);
  and (_09168_, _09166_, _08838_);
  or (_09169_, _09168_, _09167_);
  or (_09170_, _09169_, _07154_);
  and (_09171_, _09170_, _08837_);
  and (_09172_, _09171_, _08836_);
  and (_09173_, _08548_, _07152_);
  or (_09174_, _09173_, _06310_);
  or (_09175_, _09174_, _09172_);
  and (_09176_, _05449_, _05424_);
  and (_09177_, _09176_, _08433_);
  and (_09178_, _09177_, \oc8051_golden_model_1.PC [7]);
  nor (_09179_, _09177_, \oc8051_golden_model_1.PC [7]);
  nor (_09180_, _09179_, _09178_);
  not (_09181_, _09180_);
  nand (_09182_, _09181_, _06310_);
  and (_09183_, _09182_, _09175_);
  or (_09184_, _09183_, _05823_);
  and (_09185_, _08573_, _05823_);
  nor (_09186_, _09185_, _06073_);
  and (_09187_, _09186_, _09184_);
  and (_09188_, _08426_, _06073_);
  and (_09189_, _05820_, _05666_);
  nor (_09190_, _09189_, _09188_);
  not (_09191_, _09190_);
  nor (_09192_, _09191_, _09187_);
  not (_09193_, _09189_);
  nand (_09194_, _07922_, _07892_);
  and (_09195_, _07306_, _07049_);
  and (_09196_, _09195_, _07708_);
  and (_09197_, _09196_, _07544_);
  and (_09198_, _09197_, _08336_);
  and (_09199_, _09198_, _08101_);
  and (_09200_, _09199_, _08012_);
  nor (_09201_, _09200_, _09194_);
  and (_09202_, _09200_, _09194_);
  or (_09203_, _09202_, _09201_);
  nor (_09204_, _09203_, _09193_);
  nor (_09205_, _09204_, _09192_);
  nor (_09206_, _09205_, _07168_);
  or (_09207_, _08882_, _08860_);
  or (_09208_, _08930_, _08906_);
  or (_09209_, _08979_, _08955_);
  or (_09210_, _09024_, _09002_);
  or (_09211_, _09069_, _09047_);
  and (_09212_, _09160_, _09115_);
  and (_09213_, _09212_, _09211_);
  and (_09214_, _09213_, _09210_);
  and (_09215_, _09214_, _09209_);
  and (_09216_, _09215_, _09208_);
  and (_09217_, _09216_, _09207_);
  nor (_09218_, _09217_, _08838_);
  and (_09219_, _09217_, _08838_);
  or (_09220_, _09219_, _09218_);
  nor (_09221_, _09220_, _07169_);
  nor (_09222_, _09221_, _07167_);
  not (_09223_, _09222_);
  nor (_09224_, _09223_, _09206_);
  nor (_09225_, _09224_, _08346_);
  nor (_09226_, _09225_, _07418_);
  or (_09227_, _09226_, _07770_);
  and (_09228_, _09227_, _07769_);
  not (_09229_, \oc8051_golden_model_1.PC [15]);
  and (_09230_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and (_09231_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_09232_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_09233_, _09232_, _09231_);
  and (_09234_, _09233_, _09178_);
  and (_09235_, _09234_, _09230_);
  and (_09236_, _09235_, \oc8051_golden_model_1.PC [14]);
  and (_09237_, _09236_, _09229_);
  nor (_09238_, _09236_, _09229_);
  or (_09239_, _09238_, _09237_);
  not (_09240_, _09239_);
  nand (_09241_, _09240_, _06310_);
  and (_09242_, _09231_, \oc8051_golden_model_1.PC [10]);
  and (_09243_, _09242_, _08435_);
  and (_09244_, _09243_, \oc8051_golden_model_1.PC [11]);
  and (_09245_, _09244_, \oc8051_golden_model_1.PC [12]);
  and (_09246_, _09245_, \oc8051_golden_model_1.PC [13]);
  and (_09247_, _09246_, \oc8051_golden_model_1.PC [14]);
  nor (_09248_, _09247_, \oc8051_golden_model_1.PC [15]);
  and (_09249_, _09231_, _08435_);
  and (_09250_, _09249_, \oc8051_golden_model_1.PC [10]);
  and (_09251_, _09250_, \oc8051_golden_model_1.PC [11]);
  and (_09252_, _09251_, \oc8051_golden_model_1.PC [12]);
  and (_09253_, _09252_, \oc8051_golden_model_1.PC [13]);
  and (_09254_, _09253_, \oc8051_golden_model_1.PC [14]);
  and (_09255_, _09254_, \oc8051_golden_model_1.PC [15]);
  nor (_09256_, _09255_, _09248_);
  or (_09257_, _09256_, _06310_);
  and (_09258_, _09257_, _09241_);
  and (_09259_, _09258_, _07764_);
  and (_09260_, _09259_, _07767_);
  or (_40979_, _09260_, _09228_);
  not (_09261_, \oc8051_golden_model_1.B [7]);
  nor (_09262_, _01317_, _09261_);
  nor (_09263_, _07841_, _09261_);
  and (_09264_, _07923_, _07841_);
  or (_09265_, _09264_, _09263_);
  or (_09266_, _09265_, _06132_);
  nor (_09267_, _08420_, _09261_);
  and (_09268_, _08426_, _08420_);
  or (_09269_, _09268_, _09267_);
  and (_09270_, _09269_, _06152_);
  and (_09271_, _08548_, _07841_);
  or (_09272_, _09271_, _09263_);
  or (_09273_, _09272_, _06161_);
  and (_09274_, _07841_, \oc8051_golden_model_1.ACC [7]);
  or (_09275_, _09274_, _09263_);
  and (_09276_, _09275_, _07056_);
  nor (_09277_, _07056_, _09261_);
  or (_09278_, _09277_, _06160_);
  or (_09279_, _09278_, _09276_);
  and (_09280_, _09279_, _06157_);
  and (_09281_, _09280_, _09273_);
  and (_09282_, _08552_, _08420_);
  or (_09283_, _09282_, _09267_);
  and (_09284_, _09283_, _06156_);
  or (_09285_, _09284_, _06217_);
  or (_09286_, _09285_, _09281_);
  or (_09287_, _09265_, _07075_);
  and (_09288_, _09287_, _09286_);
  or (_09289_, _09288_, _06220_);
  or (_09290_, _09275_, _06229_);
  and (_09291_, _09290_, _06153_);
  and (_09292_, _09291_, _09289_);
  or (_09293_, _09292_, _09270_);
  and (_09294_, _09293_, _06146_);
  and (_09295_, _06294_, _06245_);
  or (_09296_, _09267_, _08568_);
  and (_09297_, _09283_, _06145_);
  and (_09298_, _09297_, _09296_);
  or (_09299_, _09298_, _09295_);
  or (_09300_, _09299_, _09294_);
  not (_09301_, _09295_);
  and (_09302_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_09303_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_09304_, _09303_, _09302_);
  and (_09305_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [2]);
  and (_09306_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  and (_09307_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_09308_, _09307_, _09306_);
  nor (_09309_, _09308_, _09304_);
  and (_09310_, _09309_, _09305_);
  nor (_09311_, _09310_, _09304_);
  and (_09312_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_09313_, _09312_, _09306_);
  and (_09314_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_09315_, _09314_, _09302_);
  nor (_09316_, _09315_, _09313_);
  not (_09317_, _09316_);
  nor (_09318_, _09317_, _09311_);
  and (_09319_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_09320_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [3]);
  and (_09321_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [4]);
  and (_09322_, _09321_, _09320_);
  nor (_09323_, _09321_, _09320_);
  nor (_09324_, _09323_, _09322_);
  and (_09325_, _09324_, _09319_);
  nor (_09326_, _09324_, _09319_);
  nor (_09327_, _09326_, _09325_);
  and (_09328_, _09317_, _09311_);
  nor (_09329_, _09328_, _09318_);
  and (_09330_, _09329_, _09327_);
  nor (_09331_, _09330_, _09318_);
  not (_09332_, _09306_);
  and (_09333_, _09312_, _09332_);
  and (_09334_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [5]);
  and (_09335_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_09336_, _09335_, _09320_);
  and (_09337_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [4]);
  and (_09338_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_09339_, _09338_, _09337_);
  nor (_09340_, _09339_, _09336_);
  and (_09341_, _09340_, _09334_);
  nor (_09342_, _09340_, _09334_);
  nor (_09343_, _09342_, _09341_);
  and (_09344_, _09343_, _09333_);
  nor (_09345_, _09343_, _09333_);
  nor (_09346_, _09345_, _09344_);
  not (_09347_, _09346_);
  nor (_09348_, _09347_, _09331_);
  and (_09349_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_09350_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [7]);
  and (_09351_, _09350_, _09349_);
  nor (_09352_, _09325_, _09322_);
  and (_09353_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.B [7]);
  and (_09354_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_09355_, _09354_, _09353_);
  nor (_09356_, _09354_, _09353_);
  nor (_09357_, _09356_, _09355_);
  not (_09358_, _09357_);
  nor (_09359_, _09358_, _09352_);
  and (_09360_, _09358_, _09352_);
  nor (_09361_, _09360_, _09359_);
  and (_09362_, _09361_, _09351_);
  nor (_09363_, _09361_, _09351_);
  nor (_09364_, _09363_, _09362_);
  and (_09365_, _09347_, _09331_);
  nor (_09366_, _09365_, _09348_);
  and (_09367_, _09366_, _09364_);
  nor (_09368_, _09367_, _09348_);
  nor (_09369_, _09341_, _09336_);
  and (_09370_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.B [7]);
  and (_09371_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [6]);
  and (_09372_, _09371_, _09370_);
  nor (_09373_, _09371_, _09370_);
  nor (_09374_, _09373_, _09372_);
  not (_09375_, _09374_);
  nor (_09376_, _09375_, _09369_);
  and (_09377_, _09375_, _09369_);
  nor (_09378_, _09377_, _09376_);
  and (_09379_, _09378_, _09355_);
  nor (_09380_, _09378_, _09355_);
  nor (_09381_, _09380_, _09379_);
  nor (_09382_, _09344_, _09313_);
  and (_09383_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [5]);
  and (_09384_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_09385_, _09384_, _09335_);
  nor (_09386_, _09384_, _09335_);
  nor (_09387_, _09386_, _09385_);
  and (_09388_, _09387_, _09383_);
  nor (_09389_, _09387_, _09383_);
  nor (_09390_, _09389_, _09388_);
  not (_09391_, _09390_);
  nor (_09392_, _09391_, _09382_);
  and (_09393_, _09391_, _09382_);
  nor (_09394_, _09393_, _09392_);
  and (_09395_, _09394_, _09381_);
  nor (_09396_, _09394_, _09381_);
  nor (_09397_, _09396_, _09395_);
  not (_09398_, _09397_);
  nor (_09399_, _09398_, _09368_);
  nor (_09400_, _09362_, _09359_);
  not (_09401_, _09400_);
  and (_09402_, _09398_, _09368_);
  nor (_09403_, _09402_, _09399_);
  and (_09404_, _09403_, _09401_);
  nor (_09405_, _09404_, _09399_);
  nor (_09406_, _09379_, _09376_);
  not (_09407_, _09406_);
  nor (_09408_, _09395_, _09392_);
  not (_09409_, _09408_);
  and (_09410_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_09411_, _09410_, _09335_);
  and (_09412_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_09413_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_09414_, _09413_, _09412_);
  nor (_09415_, _09414_, _09411_);
  nor (_09416_, _09388_, _09385_);
  and (_09417_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [7]);
  and (_09418_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [6]);
  and (_09419_, _09418_, _09417_);
  nor (_09420_, _09418_, _09417_);
  nor (_09421_, _09420_, _09419_);
  not (_09422_, _09421_);
  nor (_09423_, _09422_, _09416_);
  and (_09424_, _09422_, _09416_);
  nor (_09425_, _09424_, _09423_);
  and (_09426_, _09425_, _09372_);
  nor (_09427_, _09425_, _09372_);
  nor (_09428_, _09427_, _09426_);
  and (_09429_, _09428_, _09415_);
  nor (_09430_, _09428_, _09415_);
  nor (_09431_, _09430_, _09429_);
  and (_09432_, _09431_, _09409_);
  nor (_09433_, _09431_, _09409_);
  nor (_09434_, _09433_, _09432_);
  and (_09435_, _09434_, _09407_);
  nor (_09436_, _09434_, _09407_);
  nor (_09437_, _09436_, _09435_);
  not (_09438_, _09437_);
  nor (_09439_, _09438_, _09405_);
  nor (_09440_, _09435_, _09432_);
  nor (_09441_, _09426_, _09423_);
  not (_09442_, _09441_);
  and (_09443_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [7]);
  and (_09444_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_09445_, _09444_, _09443_);
  nor (_09446_, _09444_, _09443_);
  nor (_09447_, _09446_, _09445_);
  and (_09448_, _09447_, _09411_);
  nor (_09449_, _09447_, _09411_);
  nor (_09450_, _09449_, _09448_);
  and (_09451_, _09450_, _09419_);
  nor (_09452_, _09450_, _09419_);
  nor (_09453_, _09452_, _09451_);
  and (_09454_, _09453_, _09410_);
  nor (_09455_, _09453_, _09410_);
  nor (_09456_, _09455_, _09454_);
  and (_09457_, _09456_, _09429_);
  nor (_09458_, _09456_, _09429_);
  nor (_09459_, _09458_, _09457_);
  and (_09460_, _09459_, _09442_);
  nor (_09461_, _09459_, _09442_);
  nor (_09462_, _09461_, _09460_);
  not (_09463_, _09462_);
  nor (_09464_, _09463_, _09440_);
  and (_09465_, _09463_, _09440_);
  nor (_09466_, _09465_, _09464_);
  and (_09467_, _09466_, _09439_);
  nor (_09468_, _09460_, _09457_);
  nor (_09469_, _09451_, _09448_);
  not (_09470_, _09469_);
  and (_09471_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.B [7]);
  and (_09472_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_09473_, _09472_, _09471_);
  nor (_09474_, _09472_, _09471_);
  nor (_09475_, _09474_, _09473_);
  and (_09476_, _09475_, _09445_);
  nor (_09477_, _09475_, _09445_);
  nor (_09478_, _09477_, _09476_);
  and (_09479_, _09478_, _09454_);
  nor (_09480_, _09478_, _09454_);
  nor (_09481_, _09480_, _09479_);
  and (_09482_, _09481_, _09470_);
  nor (_09483_, _09481_, _09470_);
  nor (_09484_, _09483_, _09482_);
  not (_09485_, _09484_);
  nor (_09486_, _09485_, _09468_);
  and (_09487_, _09485_, _09468_);
  nor (_09488_, _09487_, _09486_);
  and (_09489_, _09488_, _09464_);
  nor (_09490_, _09488_, _09464_);
  nor (_09491_, _09490_, _09489_);
  and (_09492_, _09491_, _09467_);
  nor (_09493_, _09491_, _09467_);
  and (_09494_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  and (_09495_, _09494_, _09306_);
  and (_09496_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [2]);
  and (_09497_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [1]);
  nor (_09498_, _09497_, _09303_);
  nor (_09499_, _09498_, _09495_);
  and (_09500_, _09499_, _09496_);
  nor (_09501_, _09500_, _09495_);
  not (_09502_, _09501_);
  nor (_09503_, _09309_, _09305_);
  nor (_09504_, _09503_, _09310_);
  and (_09505_, _09504_, _09502_);
  and (_09506_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_09507_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [3]);
  and (_09508_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_09509_, _09508_, _09507_);
  nor (_09510_, _09508_, _09507_);
  nor (_09511_, _09510_, _09509_);
  and (_09512_, _09511_, _09506_);
  nor (_09513_, _09511_, _09506_);
  nor (_09514_, _09513_, _09512_);
  nor (_09515_, _09504_, _09502_);
  nor (_09516_, _09515_, _09505_);
  and (_09517_, _09516_, _09514_);
  nor (_09518_, _09517_, _09505_);
  nor (_09519_, _09329_, _09327_);
  nor (_09520_, _09519_, _09330_);
  not (_09522_, _09520_);
  nor (_09523_, _09522_, _09518_);
  and (_09524_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_09525_, _09524_, _09350_);
  nor (_09526_, _09512_, _09509_);
  nor (_09527_, _09350_, _09349_);
  nor (_09528_, _09527_, _09351_);
  not (_09529_, _09528_);
  nor (_09530_, _09529_, _09526_);
  and (_09531_, _09529_, _09526_);
  nor (_09532_, _09531_, _09530_);
  and (_09533_, _09532_, _09525_);
  nor (_09534_, _09532_, _09525_);
  nor (_09535_, _09534_, _09533_);
  and (_09536_, _09522_, _09518_);
  nor (_09537_, _09536_, _09523_);
  and (_09538_, _09537_, _09535_);
  nor (_09539_, _09538_, _09523_);
  nor (_09540_, _09366_, _09364_);
  nor (_09541_, _09540_, _09367_);
  not (_09543_, _09541_);
  nor (_09544_, _09543_, _09539_);
  nor (_09545_, _09533_, _09530_);
  not (_09546_, _09545_);
  and (_09547_, _09543_, _09539_);
  nor (_09548_, _09547_, _09544_);
  and (_09549_, _09548_, _09546_);
  nor (_09550_, _09549_, _09544_);
  nor (_09551_, _09403_, _09401_);
  nor (_09552_, _09551_, _09404_);
  not (_09553_, _09552_);
  nor (_09554_, _09553_, _09550_);
  and (_09555_, _09438_, _09405_);
  nor (_09556_, _09555_, _09439_);
  and (_09557_, _09556_, _09554_);
  nor (_09558_, _09466_, _09439_);
  nor (_09559_, _09558_, _09467_);
  nand (_09560_, _09559_, _09557_);
  and (_09561_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [1]);
  and (_09562_, _09561_, _09494_);
  and (_09563_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_09564_, _09561_, _09494_);
  nor (_09565_, _09564_, _09562_);
  and (_09566_, _09565_, _09563_);
  nor (_09567_, _09566_, _09562_);
  not (_09568_, _09567_);
  nor (_09569_, _09499_, _09496_);
  nor (_09570_, _09569_, _09500_);
  and (_09571_, _09570_, _09568_);
  and (_09572_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [5]);
  and (_09573_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_09574_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_09575_, _09574_, _09573_);
  nor (_09576_, _09574_, _09573_);
  nor (_09577_, _09576_, _09575_);
  and (_09578_, _09577_, _09572_);
  nor (_09579_, _09577_, _09572_);
  nor (_09580_, _09579_, _09578_);
  nor (_09581_, _09570_, _09568_);
  nor (_09582_, _09581_, _09571_);
  and (_09583_, _09582_, _09580_);
  nor (_09584_, _09583_, _09571_);
  not (_09585_, _09584_);
  nor (_09586_, _09516_, _09514_);
  nor (_09587_, _09586_, _09517_);
  and (_09588_, _09587_, _09585_);
  nor (_09589_, _09578_, _09575_);
  and (_09590_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [6]);
  and (_09591_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.B [7]);
  nor (_09592_, _09591_, _09590_);
  nor (_09593_, _09592_, _09525_);
  not (_09594_, _09593_);
  nor (_09595_, _09594_, _09589_);
  and (_09596_, _09594_, _09589_);
  nor (_09597_, _09596_, _09595_);
  nor (_09598_, _09587_, _09585_);
  nor (_09599_, _09598_, _09588_);
  and (_09600_, _09599_, _09597_);
  nor (_09601_, _09600_, _09588_);
  nor (_09602_, _09537_, _09535_);
  nor (_09603_, _09602_, _09538_);
  not (_09604_, _09603_);
  nor (_09605_, _09604_, _09601_);
  and (_09606_, _09604_, _09601_);
  nor (_09607_, _09606_, _09605_);
  and (_09608_, _09607_, _09595_);
  nor (_09609_, _09608_, _09605_);
  nor (_09610_, _09548_, _09546_);
  nor (_09611_, _09610_, _09549_);
  not (_09612_, _09611_);
  nor (_09613_, _09612_, _09609_);
  and (_09614_, _09553_, _09550_);
  nor (_09615_, _09614_, _09554_);
  and (_09616_, _09615_, _09613_);
  nor (_09617_, _09556_, _09554_);
  nor (_09618_, _09617_, _09557_);
  and (_09619_, _09618_, _09616_);
  nor (_09620_, _09618_, _09616_);
  nor (_09621_, _09620_, _09619_);
  and (_09622_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [0]);
  and (_09623_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_09624_, _09623_, _09622_);
  and (_09625_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_09626_, _09623_, _09622_);
  nor (_09627_, _09626_, _09624_);
  and (_09628_, _09627_, _09625_);
  nor (_09629_, _09628_, _09624_);
  not (_09630_, _09629_);
  nor (_09631_, _09565_, _09563_);
  nor (_09632_, _09631_, _09566_);
  and (_09633_, _09632_, _09630_);
  and (_09634_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_09635_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_09636_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [4]);
  and (_09637_, _09636_, _09635_);
  nor (_09638_, _09636_, _09635_);
  nor (_09639_, _09638_, _09637_);
  and (_09640_, _09639_, _09634_);
  nor (_09641_, _09639_, _09634_);
  nor (_09642_, _09641_, _09640_);
  nor (_09643_, _09632_, _09630_);
  nor (_09644_, _09643_, _09633_);
  and (_09645_, _09644_, _09642_);
  nor (_09646_, _09645_, _09633_);
  not (_09647_, _09646_);
  nor (_09648_, _09582_, _09580_);
  nor (_09649_, _09648_, _09583_);
  and (_09650_, _09649_, _09647_);
  not (_09651_, _09524_);
  nor (_09652_, _09640_, _09637_);
  nor (_09653_, _09652_, _09651_);
  and (_09654_, _09652_, _09651_);
  nor (_09655_, _09654_, _09653_);
  nor (_09656_, _09649_, _09647_);
  nor (_09657_, _09656_, _09650_);
  and (_09658_, _09657_, _09655_);
  nor (_09659_, _09658_, _09650_);
  not (_09660_, _09659_);
  nor (_09661_, _09599_, _09597_);
  nor (_09662_, _09661_, _09600_);
  and (_09663_, _09662_, _09660_);
  nor (_09664_, _09662_, _09660_);
  nor (_09665_, _09664_, _09663_);
  and (_09666_, _09665_, _09653_);
  nor (_09667_, _09666_, _09663_);
  nor (_09668_, _09607_, _09595_);
  nor (_09669_, _09668_, _09608_);
  not (_09670_, _09669_);
  nor (_09671_, _09670_, _09667_);
  and (_09672_, _09612_, _09609_);
  nor (_09673_, _09672_, _09613_);
  and (_09674_, _09673_, _09671_);
  nor (_09675_, _09615_, _09613_);
  nor (_09676_, _09675_, _09616_);
  nand (_09677_, _09676_, _09674_);
  or (_09678_, _09676_, _09674_);
  and (_09679_, _09678_, _09677_);
  and (_09680_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_09681_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_09682_, _09681_, _09680_);
  and (_09683_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [2]);
  nor (_09684_, _09681_, _09680_);
  nor (_09685_, _09684_, _09682_);
  and (_09686_, _09685_, _09683_);
  nor (_09687_, _09686_, _09682_);
  not (_09688_, _09687_);
  nor (_09689_, _09627_, _09625_);
  nor (_09690_, _09689_, _09628_);
  and (_09691_, _09690_, _09688_);
  and (_09692_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_09693_, _09692_, _09636_);
  and (_09694_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [3]);
  and (_09695_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_09696_, _09695_, _09694_);
  nor (_09698_, _09696_, _09693_);
  nor (_09699_, _09690_, _09688_);
  nor (_09701_, _09699_, _09691_);
  and (_09702_, _09701_, _09698_);
  nor (_09704_, _09702_, _09691_);
  not (_09705_, _09704_);
  nor (_09707_, _09644_, _09642_);
  nor (_09708_, _09707_, _09645_);
  and (_09710_, _09708_, _09705_);
  nor (_09711_, _09708_, _09705_);
  nor (_09713_, _09711_, _09710_);
  and (_09714_, _09713_, _09693_);
  nor (_09716_, _09714_, _09710_);
  not (_09717_, _09716_);
  nor (_09719_, _09657_, _09655_);
  nor (_09720_, _09719_, _09658_);
  and (_09722_, _09720_, _09717_);
  nor (_09723_, _09665_, _09653_);
  nor (_09725_, _09723_, _09666_);
  and (_09726_, _09725_, _09722_);
  and (_09728_, _09670_, _09667_);
  nor (_09729_, _09728_, _09671_);
  and (_09731_, _09729_, _09726_);
  nor (_09732_, _09673_, _09671_);
  nor (_09734_, _09732_, _09674_);
  and (_09735_, _09734_, _09731_);
  nor (_09736_, _09734_, _09731_);
  nor (_09737_, _09736_, _09735_);
  and (_09738_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_09739_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [1]);
  and (_09740_, _09739_, _09738_);
  and (_09741_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_09742_, _09739_, _09738_);
  nor (_09743_, _09742_, _09740_);
  and (_09744_, _09743_, _09741_);
  nor (_09745_, _09744_, _09740_);
  not (_09746_, _09745_);
  nor (_09747_, _09685_, _09683_);
  nor (_09748_, _09747_, _09686_);
  and (_09749_, _09748_, _09746_);
  nor (_09750_, _09748_, _09746_);
  nor (_09751_, _09750_, _09749_);
  and (_09752_, _09751_, _09692_);
  nor (_09753_, _09752_, _09749_);
  not (_09754_, _09753_);
  nor (_09755_, _09701_, _09698_);
  nor (_09756_, _09755_, _09702_);
  and (_09757_, _09756_, _09754_);
  nor (_09758_, _09713_, _09693_);
  nor (_09759_, _09758_, _09714_);
  and (_09760_, _09759_, _09757_);
  nor (_09761_, _09720_, _09717_);
  nor (_09762_, _09761_, _09722_);
  and (_09763_, _09762_, _09760_);
  nor (_09764_, _09725_, _09722_);
  nor (_09765_, _09764_, _09726_);
  and (_09766_, _09765_, _09763_);
  nor (_09767_, _09729_, _09726_);
  nor (_09768_, _09767_, _09731_);
  and (_09769_, _09768_, _09766_);
  and (_09770_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  and (_09771_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  and (_09772_, _09771_, _09770_);
  nor (_09773_, _09743_, _09741_);
  nor (_09774_, _09773_, _09744_);
  and (_09775_, _09774_, _09772_);
  nor (_09776_, _09751_, _09692_);
  nor (_09777_, _09776_, _09752_);
  and (_09778_, _09777_, _09775_);
  nor (_09779_, _09756_, _09754_);
  nor (_09780_, _09779_, _09757_);
  and (_09781_, _09780_, _09778_);
  nor (_09782_, _09759_, _09757_);
  nor (_09783_, _09782_, _09760_);
  and (_09784_, _09783_, _09781_);
  nor (_09785_, _09762_, _09760_);
  nor (_09786_, _09785_, _09763_);
  and (_09787_, _09786_, _09784_);
  nor (_09788_, _09765_, _09763_);
  nor (_09789_, _09788_, _09766_);
  and (_09790_, _09789_, _09787_);
  nor (_09791_, _09768_, _09766_);
  nor (_09793_, _09791_, _09769_);
  and (_09795_, _09793_, _09790_);
  nor (_09796_, _09795_, _09769_);
  not (_09798_, _09796_);
  and (_09799_, _09798_, _09737_);
  or (_09801_, _09799_, _09735_);
  nand (_09802_, _09801_, _09679_);
  and (_09804_, _09802_, _09677_);
  not (_09805_, _09804_);
  and (_09807_, _09805_, _09621_);
  or (_09808_, _09807_, _09619_);
  or (_09810_, _09559_, _09557_);
  and (_09811_, _09810_, _09560_);
  nand (_09813_, _09811_, _09808_);
  and (_09814_, _09813_, _09560_);
  nor (_09816_, _09814_, _09493_);
  or (_09817_, _09816_, _09492_);
  and (_09819_, \oc8051_golden_model_1.ACC [7], \oc8051_golden_model_1.B [7]);
  not (_09820_, _09819_);
  nor (_09822_, _09820_, _09444_);
  nor (_09823_, _09822_, _09476_);
  nor (_09825_, _09482_, _09479_);
  nor (_09826_, _09825_, _09823_);
  and (_09828_, _09825_, _09823_);
  nor (_09829_, _09828_, _09826_);
  nor (_09830_, _09489_, _09486_);
  not (_09831_, _09830_);
  and (_09832_, _09831_, _09829_);
  nor (_09833_, _09831_, _09829_);
  nor (_09834_, _09833_, _09832_);
  and (_09835_, _09834_, _09817_);
  or (_09836_, _09826_, _09473_);
  or (_09837_, _09836_, _09832_);
  or (_09838_, _09837_, _09835_);
  or (_09839_, _09838_, _09301_);
  and (_09840_, _09839_, _06140_);
  and (_09841_, _09840_, _09300_);
  not (_09842_, _06132_);
  and (_09843_, _08587_, _08420_);
  or (_09844_, _09843_, _09267_);
  and (_09845_, _09844_, _06139_);
  or (_09846_, _09845_, _09842_);
  or (_09847_, _09846_, _09841_);
  and (_09848_, _09847_, _09266_);
  or (_09849_, _09848_, _06116_);
  and (_09850_, _08535_, _07841_);
  or (_09851_, _09263_, _06117_);
  or (_09852_, _09851_, _09850_);
  and (_09853_, _09852_, _06114_);
  and (_09854_, _09853_, _09849_);
  and (_09855_, _06294_, _05781_);
  and (_09856_, _08782_, _07841_);
  or (_09857_, _09856_, _09263_);
  and (_09858_, _09857_, _05787_);
  or (_09859_, _09858_, _09855_);
  or (_09860_, _09859_, _09854_);
  not (_09861_, _09855_);
  nor (_09862_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_09863_, _09862_, _09307_);
  not (_09864_, \oc8051_golden_model_1.B [1]);
  nor (_09865_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor (_09866_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and (_09867_, _09866_, _09865_);
  and (_09868_, _09867_, _09864_);
  nor (_09869_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not (_09870_, _09869_);
  and (_09871_, \oc8051_golden_model_1.B [0], _08430_);
  nor (_09872_, _09871_, _09870_);
  and (_09873_, _09872_, _09868_);
  and (_09874_, _09873_, _09863_);
  or (_09875_, _09873_, _08430_);
  not (_09876_, \oc8051_golden_model_1.B [4]);
  not (_09877_, \oc8051_golden_model_1.B [5]);
  nor (_09878_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_09879_, _09878_, _09877_);
  and (_09880_, _09879_, _09876_);
  nor (_09881_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.B [2]);
  and (_09882_, _09881_, _09880_);
  not (_09883_, \oc8051_golden_model_1.ACC [6]);
  and (_09884_, \oc8051_golden_model_1.B [0], _09883_);
  nor (_09885_, _09884_, _08430_);
  nor (_09886_, _09885_, _09864_);
  not (_09887_, _09886_);
  and (_09888_, _09887_, _09882_);
  nor (_09889_, _09888_, _09875_);
  nor (_09890_, _09889_, _09874_);
  and (_09891_, _09888_, \oc8051_golden_model_1.B [0]);
  nor (_09892_, _09891_, _09883_);
  and (_09893_, _09892_, _09864_);
  nor (_09894_, _09892_, _09864_);
  nor (_09895_, _09894_, _09893_);
  nor (_09896_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  nor (_09897_, _09896_, _09494_);
  nor (_09898_, _09897_, \oc8051_golden_model_1.ACC [4]);
  not (_09899_, \oc8051_golden_model_1.B [0]);
  and (_09900_, \oc8051_golden_model_1.ACC [4], _09899_);
  nor (_09901_, _09900_, \oc8051_golden_model_1.ACC [5]);
  not (_09902_, \oc8051_golden_model_1.ACC [4]);
  and (_09903_, _09902_, \oc8051_golden_model_1.B [0]);
  nor (_09904_, _09903_, _09901_);
  nor (_09905_, _09904_, _09898_);
  not (_09906_, _09905_);
  and (_09907_, _09906_, _09895_);
  nor (_09908_, _09890_, \oc8051_golden_model_1.B [2]);
  nor (_09909_, _09908_, _09893_);
  not (_09910_, _09909_);
  nor (_09911_, _09910_, _09907_);
  and (_09912_, \oc8051_golden_model_1.B [2], _08430_);
  nor (_09913_, _09912_, \oc8051_golden_model_1.B [7]);
  and (_09914_, _09913_, _09867_);
  not (_09915_, _09914_);
  nor (_09916_, _09915_, _09911_);
  nor (_09917_, _09916_, _09890_);
  nor (_09918_, _09917_, _09874_);
  not (_09919_, \oc8051_golden_model_1.B [2]);
  nor (_09920_, _09906_, _09895_);
  nor (_09921_, _09920_, _09907_);
  not (_09922_, _09921_);
  and (_09923_, _09922_, _09916_);
  nor (_09924_, _09916_, _09892_);
  nor (_09925_, _09924_, _09923_);
  and (_09926_, _09925_, _09919_);
  nor (_09927_, _09925_, _09919_);
  nor (_09928_, _09927_, _09926_);
  not (_09929_, _09928_);
  not (_09930_, \oc8051_golden_model_1.ACC [5]);
  nor (_09931_, _09916_, _09930_);
  and (_09932_, _09916_, _09897_);
  or (_09933_, _09932_, _09931_);
  and (_09934_, _09933_, _09864_);
  nor (_09935_, _09933_, _09864_);
  nor (_09936_, _09935_, _09903_);
  nor (_09937_, _09936_, _09934_);
  nor (_09938_, _09937_, _09929_);
  nor (_09939_, _09918_, \oc8051_golden_model_1.B [3]);
  nor (_09940_, _09939_, _09926_);
  not (_09941_, _09940_);
  nor (_09942_, _09941_, _09938_);
  not (_09943_, _09942_);
  and (_09944_, \oc8051_golden_model_1.B [3], _08430_);
  not (_09945_, _09944_);
  and (_09946_, _09945_, _09880_);
  and (_09947_, _09946_, _09943_);
  nor (_09948_, _09947_, _09918_);
  nor (_09949_, _09948_, _09874_);
  nor (_09950_, _09949_, \oc8051_golden_model_1.B [4]);
  not (_09951_, \oc8051_golden_model_1.B [3]);
  not (_09952_, _09947_);
  and (_09953_, _09937_, _09929_);
  nor (_09954_, _09953_, _09938_);
  nor (_09955_, _09954_, _09952_);
  nor (_09956_, _09947_, _09925_);
  nor (_09957_, _09956_, _09955_);
  and (_09958_, _09957_, _09951_);
  nor (_09959_, _09957_, _09951_);
  nor (_09960_, _09959_, _09958_);
  not (_09961_, _09960_);
  nor (_09962_, _09947_, _09933_);
  nor (_09963_, _09935_, _09934_);
  and (_09964_, _09963_, _09903_);
  nor (_09965_, _09963_, _09903_);
  nor (_09966_, _09965_, _09964_);
  and (_09967_, _09966_, _09947_);
  or (_09968_, _09967_, _09962_);
  nor (_09969_, _09968_, \oc8051_golden_model_1.B [2]);
  and (_09970_, _09968_, \oc8051_golden_model_1.B [2]);
  nor (_09971_, _09903_, _09900_);
  and (_09972_, _09947_, _09971_);
  nor (_09973_, _09947_, \oc8051_golden_model_1.ACC [4]);
  nor (_09974_, _09973_, _09972_);
  and (_09975_, _09974_, _09864_);
  nor (_09976_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_09977_, _09976_, _09680_);
  nor (_09978_, _09977_, \oc8051_golden_model_1.ACC [2]);
  and (_09979_, _09899_, \oc8051_golden_model_1.ACC [2]);
  nor (_09980_, _09979_, \oc8051_golden_model_1.ACC [3]);
  not (_09981_, \oc8051_golden_model_1.ACC [2]);
  and (_09982_, \oc8051_golden_model_1.B [0], _09981_);
  nor (_09983_, _09982_, _09980_);
  nor (_09984_, _09983_, _09978_);
  not (_09985_, _09984_);
  nor (_09986_, _09974_, _09864_);
  nor (_09987_, _09986_, _09975_);
  and (_09988_, _09987_, _09985_);
  nor (_09989_, _09988_, _09975_);
  nor (_09990_, _09989_, _09970_);
  nor (_09991_, _09990_, _09969_);
  nor (_09992_, _09991_, _09961_);
  or (_09993_, _09992_, _09958_);
  nor (_09994_, _09993_, _09950_);
  and (_09995_, _09879_, \oc8051_golden_model_1.ACC [7]);
  or (_09996_, _09995_, _09880_);
  not (_09997_, _09996_);
  nor (_09998_, _09997_, _09994_);
  nor (_09999_, _09998_, _09949_);
  nor (_10000_, _09999_, _09874_);
  and (_10001_, _09991_, _09961_);
  nor (_10002_, _10001_, _09992_);
  not (_10003_, _10002_);
  and (_10004_, _10003_, _09998_);
  nor (_10005_, _09998_, _09957_);
  nor (_10006_, _10005_, _10004_);
  and (_10007_, _10006_, _09876_);
  nor (_10008_, _10006_, _09876_);
  nor (_10009_, _10008_, _10007_);
  not (_10010_, _10009_);
  nor (_10011_, _09998_, _09968_);
  nor (_10012_, _09970_, _09969_);
  and (_10013_, _10012_, _09989_);
  nor (_10014_, _10012_, _09989_);
  nor (_10015_, _10014_, _10013_);
  not (_10016_, _10015_);
  and (_10017_, _10016_, _09998_);
  nor (_10018_, _10017_, _10011_);
  nor (_10019_, _10018_, \oc8051_golden_model_1.B [3]);
  and (_10020_, _10018_, \oc8051_golden_model_1.B [3]);
  nor (_10021_, _09987_, _09985_);
  nor (_10022_, _10021_, _09988_);
  not (_10023_, _10022_);
  and (_10024_, _10023_, _09998_);
  nor (_10025_, _09998_, _09974_);
  nor (_10026_, _10025_, _10024_);
  and (_10027_, _10026_, _09919_);
  not (_10028_, \oc8051_golden_model_1.ACC [3]);
  nor (_10029_, _09998_, _10028_);
  and (_10030_, _09998_, _09977_);
  or (_10031_, _10030_, _10029_);
  and (_10032_, _10031_, _09864_);
  nor (_10033_, _10031_, _09864_);
  nor (_10034_, _10033_, _09982_);
  nor (_10035_, _10034_, _10032_);
  nor (_10036_, _10026_, _09919_);
  nor (_10037_, _10036_, _10027_);
  not (_10038_, _10037_);
  nor (_10039_, _10038_, _10035_);
  nor (_10040_, _10039_, _10027_);
  nor (_10041_, _10040_, _10020_);
  nor (_10042_, _10041_, _10019_);
  nor (_10043_, _10042_, _10010_);
  nor (_10044_, _10000_, \oc8051_golden_model_1.B [5]);
  nor (_10045_, _10044_, _10007_);
  not (_10046_, _10045_);
  nor (_10047_, _10046_, _10043_);
  not (_10048_, _10047_);
  not (_10049_, _09878_);
  and (_10050_, \oc8051_golden_model_1.B [5], _08430_);
  nor (_10051_, _10050_, _10049_);
  and (_10052_, _10051_, _10048_);
  nor (_10053_, _10052_, _10000_);
  nor (_10054_, _10053_, _09874_);
  not (_10055_, _10052_);
  and (_10056_, _10042_, _10010_);
  nor (_10057_, _10056_, _10043_);
  nor (_10058_, _10057_, _10055_);
  nor (_10059_, _10052_, _10006_);
  nor (_10060_, _10059_, _10058_);
  and (_10061_, _10060_, _09877_);
  nor (_10062_, _10060_, _09877_);
  nor (_10063_, _10062_, _10061_);
  not (_10064_, _10063_);
  nor (_10065_, _10052_, _10018_);
  nor (_10066_, _10020_, _10019_);
  nor (_10067_, _10066_, _10040_);
  and (_10068_, _10066_, _10040_);
  or (_10069_, _10068_, _10067_);
  and (_10070_, _10069_, _10052_);
  or (_10071_, _10070_, _10065_);
  and (_10072_, _10071_, _09876_);
  nor (_10073_, _10071_, _09876_);
  and (_10074_, _10038_, _10035_);
  nor (_10075_, _10074_, _10039_);
  nor (_10076_, _10075_, _10055_);
  nor (_10077_, _10052_, _10026_);
  nor (_10078_, _10077_, _10076_);
  and (_10079_, _10078_, _09951_);
  nor (_10080_, _10033_, _10032_);
  nor (_10081_, _10080_, _09982_);
  and (_10082_, _10080_, _09982_);
  or (_10083_, _10082_, _10081_);
  nor (_10084_, _10083_, _10055_);
  nor (_10085_, _10052_, _10031_);
  nor (_10086_, _10085_, _10084_);
  and (_10087_, _10086_, _09919_);
  nor (_10088_, _10086_, _09919_);
  nor (_10089_, _09982_, _09979_);
  and (_10090_, _10052_, _10089_);
  nor (_10091_, _10052_, \oc8051_golden_model_1.ACC [2]);
  nor (_10092_, _10091_, _10090_);
  and (_10093_, _10092_, _09864_);
  and (_10094_, _05887_, \oc8051_golden_model_1.B [0]);
  not (_10095_, _10094_);
  nor (_10096_, _10092_, _09864_);
  nor (_10097_, _10096_, _10093_);
  and (_10098_, _10097_, _10095_);
  nor (_10099_, _10098_, _10093_);
  nor (_10100_, _10099_, _10088_);
  nor (_10101_, _10100_, _10087_);
  nor (_10102_, _10078_, _09951_);
  nor (_10103_, _10102_, _10079_);
  not (_10104_, _10103_);
  nor (_10105_, _10104_, _10101_);
  nor (_10106_, _10105_, _10079_);
  nor (_10107_, _10106_, _10073_);
  nor (_10108_, _10107_, _10072_);
  nor (_10109_, _10108_, _10064_);
  nor (_10110_, _10054_, \oc8051_golden_model_1.B [6]);
  or (_10111_, _10110_, _10061_);
  or (_10112_, _10111_, _10109_);
  and (_10113_, \oc8051_golden_model_1.B [6], _08430_);
  nor (_10114_, _10113_, \oc8051_golden_model_1.B [7]);
  and (_10115_, _10114_, _10112_);
  nor (_10116_, _10115_, _10054_);
  or (_10117_, _10116_, _09874_);
  nor (_10118_, _10117_, \oc8051_golden_model_1.B [7]);
  nor (_10119_, _10118_, _09819_);
  not (_10120_, \oc8051_golden_model_1.B [6]);
  and (_10121_, _10108_, _10064_);
  nor (_10122_, _10121_, _10109_);
  not (_10123_, _10122_);
  and (_10124_, _10123_, _10115_);
  nor (_10125_, _10115_, _10060_);
  nor (_10126_, _10125_, _10124_);
  nor (_10127_, _10126_, _10120_);
  not (_10128_, _10127_);
  nor (_10129_, _10128_, _10119_);
  nor (_10130_, _10088_, _10087_);
  nor (_10131_, _10130_, _10099_);
  and (_10132_, _10130_, _10099_);
  or (_10133_, _10132_, _10131_);
  not (_10134_, _10133_);
  and (_10135_, _10134_, _10115_);
  nor (_10136_, _10115_, _10086_);
  nor (_10137_, _10136_, _10135_);
  and (_10138_, _10137_, _09951_);
  nor (_10139_, _10137_, _09951_);
  nor (_10140_, _10139_, _10138_);
  nor (_10141_, _10097_, _10095_);
  nor (_10142_, _10141_, _10098_);
  and (_10143_, _10142_, _10115_);
  not (_10144_, _10092_);
  nor (_10145_, _10115_, _10144_);
  nor (_10146_, _10145_, _10143_);
  and (_10147_, _10146_, \oc8051_golden_model_1.B [2]);
  nor (_10148_, _10146_, \oc8051_golden_model_1.B [2]);
  nor (_10149_, _10148_, _10147_);
  and (_10150_, _10149_, _10140_);
  nor (_10151_, _10115_, \oc8051_golden_model_1.ACC [1]);
  nor (_10152_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  or (_10153_, _10152_, _09770_);
  and (_10154_, _10115_, _10153_);
  nor (_10155_, _10154_, _10151_);
  and (_10156_, _10155_, _09864_);
  nor (_10157_, _10155_, _09864_);
  and (_10158_, _09899_, \oc8051_golden_model_1.ACC [0]);
  not (_10159_, _10158_);
  nor (_10160_, _10159_, _10157_);
  nor (_10161_, _10160_, _10156_);
  and (_10162_, _10161_, _10150_);
  not (_10163_, _10162_);
  and (_10164_, _10147_, _10140_);
  nor (_10165_, _10164_, _10139_);
  and (_10166_, _10165_, _10163_);
  and (_10167_, _10126_, _10120_);
  nor (_10168_, _10167_, _10127_);
  not (_10169_, _10168_);
  nor (_10170_, _10169_, _10119_);
  and (_10171_, _10104_, _10101_);
  or (_10172_, _10171_, _10105_);
  and (_10173_, _10172_, _10115_);
  nor (_10174_, _10115_, _10078_);
  nor (_10175_, _10174_, _10173_);
  nor (_10176_, _10175_, _09876_);
  and (_10177_, _10175_, _09876_);
  nor (_10178_, _10177_, _10176_);
  nor (_10179_, _10073_, _10072_);
  nor (_10180_, _10179_, _10106_);
  and (_10181_, _10179_, _10106_);
  or (_10182_, _10181_, _10180_);
  not (_10183_, _10182_);
  and (_10184_, _10183_, _10115_);
  nor (_10185_, _10115_, _10071_);
  nor (_10186_, _10185_, _10184_);
  nor (_10187_, _10186_, _09877_);
  and (_10188_, _10186_, _09877_);
  nor (_10189_, _10188_, _10187_);
  and (_10190_, _10189_, _10178_);
  and (_10191_, _10190_, _10170_);
  not (_10192_, _10191_);
  nor (_10193_, _10192_, _10166_);
  and (_10194_, _10054_, \oc8051_golden_model_1.B [7]);
  and (_10195_, _10189_, _10176_);
  nor (_10196_, _10195_, _10187_);
  not (_10197_, _10196_);
  and (_10198_, _10197_, _10170_);
  or (_10199_, _10198_, _10194_);
  or (_10200_, _10199_, _10193_);
  nor (_10201_, _10200_, _10129_);
  and (_10202_, \oc8051_golden_model_1.B [0], _05855_);
  not (_10203_, _10202_);
  nor (_10204_, _10157_, _10156_);
  and (_10205_, _10204_, _10203_);
  and (_10206_, _10205_, _10159_);
  and (_10207_, _10206_, _10150_);
  and (_10208_, _10207_, _10191_);
  nor (_10209_, _10208_, _10201_);
  and (_10210_, _10209_, _10117_);
  or (_10211_, _10210_, _09874_);
  or (_10212_, _10211_, _09861_);
  and (_10213_, _10212_, _06298_);
  and (_10214_, _10213_, _09860_);
  and (_10215_, _08802_, _07841_);
  or (_10216_, _10215_, _09263_);
  and (_10217_, _10216_, _06297_);
  and (_10218_, _08607_, _07841_);
  or (_10219_, _10218_, _09263_);
  and (_10220_, _10219_, _06110_);
  or (_10221_, _10220_, _06402_);
  or (_10222_, _10221_, _10217_);
  or (_10223_, _10222_, _10214_);
  and (_10224_, _08810_, _07841_);
  or (_10225_, _09263_, _07125_);
  or (_10226_, _10225_, _10224_);
  and (_10227_, _10226_, _07132_);
  and (_10228_, _10227_, _10223_);
  or (_10229_, _09263_, _07926_);
  and (_10230_, _10219_, _06306_);
  and (_10231_, _10230_, _10229_);
  or (_10232_, _10231_, _10228_);
  and (_10233_, _10232_, _07130_);
  and (_10234_, _09275_, _06411_);
  and (_10235_, _10234_, _10229_);
  or (_10236_, _10235_, _06303_);
  or (_10237_, _10236_, _10233_);
  and (_10238_, _08801_, _07841_);
  or (_10239_, _09263_, _08819_);
  or (_10240_, _10239_, _10238_);
  and (_10241_, _10240_, _08824_);
  and (_10242_, _10241_, _10237_);
  not (_10243_, _07841_);
  nor (_10244_, _08809_, _10243_);
  or (_10245_, _10244_, _09263_);
  and (_10246_, _10245_, _06396_);
  or (_10247_, _10246_, _06433_);
  or (_10248_, _10247_, _10242_);
  or (_10249_, _09272_, _06829_);
  and (_10250_, _10249_, _05749_);
  and (_10251_, _10250_, _10248_);
  and (_10252_, _09269_, _05748_);
  or (_10253_, _10252_, _06440_);
  or (_10254_, _10253_, _10251_);
  and (_10255_, _08345_, _07841_);
  or (_10256_, _09263_, _06444_);
  or (_10257_, _10256_, _10255_);
  and (_10258_, _10257_, _01317_);
  and (_10259_, _10258_, _10254_);
  or (_10260_, _10259_, _09262_);
  and (_40980_, _10260_, _43100_);
  nor (_10261_, _01317_, _08430_);
  and (_10262_, _05825_, _06302_);
  nand (_10263_, _10262_, _09883_);
  and (_10264_, _06294_, _05825_);
  not (_10265_, _10264_);
  nor (_10266_, _08014_, _09883_);
  not (_10267_, _10266_);
  nor (_10268_, _08103_, _09930_);
  and (_10269_, _08103_, _09930_);
  nor (_10270_, _08338_, _09902_);
  not (_10271_, _10270_);
  nor (_10272_, _08139_, _10028_);
  and (_10273_, _08139_, _10028_);
  nor (_10274_, _08247_, _09981_);
  nor (_10275_, _08175_, _05887_);
  and (_10276_, _08211_, \oc8051_golden_model_1.ACC [0]);
  and (_10277_, _08175_, _05887_);
  nor (_10278_, _10277_, _10275_);
  and (_10279_, _10278_, _10276_);
  nor (_10280_, _10279_, _10275_);
  and (_10281_, _08247_, _09981_);
  nor (_10282_, _10281_, _10274_);
  not (_10283_, _10282_);
  nor (_10284_, _10283_, _10280_);
  nor (_10285_, _10284_, _10274_);
  nor (_10286_, _10285_, _10273_);
  or (_10287_, _10286_, _10272_);
  and (_10288_, _08338_, _09902_);
  nor (_10289_, _10288_, _10270_);
  nand (_10290_, _10289_, _10287_);
  and (_10291_, _10290_, _10271_);
  nor (_10292_, _10291_, _10269_);
  or (_10293_, _10292_, _10268_);
  and (_10294_, _08014_, _09883_);
  nor (_10295_, _10294_, _10266_);
  nand (_10296_, _10295_, _10293_);
  and (_10297_, _10296_, _10267_);
  nor (_10298_, _10297_, _08810_);
  and (_10299_, _10297_, _08810_);
  or (_10300_, _10299_, _10298_);
  and (_10301_, _10300_, _06169_);
  and (_10302_, _09200_, \oc8051_golden_model_1.PSW [7]);
  nor (_10303_, _10302_, _09194_);
  and (_10304_, _10302_, _09194_);
  nor (_10305_, _10304_, _10303_);
  and (_10306_, _10305_, \oc8051_golden_model_1.ACC [7]);
  nor (_10307_, _10305_, \oc8051_golden_model_1.ACC [7]);
  nor (_10308_, _10307_, _10306_);
  and (_10309_, _09199_, \oc8051_golden_model_1.PSW [7]);
  nor (_10310_, _10309_, _08012_);
  nor (_10311_, _10310_, _10302_);
  nand (_10312_, _10311_, \oc8051_golden_model_1.ACC [6]);
  nor (_10313_, _10311_, _09883_);
  and (_10314_, _10311_, _09883_);
  nor (_10315_, _10314_, _10313_);
  not (_10316_, _10315_);
  and (_10317_, _09198_, \oc8051_golden_model_1.PSW [7]);
  nor (_10318_, _10317_, _08101_);
  nor (_10319_, _10318_, _10309_);
  and (_10320_, _10319_, \oc8051_golden_model_1.ACC [5]);
  nor (_10321_, _10319_, _09930_);
  and (_10322_, _10319_, _09930_);
  nor (_10323_, _10322_, _10321_);
  and (_10324_, _09197_, \oc8051_golden_model_1.PSW [7]);
  nor (_10325_, _10324_, _08336_);
  nor (_10326_, _10325_, _10317_);
  nand (_10327_, _10326_, \oc8051_golden_model_1.ACC [4]);
  nor (_10328_, _10326_, _09902_);
  and (_10329_, _10326_, _09902_);
  or (_10330_, _10329_, _10328_);
  and (_10331_, _09196_, \oc8051_golden_model_1.PSW [7]);
  nor (_10332_, _10331_, _07544_);
  nor (_10333_, _10332_, _10324_);
  and (_10334_, _10333_, \oc8051_golden_model_1.ACC [3]);
  nor (_10335_, _10333_, _10028_);
  and (_10336_, _10333_, _10028_);
  nor (_10337_, _10336_, _10335_);
  and (_10338_, _09195_, \oc8051_golden_model_1.PSW [7]);
  nor (_10339_, _10338_, _07708_);
  nor (_10340_, _10339_, _10331_);
  and (_10341_, _10340_, \oc8051_golden_model_1.ACC [2]);
  nor (_10342_, _10340_, _09981_);
  and (_10343_, _10340_, _09981_);
  nor (_10344_, _10343_, _10342_);
  and (_10345_, _07049_, \oc8051_golden_model_1.PSW [7]);
  nor (_10346_, _10345_, _07306_);
  nor (_10347_, _10346_, _10338_);
  and (_10348_, _10347_, \oc8051_golden_model_1.ACC [1]);
  and (_10349_, _10347_, _05887_);
  nor (_10350_, _10347_, _05887_);
  nor (_10351_, _10350_, _10349_);
  not (_10352_, _10351_);
  nor (_10353_, _07049_, \oc8051_golden_model_1.PSW [7]);
  nor (_10354_, _10353_, _10345_);
  and (_10355_, _10354_, \oc8051_golden_model_1.ACC [0]);
  and (_10356_, _10355_, _10352_);
  nor (_10357_, _10356_, _10348_);
  nor (_10358_, _10357_, _10344_);
  nor (_10359_, _10358_, _10341_);
  nor (_10360_, _10359_, _10337_);
  or (_10361_, _10360_, _10334_);
  nand (_10362_, _10361_, _10330_);
  and (_10363_, _10362_, _10327_);
  nor (_10364_, _10363_, _10323_);
  or (_10365_, _10364_, _10320_);
  nand (_10366_, _10365_, _10316_);
  and (_10367_, _10366_, _10312_);
  nor (_10368_, _10367_, _10308_);
  and (_10369_, _10367_, _10308_);
  nor (_10370_, _10369_, _10368_);
  and (_10371_, _06123_, _06300_);
  nor (_10372_, _10371_, _06523_);
  and (_10373_, _06119_, _06300_);
  not (_10374_, _10373_);
  not (_10375_, _06794_);
  and (_10376_, _06957_, _06300_);
  nor (_10377_, _10376_, _06795_);
  and (_10378_, _10377_, _10375_);
  and (_10379_, _10378_, _10374_);
  and (_10380_, _10379_, _10372_);
  or (_10381_, _10380_, _10370_);
  or (_10382_, _06039_, _05802_);
  nor (_10383_, _07809_, _08430_);
  and (_10384_, _07923_, _07809_);
  or (_10385_, _10384_, _10383_);
  or (_10386_, _10385_, _06132_);
  and (_10387_, _06294_, _05790_);
  not (_10388_, _10387_);
  and (_10389_, _08211_, \oc8051_golden_model_1.PSW [7]);
  and (_10390_, _10389_, _08176_);
  and (_10391_, _10390_, _08248_);
  and (_10392_, _10391_, _08140_);
  and (_10393_, _10392_, _08339_);
  and (_10394_, _10393_, _08104_);
  and (_10395_, _10394_, _08015_);
  nor (_10396_, _10395_, _07925_);
  and (_10397_, _10395_, _07925_);
  nor (_10398_, _10397_, _10396_);
  and (_10399_, _10398_, \oc8051_golden_model_1.ACC [7]);
  nor (_10400_, _10398_, \oc8051_golden_model_1.ACC [7]);
  nor (_10401_, _10400_, _10399_);
  not (_10402_, _10401_);
  nor (_10403_, _10394_, _08015_);
  nor (_10404_, _10403_, _10395_);
  nor (_10405_, _10404_, _09883_);
  nor (_10406_, _10393_, _08104_);
  nor (_10407_, _10406_, _10394_);
  nor (_10408_, _10407_, _09930_);
  and (_10409_, _10407_, _09930_);
  nor (_10410_, _10409_, _10408_);
  not (_10411_, _10410_);
  nor (_10412_, _10392_, _08339_);
  nor (_10413_, _10412_, _10393_);
  nor (_10414_, _10413_, _09902_);
  and (_10415_, _10413_, _09902_);
  or (_10416_, _10415_, _10414_);
  or (_10417_, _10416_, _10411_);
  nor (_10418_, _10391_, _08140_);
  nor (_10419_, _10418_, _10392_);
  nor (_10420_, _10419_, _10028_);
  and (_10421_, _10419_, _10028_);
  nor (_10422_, _10421_, _10420_);
  nor (_10423_, _10390_, _08248_);
  nor (_10424_, _10423_, _10391_);
  nor (_10425_, _10424_, _09981_);
  and (_10426_, _10424_, _09981_);
  nor (_10427_, _10426_, _10425_);
  and (_10428_, _10427_, _10422_);
  nor (_10429_, _10389_, _08176_);
  nor (_10430_, _10429_, _10390_);
  nor (_10431_, _10430_, _05887_);
  and (_10432_, _10430_, _05887_);
  nor (_10433_, _08211_, \oc8051_golden_model_1.PSW [7]);
  nor (_10434_, _10433_, _10389_);
  and (_10435_, _10434_, _05855_);
  nor (_10436_, _10435_, _10432_);
  or (_10437_, _10436_, _10431_);
  nand (_10438_, _10437_, _10428_);
  nor (_10439_, _10425_, _10420_);
  or (_10440_, _10439_, _10421_);
  and (_10441_, _10440_, _10438_);
  nor (_10442_, _10441_, _10417_);
  nor (_10443_, _10414_, _10408_);
  nor (_10444_, _10443_, _10409_);
  nor (_10445_, _10444_, _10442_);
  and (_10446_, _10404_, _09883_);
  nor (_10447_, _10405_, _10446_);
  not (_10448_, _10447_);
  nor (_10449_, _10448_, _10445_);
  or (_10450_, _10449_, _10405_);
  and (_10451_, _10450_, _10402_);
  nor (_10452_, _10450_, _10402_);
  or (_10453_, _10452_, _10451_);
  or (_10454_, _10453_, _06265_);
  and (_10455_, _10454_, _10388_);
  not (_10456_, _06529_);
  nor (_10457_, _07678_, _06538_);
  and (_10458_, _10457_, _10456_);
  or (_10459_, _10458_, _07923_);
  nor (_10460_, _08409_, _08430_);
  and (_10461_, _08552_, _08409_);
  or (_10462_, _10461_, _10460_);
  or (_10463_, _10462_, _06157_);
  and (_10464_, _10463_, _07075_);
  not (_10465_, _06658_);
  nor (_10466_, _06119_, _06284_);
  nor (_10467_, _10466_, _05771_);
  nor (_10468_, _10467_, _10465_);
  nor (_10469_, _06129_, _05771_);
  not (_10470_, _10469_);
  and (_10471_, _10470_, _10468_);
  or (_10472_, _10471_, _07923_);
  and (_10473_, _06294_, _06222_);
  not (_10474_, _10473_);
  nor (_10475_, _06653_, _08430_);
  and (_10476_, _06653_, _08430_);
  nor (_10477_, _10476_, _10475_);
  nand (_10478_, _10477_, _10471_);
  and (_10479_, _10478_, _10474_);
  and (_10480_, _10479_, _10472_);
  and (_10481_, _10473_, _08535_);
  or (_10482_, _10481_, _10480_);
  not (_10483_, _05772_);
  nor (_10484_, _06160_, _10483_);
  and (_10485_, _10484_, _10482_);
  and (_10486_, _08548_, _07809_);
  or (_10487_, _10486_, _10383_);
  and (_10488_, _10487_, _06160_);
  or (_10489_, _10488_, _10485_);
  and (_10490_, _06294_, _06155_);
  not (_10491_, _10490_);
  and (_10492_, _10491_, _10489_);
  nor (_10493_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [2]);
  nor (_10494_, _10493_, _10028_);
  and (_10495_, _10494_, \oc8051_golden_model_1.ACC [4]);
  and (_10496_, _10495_, \oc8051_golden_model_1.ACC [5]);
  and (_10497_, _10496_, \oc8051_golden_model_1.ACC [6]);
  and (_10498_, _10497_, \oc8051_golden_model_1.ACC [7]);
  nor (_10499_, _10497_, \oc8051_golden_model_1.ACC [7]);
  nor (_10500_, _10499_, _10498_);
  nor (_10501_, _10495_, \oc8051_golden_model_1.ACC [5]);
  nor (_10502_, _10501_, _10496_);
  nor (_10503_, _10496_, \oc8051_golden_model_1.ACC [6]);
  nor (_10504_, _10503_, _10497_);
  nor (_10505_, _10504_, _10502_);
  not (_10506_, _10505_);
  and (_10507_, _10506_, _10500_);
  or (_10508_, _10498_, \oc8051_golden_model_1.PSW [7]);
  and (_10509_, _10508_, _10506_);
  nor (_10510_, _10509_, _10500_);
  nor (_10511_, _10510_, _10507_);
  and (_10512_, _10511_, _10490_);
  or (_10513_, _10512_, _06156_);
  or (_10514_, _10513_, _10492_);
  and (_10515_, _10514_, _10464_);
  not (_10516_, _10458_);
  and (_10517_, _10385_, _06217_);
  or (_10518_, _10517_, _10516_);
  or (_10519_, _10518_, _10515_);
  and (_10520_, _10519_, _10459_);
  or (_10521_, _10520_, _07081_);
  or (_10522_, _08535_, _07082_);
  and (_10523_, _10522_, _06229_);
  and (_10524_, _10523_, _10521_);
  and (_10525_, _06294_, _06150_);
  nor (_10526_, _07925_, _06229_);
  or (_10527_, _10526_, _10525_);
  or (_10528_, _10527_, _10524_);
  nand (_10529_, _10525_, _10028_);
  and (_10530_, _10529_, _10528_);
  or (_10531_, _10530_, _06152_);
  and (_10532_, _08426_, _08409_);
  or (_10533_, _10532_, _10460_);
  or (_10534_, _10533_, _06153_);
  and (_10535_, _10534_, _06146_);
  and (_10536_, _10535_, _10531_);
  or (_10537_, _10460_, _08568_);
  and (_10538_, _10462_, _06145_);
  and (_10539_, _10538_, _10537_);
  or (_10540_, _10539_, _09295_);
  or (_10541_, _10540_, _10536_);
  nor (_10542_, _09789_, _09787_);
  nor (_10543_, _10542_, _09790_);
  or (_10544_, _10543_, _09301_);
  and (_10545_, _06273_, _05790_);
  not (_10546_, _10545_);
  and (_10547_, _06125_, _05790_);
  nor (_10548_, _10547_, _06536_);
  and (_10549_, _06118_, _05790_);
  or (_10550_, _06971_, _06276_);
  and (_10551_, _10550_, _10549_);
  not (_10552_, _10551_);
  and (_10553_, _10552_, _10548_);
  and (_10554_, _10553_, _10546_);
  and (_10555_, _10554_, _10544_);
  and (_10556_, _10555_, _10541_);
  not (_10557_, _10554_);
  not (_10558_, _10308_);
  not (_10559_, _10323_);
  or (_10560_, _10330_, _10559_);
  and (_10561_, _10344_, _10337_);
  and (_10562_, _10354_, _05855_);
  nor (_10563_, _10562_, _10349_);
  or (_10564_, _10563_, _10350_);
  nand (_10565_, _10564_, _10561_);
  nor (_10566_, _10342_, _10335_);
  or (_10567_, _10566_, _10336_);
  and (_10568_, _10567_, _10565_);
  nor (_10569_, _10568_, _10560_);
  nor (_10570_, _10328_, _10321_);
  nor (_10571_, _10570_, _10322_);
  nor (_10572_, _10571_, _10569_);
  nor (_10573_, _10572_, _10316_);
  or (_10574_, _10573_, _10313_);
  and (_10575_, _10574_, _10558_);
  nor (_10576_, _10574_, _10558_);
  or (_10577_, _10576_, _10575_);
  and (_10578_, _10577_, _10557_);
  or (_10579_, _10578_, _10556_);
  and (_10580_, _06284_, _05790_);
  not (_10581_, _10580_);
  and (_10582_, _10581_, _10579_);
  and (_10583_, _09217_, \oc8051_golden_model_1.PSW [7]);
  nor (_10584_, _10583_, _08838_);
  and (_10585_, _10583_, _08838_);
  nor (_10586_, _10585_, _10584_);
  and (_10587_, _10586_, \oc8051_golden_model_1.ACC [7]);
  nor (_10588_, _10586_, \oc8051_golden_model_1.ACC [7]);
  nor (_10589_, _10588_, _10587_);
  and (_10590_, _09216_, \oc8051_golden_model_1.PSW [7]);
  nor (_10591_, _10590_, _09207_);
  nor (_10592_, _10591_, _10583_);
  nor (_10593_, _10592_, _09883_);
  and (_10594_, _09215_, \oc8051_golden_model_1.PSW [7]);
  nor (_10595_, _10594_, _09208_);
  nor (_10596_, _10595_, _10590_);
  nor (_10597_, _10596_, _09930_);
  and (_10598_, _10596_, _09930_);
  nor (_10599_, _10598_, _10597_);
  not (_10600_, _10599_);
  and (_10601_, _09214_, \oc8051_golden_model_1.PSW [7]);
  nor (_10602_, _10601_, _09209_);
  nor (_10603_, _10602_, _10594_);
  nor (_10604_, _10603_, _09902_);
  and (_10605_, _10603_, _09902_);
  or (_10606_, _10605_, _10604_);
  or (_10607_, _10606_, _10600_);
  and (_10608_, _09213_, \oc8051_golden_model_1.PSW [7]);
  nor (_10609_, _10608_, _09210_);
  nor (_10610_, _10609_, _10601_);
  nor (_10611_, _10610_, _10028_);
  and (_10612_, _10610_, _10028_);
  nor (_10613_, _10612_, _10611_);
  and (_10614_, _09212_, \oc8051_golden_model_1.PSW [7]);
  nor (_10615_, _10614_, _09211_);
  nor (_10616_, _10615_, _10608_);
  nor (_10617_, _10616_, _09981_);
  and (_10618_, _10616_, _09981_);
  nor (_10619_, _10618_, _10617_);
  and (_10620_, _10619_, _10613_);
  and (_10621_, _09160_, \oc8051_golden_model_1.PSW [7]);
  nor (_10622_, _10621_, _09115_);
  nor (_10623_, _10622_, _10614_);
  nor (_10624_, _10623_, _05887_);
  and (_10625_, _10623_, _05887_);
  nor (_10626_, _09160_, \oc8051_golden_model_1.PSW [7]);
  nor (_10627_, _10626_, _10621_);
  and (_10628_, _10627_, _05855_);
  nor (_10629_, _10628_, _10625_);
  or (_10630_, _10629_, _10624_);
  nand (_10631_, _10630_, _10620_);
  nor (_10632_, _10617_, _10611_);
  or (_10633_, _10632_, _10612_);
  and (_10634_, _10633_, _10631_);
  nor (_10635_, _10634_, _10607_);
  nor (_10636_, _10604_, _10597_);
  nor (_10637_, _10636_, _10598_);
  nor (_10638_, _10637_, _10635_);
  and (_10639_, _10592_, _09883_);
  nor (_10640_, _10593_, _10639_);
  not (_10641_, _10640_);
  nor (_10642_, _10641_, _10638_);
  or (_10643_, _10642_, _10593_);
  nor (_10644_, _10643_, _10589_);
  and (_10645_, _10643_, _10589_);
  or (_10646_, _10645_, _10644_);
  nor (_10647_, _10646_, _10581_);
  or (_10648_, _10647_, _10582_);
  and (_10649_, _10648_, _06710_);
  nor (_10650_, _10646_, _06710_);
  or (_10651_, _10650_, _10649_);
  or (_10652_, _10651_, _06260_);
  and (_10653_, _10652_, _10455_);
  and (_10654_, _08586_, _06228_);
  and (_10655_, _10654_, _07839_);
  and (_10656_, _10654_, _07828_);
  and (_10657_, _10656_, _07482_);
  nor (_10658_, _10657_, _06039_);
  nor (_10659_, _10658_, _10655_);
  nor (_10660_, _10659_, _08430_);
  and (_10661_, _10659_, _08430_);
  nor (_10662_, _10661_, _10660_);
  nor (_10663_, _10656_, _07482_);
  nor (_10664_, _10663_, _10657_);
  nor (_10665_, _10664_, _09883_);
  and (_10666_, _10654_, _07775_);
  nor (_10667_, _10666_, _07805_);
  nor (_10668_, _10667_, _10656_);
  and (_10669_, _10668_, _09930_);
  nor (_10670_, _10668_, _09930_);
  nor (_10671_, _10654_, _07775_);
  nor (_10672_, _10671_, _10666_);
  nor (_10673_, _10672_, _09902_);
  nor (_10674_, _10673_, _10670_);
  nor (_10675_, _10674_, _10669_);
  nor (_10676_, _10670_, _10669_);
  not (_10677_, _10676_);
  and (_10678_, _10672_, _09902_);
  or (_10679_, _10678_, _10673_);
  or (_10680_, _10679_, _10677_);
  nor (_10681_, _08586_, _06228_);
  nor (_10682_, _10681_, _10654_);
  and (_10683_, _10682_, _10028_);
  nor (_10684_, _10682_, _10028_);
  nor (_10685_, _10684_, _10683_);
  and (_10686_, _07834_, \oc8051_golden_model_1.PSW [7]);
  nor (_10687_, _10686_, _06626_);
  nor (_10688_, _10687_, _08586_);
  and (_10689_, _10688_, _09981_);
  nor (_10690_, _10688_, _09981_);
  nor (_10691_, _10690_, _10689_);
  and (_10692_, _10691_, _10685_);
  not (_10693_, \oc8051_golden_model_1.PSW [7]);
  nor (_10694_, _06107_, _10693_);
  nor (_10695_, _10694_, _06913_);
  nor (_10696_, _10695_, _10686_);
  nor (_10697_, _10696_, _05887_);
  and (_10699_, _10696_, _05887_);
  and (_10700_, _06107_, _10693_);
  nor (_10701_, _10700_, _10694_);
  and (_10702_, _10701_, _05855_);
  nor (_10703_, _10702_, _10699_);
  or (_10704_, _10703_, _10697_);
  nand (_10705_, _10704_, _10692_);
  and (_10706_, _10690_, _10685_);
  nor (_10707_, _10706_, _10684_);
  and (_10708_, _10707_, _10705_);
  nor (_10710_, _10708_, _10680_);
  nor (_10711_, _10710_, _10675_);
  and (_10712_, _10664_, _09883_);
  nor (_10713_, _10665_, _10712_);
  not (_10714_, _10713_);
  nor (_10715_, _10714_, _10711_);
  or (_10716_, _10715_, _10665_);
  nor (_10717_, _10716_, _10662_);
  and (_10718_, _10716_, _10662_);
  or (_10719_, _10718_, _10717_);
  nor (_10721_, _10719_, _10388_);
  or (_10722_, _10721_, _10653_);
  and (_10723_, _10722_, _05805_);
  and (_10724_, _06039_, _05870_);
  or (_10725_, _10724_, _10723_);
  and (_10726_, _10725_, _06140_);
  and (_10727_, _08587_, _08409_);
  or (_10728_, _10727_, _10460_);
  and (_10729_, _10728_, _06139_);
  or (_10730_, _10729_, _09842_);
  or (_10732_, _10730_, _10726_);
  and (_10733_, _10732_, _10386_);
  or (_10734_, _10733_, _06116_);
  and (_10735_, _08535_, _07809_);
  or (_10736_, _10383_, _06117_);
  or (_10737_, _10736_, _10735_);
  and (_10738_, _10737_, _06114_);
  and (_10739_, _10738_, _10734_);
  and (_10740_, _08782_, _07809_);
  or (_10741_, _10740_, _10383_);
  and (_10743_, _10741_, _05787_);
  or (_10744_, _10743_, _09855_);
  or (_10745_, _10744_, _10739_);
  or (_10746_, _09873_, _09861_);
  and (_10747_, _10746_, _10745_);
  or (_10748_, _10747_, _05801_);
  and (_10749_, _10748_, _10382_);
  or (_10750_, _10749_, _06110_);
  and (_10751_, _06294_, _06109_);
  not (_10752_, _10751_);
  and (_10754_, _08607_, _07809_);
  or (_10755_, _10754_, _10383_);
  or (_10756_, _10755_, _06111_);
  and (_10757_, _10756_, _10752_);
  and (_10758_, _10757_, _10750_);
  and (_10759_, _10751_, _06039_);
  or (_10760_, _10759_, _06558_);
  or (_10761_, _10760_, _10758_);
  not (_10762_, _06558_);
  and (_10763_, _09194_, _08430_);
  and (_10765_, _07923_, \oc8051_golden_model_1.ACC [7]);
  nor (_10766_, _10765_, _10763_);
  nor (_10767_, _10766_, _10762_);
  nor (_10768_, _06129_, _05833_);
  nor (_10769_, _10768_, _10767_);
  and (_10770_, _10769_, _10761_);
  and (_10771_, _10768_, _10766_);
  and (_10772_, _06119_, _06399_);
  or (_10773_, _10772_, _10771_);
  or (_10774_, _10773_, _10770_);
  and (_10775_, _06115_, _06399_);
  not (_10776_, _10775_);
  nand (_10777_, _10776_, _10766_);
  nor (_10778_, _07365_, _05833_);
  nand (_10779_, _10778_, _10777_);
  and (_10780_, _10779_, _10774_);
  and (_10781_, _08838_, _08430_);
  and (_10782_, _08535_, \oc8051_golden_model_1.ACC [7]);
  nor (_10783_, _10782_, _10781_);
  and (_10784_, _10775_, _10783_);
  or (_10785_, _10784_, _06400_);
  or (_10786_, _10785_, _10780_);
  and (_10787_, _06294_, _06399_);
  not (_10788_, _10787_);
  or (_10789_, _08810_, _06401_);
  and (_10790_, _10789_, _10788_);
  and (_10791_, _10790_, _10786_);
  nor (_10792_, _06039_, \oc8051_golden_model_1.ACC [7]);
  and (_10793_, _06039_, \oc8051_golden_model_1.ACC [7]);
  nor (_10794_, _10793_, _10792_);
  and (_10795_, _10787_, _10794_);
  or (_10796_, _10795_, _06297_);
  or (_10797_, _10796_, _10791_);
  and (_10798_, _08802_, _07809_);
  or (_10799_, _10798_, _10383_);
  or (_10800_, _10799_, _07127_);
  and (_10801_, _10800_, _10797_);
  or (_10802_, _10801_, _06402_);
  or (_10803_, _10383_, _07125_);
  nor (_10804_, _06129_, _05847_);
  and (_10805_, _06125_, _06408_);
  or (_10806_, _10805_, _10804_);
  and (_10807_, _06119_, _06408_);
  nor (_10808_, _10807_, _10806_);
  and (_10809_, _10808_, _10803_);
  and (_10810_, _10809_, _10802_);
  and (_10811_, _06115_, _06408_);
  not (_10812_, _10808_);
  and (_10813_, _10812_, _10765_);
  or (_10814_, _10813_, _10811_);
  or (_10815_, _10814_, _10810_);
  not (_10816_, _10811_);
  or (_10817_, _10816_, _10782_);
  and (_10818_, _10817_, _06410_);
  and (_10819_, _10818_, _10815_);
  and (_10820_, _06294_, _06408_);
  nor (_10821_, _10820_, _06409_);
  not (_10822_, _10821_);
  or (_10823_, _10820_, _08808_);
  and (_10824_, _10823_, _10822_);
  or (_10825_, _10824_, _10819_);
  not (_10826_, _10820_);
  or (_10827_, _10826_, _10793_);
  and (_10828_, _10827_, _07132_);
  and (_10829_, _10828_, _10825_);
  nand (_10830_, _10755_, _06306_);
  nor (_10831_, _10830_, _08809_);
  or (_10832_, _10831_, _06524_);
  or (_10833_, _10832_, _10829_);
  not (_10834_, _06555_);
  and (_10835_, _06119_, _05840_);
  nor (_10836_, _10835_, _06975_);
  and (_10837_, _10836_, _10834_);
  nand (_10838_, _10763_, _06524_);
  and (_10839_, _10838_, _10837_);
  and (_10840_, _10839_, _10833_);
  and (_10841_, _06115_, _05840_);
  nor (_10842_, _10837_, _10763_);
  or (_10843_, _10842_, _10841_);
  or (_10844_, _10843_, _10840_);
  nand (_10845_, _10841_, _10781_);
  and (_10846_, _10845_, _06395_);
  and (_10847_, _10846_, _10844_);
  and (_10848_, _06294_, _05840_);
  nor (_10849_, _10848_, _06394_);
  not (_10850_, _10849_);
  not (_10851_, _10848_);
  nand (_10852_, _10851_, _08809_);
  and (_10853_, _10852_, _10850_);
  or (_10854_, _10853_, _10847_);
  nand (_10855_, _10848_, _10792_);
  and (_10856_, _10855_, _08819_);
  and (_10857_, _10856_, _10854_);
  not (_10858_, _10380_);
  and (_10859_, _08801_, _07809_);
  or (_10860_, _10859_, _10383_);
  and (_10861_, _10860_, _06303_);
  or (_10862_, _10861_, _10858_);
  or (_10863_, _10862_, _10857_);
  and (_10864_, _10863_, _10381_);
  and (_10865_, _06115_, _06300_);
  or (_10866_, _10865_, _10864_);
  not (_10867_, _10865_);
  nand (_10868_, _10592_, \oc8051_golden_model_1.ACC [6]);
  and (_10869_, _10596_, \oc8051_golden_model_1.ACC [5]);
  nand (_10870_, _10603_, \oc8051_golden_model_1.ACC [4]);
  and (_10871_, _10610_, \oc8051_golden_model_1.ACC [3]);
  and (_10872_, _10616_, \oc8051_golden_model_1.ACC [2]);
  and (_10873_, _10623_, \oc8051_golden_model_1.ACC [1]);
  nor (_10874_, _10625_, _10624_);
  not (_10875_, _10874_);
  and (_10876_, _10627_, \oc8051_golden_model_1.ACC [0]);
  and (_10877_, _10876_, _10875_);
  nor (_10878_, _10877_, _10873_);
  nor (_10879_, _10878_, _10619_);
  nor (_10880_, _10879_, _10872_);
  nor (_10881_, _10880_, _10613_);
  or (_10882_, _10881_, _10871_);
  nand (_10883_, _10882_, _10606_);
  and (_10884_, _10883_, _10870_);
  nor (_10885_, _10884_, _10599_);
  or (_10886_, _10885_, _10869_);
  nand (_10887_, _10886_, _10641_);
  and (_10888_, _10887_, _10868_);
  nor (_10889_, _10888_, _10589_);
  and (_10890_, _10888_, _10589_);
  nor (_10891_, _10890_, _10889_);
  or (_10892_, _10891_, _10867_);
  and (_10893_, _10892_, _06407_);
  and (_10894_, _10893_, _10866_);
  and (_10895_, _06294_, _06300_);
  nor (_10896_, _10895_, _06406_);
  not (_10897_, _10896_);
  and (_10898_, _10404_, \oc8051_golden_model_1.ACC [6]);
  and (_10899_, _10407_, \oc8051_golden_model_1.ACC [5]);
  nand (_10900_, _10413_, \oc8051_golden_model_1.ACC [4]);
  and (_10901_, _10419_, \oc8051_golden_model_1.ACC [3]);
  and (_10902_, _10424_, \oc8051_golden_model_1.ACC [2]);
  and (_10903_, _10430_, \oc8051_golden_model_1.ACC [1]);
  nor (_10904_, _10432_, _10431_);
  not (_10905_, _10904_);
  and (_10906_, _10434_, \oc8051_golden_model_1.ACC [0]);
  and (_10907_, _10906_, _10905_);
  nor (_10908_, _10907_, _10903_);
  nor (_10909_, _10908_, _10427_);
  nor (_10910_, _10909_, _10902_);
  nor (_10911_, _10910_, _10422_);
  or (_10912_, _10911_, _10901_);
  nand (_10913_, _10912_, _10416_);
  and (_10914_, _10913_, _10900_);
  nor (_10915_, _10914_, _10410_);
  or (_10916_, _10915_, _10899_);
  and (_10917_, _10916_, _10448_);
  nor (_10918_, _10917_, _10898_);
  nor (_10919_, _10918_, _10401_);
  and (_10920_, _10918_, _10401_);
  nor (_10921_, _10920_, _10919_);
  or (_10922_, _10921_, _10895_);
  and (_10923_, _10922_, _10897_);
  or (_10924_, _10923_, _10894_);
  nor (_10925_, _05844_, _05799_);
  not (_10926_, _10925_);
  not (_10927_, _10895_);
  and (_10928_, _10664_, \oc8051_golden_model_1.ACC [6]);
  and (_10929_, _10668_, \oc8051_golden_model_1.ACC [5]);
  nand (_10930_, _10672_, \oc8051_golden_model_1.ACC [4]);
  and (_10931_, _10682_, \oc8051_golden_model_1.ACC [3]);
  and (_10932_, _10688_, \oc8051_golden_model_1.ACC [2]);
  and (_10933_, _10696_, \oc8051_golden_model_1.ACC [1]);
  nor (_10934_, _10699_, _10697_);
  not (_10935_, _10934_);
  and (_10936_, _10701_, \oc8051_golden_model_1.ACC [0]);
  and (_10937_, _10936_, _10935_);
  nor (_10938_, _10937_, _10933_);
  nor (_10939_, _10938_, _10691_);
  nor (_10940_, _10939_, _10932_);
  nor (_10941_, _10940_, _10685_);
  or (_10942_, _10941_, _10931_);
  nand (_10943_, _10942_, _10679_);
  and (_10944_, _10943_, _10930_);
  nor (_10945_, _10944_, _10676_);
  or (_10946_, _10945_, _10929_);
  and (_10947_, _10946_, _10714_);
  nor (_10948_, _10947_, _10928_);
  nor (_10949_, _10948_, _10662_);
  and (_10950_, _10948_, _10662_);
  nor (_10951_, _10950_, _10949_);
  or (_10952_, _10951_, _10927_);
  and (_10953_, _10952_, _10926_);
  and (_10954_, _10953_, _10924_);
  nand (_10955_, _10925_, \oc8051_golden_model_1.ACC [6]);
  and (_10956_, _06273_, _05825_);
  not (_10957_, _10956_);
  and (_10958_, _06288_, _05825_);
  nor (_10959_, _10958_, _06952_);
  and (_10960_, _06122_, _05825_);
  nor (_10961_, _06958_, _10960_);
  and (_10962_, _10961_, _10959_);
  and (_10963_, _10962_, _10957_);
  nand (_10964_, _10963_, _10955_);
  or (_10965_, _10964_, _10954_);
  and (_10966_, _08012_, \oc8051_golden_model_1.ACC [6]);
  or (_10967_, _08012_, \oc8051_golden_model_1.ACC [6]);
  not (_10968_, _10966_);
  and (_10969_, _10968_, _10967_);
  and (_10970_, _08101_, \oc8051_golden_model_1.ACC [5]);
  and (_10971_, _08348_, _09930_);
  and (_10972_, _08336_, \oc8051_golden_model_1.ACC [4]);
  or (_10973_, _08336_, \oc8051_golden_model_1.ACC [4]);
  not (_10974_, _10972_);
  and (_10975_, _10974_, _10973_);
  and (_10976_, _07544_, \oc8051_golden_model_1.ACC [3]);
  and (_10977_, _07474_, _10028_);
  and (_10978_, _07708_, \oc8051_golden_model_1.ACC [2]);
  and (_10979_, _07657_, _09981_);
  nor (_10980_, _10978_, _10979_);
  not (_10981_, _10980_);
  and (_10982_, _07306_, \oc8051_golden_model_1.ACC [1]);
  and (_10983_, _07252_, _05887_);
  nor (_10984_, _10982_, _10983_);
  and (_10985_, _07049_, \oc8051_golden_model_1.ACC [0]);
  and (_10986_, _10985_, _10984_);
  nor (_10987_, _10986_, _10982_);
  nor (_10988_, _10987_, _10981_);
  nor (_10989_, _10988_, _10978_);
  nor (_10990_, _10989_, _10977_);
  or (_10991_, _10990_, _10976_);
  and (_10992_, _10991_, _10975_);
  nor (_10993_, _10992_, _10972_);
  nor (_10994_, _10993_, _10971_);
  or (_10995_, _10994_, _10970_);
  and (_10996_, _10995_, _10969_);
  nor (_10997_, _10996_, _10966_);
  and (_10998_, _10997_, _10766_);
  nor (_10999_, _10997_, _10766_);
  or (_11000_, _10999_, _10998_);
  or (_11001_, _11000_, _10963_);
  and (_11002_, _11001_, _10965_);
  and (_11003_, _06115_, _05825_);
  or (_11004_, _11003_, _11002_);
  and (_11005_, _09207_, \oc8051_golden_model_1.ACC [6]);
  or (_11006_, _09207_, \oc8051_golden_model_1.ACC [6]);
  not (_11007_, _11005_);
  and (_11008_, _11007_, _11006_);
  and (_11009_, _09208_, \oc8051_golden_model_1.ACC [5]);
  and (_11010_, _08931_, _09930_);
  or (_11011_, _11010_, _11009_);
  and (_11012_, _09209_, \oc8051_golden_model_1.ACC [4]);
  not (_11013_, _11012_);
  or (_11014_, _09209_, \oc8051_golden_model_1.ACC [4]);
  and (_11015_, _11013_, _11014_);
  and (_11016_, _09210_, \oc8051_golden_model_1.ACC [3]);
  and (_11017_, _09025_, _10028_);
  and (_11018_, _09211_, \oc8051_golden_model_1.ACC [2]);
  or (_11019_, _09211_, \oc8051_golden_model_1.ACC [2]);
  not (_11020_, _11018_);
  and (_11021_, _11020_, _11019_);
  not (_11022_, _11021_);
  and (_11023_, _09115_, \oc8051_golden_model_1.ACC [1]);
  or (_11024_, _09115_, \oc8051_golden_model_1.ACC [1]);
  not (_11025_, _11023_);
  and (_11026_, _11025_, _11024_);
  and (_11027_, _09160_, \oc8051_golden_model_1.ACC [0]);
  and (_11028_, _11027_, _11026_);
  nor (_11029_, _11028_, _11023_);
  nor (_11030_, _11029_, _11022_);
  nor (_11031_, _11030_, _11018_);
  nor (_11032_, _11031_, _11017_);
  or (_11033_, _11032_, _11016_);
  nand (_11034_, _11033_, _11015_);
  and (_11035_, _11034_, _11013_);
  nor (_11036_, _11035_, _11011_);
  or (_11037_, _11036_, _11009_);
  and (_11038_, _11037_, _11008_);
  nor (_11039_, _11038_, _11005_);
  and (_11040_, _11039_, _10783_);
  not (_11041_, _11003_);
  nor (_11042_, _11039_, _10783_);
  or (_11043_, _11042_, _11041_);
  or (_11044_, _11043_, _11040_);
  and (_11045_, _11044_, _06171_);
  and (_11046_, _11045_, _11004_);
  or (_11047_, _11046_, _10301_);
  and (_11048_, _11047_, _10265_);
  nor (_11049_, _06203_, _09883_);
  not (_11050_, _11049_);
  and (_11051_, _06203_, _09883_);
  nor (_11052_, _11049_, _11051_);
  nor (_11053_, _06477_, _09930_);
  and (_11054_, _06477_, _09930_);
  nor (_11055_, _06876_, _09902_);
  not (_11056_, _11055_);
  and (_11057_, _06876_, _09902_);
  nor (_11058_, _11055_, _11057_);
  nor (_11059_, _06070_, _10028_);
  and (_11060_, _06070_, _10028_);
  nor (_11061_, _06625_, _09981_);
  and (_11062_, _06625_, _09981_);
  nor (_11063_, _11061_, _11062_);
  nor (_11064_, _06912_, _05887_);
  and (_11065_, _06912_, _05887_);
  nor (_11066_, _11064_, _11065_);
  nor (_11067_, _06107_, _05855_);
  and (_11068_, _11067_, _11066_);
  nor (_11069_, _11068_, _11064_);
  not (_11070_, _11069_);
  and (_11071_, _11070_, _11063_);
  nor (_11072_, _11071_, _11061_);
  nor (_11073_, _11072_, _11060_);
  or (_11074_, _11073_, _11059_);
  nand (_11075_, _11074_, _11058_);
  and (_11076_, _11075_, _11056_);
  nor (_11077_, _11076_, _11054_);
  or (_11078_, _11077_, _11053_);
  nand (_11079_, _11078_, _11052_);
  and (_11080_, _11079_, _11050_);
  nor (_11081_, _11080_, _10794_);
  and (_11082_, _11080_, _10794_);
  or (_11083_, _11082_, _11081_);
  and (_11084_, _11083_, _10264_);
  or (_11085_, _11084_, _10262_);
  or (_11086_, _11085_, _11048_);
  and (_11087_, _11086_, _10263_);
  or (_11088_, _11087_, _06433_);
  and (_11089_, _06294_, _05591_);
  not (_11090_, _11089_);
  or (_11091_, _10487_, _06829_);
  and (_11092_, _11091_, _11090_);
  and (_11093_, _11092_, _11088_);
  and (_11094_, _06302_, _05591_);
  and (_11095_, _10493_, _05855_);
  and (_11096_, _11095_, _10028_);
  and (_11097_, _11096_, _09902_);
  and (_11098_, _11097_, _09930_);
  and (_11099_, _11098_, _09883_);
  nor (_11100_, _11099_, _08430_);
  and (_11101_, _11099_, _08430_);
  or (_11102_, _11101_, _11100_);
  and (_11103_, _11102_, _11089_);
  or (_11104_, _11103_, _11094_);
  or (_11105_, _11104_, _11093_);
  nand (_11106_, _11094_, _10693_);
  and (_11107_, _11106_, _05749_);
  and (_11108_, _11107_, _11105_);
  and (_11109_, _10533_, _05748_);
  or (_11110_, _11109_, _06440_);
  or (_11111_, _11110_, _11108_);
  and (_11112_, _06294_, _05820_);
  not (_11113_, _11112_);
  and (_11114_, _08345_, _07809_);
  or (_11115_, _10383_, _06444_);
  or (_11116_, _11115_, _11114_);
  and (_11117_, _11116_, _11113_);
  and (_11118_, _11117_, _11111_);
  and (_11119_, _05820_, _06302_);
  and (_11120_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  and (_11121_, _11120_, \oc8051_golden_model_1.ACC [2]);
  and (_11122_, _11121_, \oc8051_golden_model_1.ACC [3]);
  and (_11123_, _11122_, \oc8051_golden_model_1.ACC [4]);
  and (_11124_, _11123_, \oc8051_golden_model_1.ACC [5]);
  and (_11125_, _11124_, \oc8051_golden_model_1.ACC [6]);
  nor (_11126_, _11125_, _08430_);
  and (_11127_, _11125_, _08430_);
  or (_11128_, _11127_, _11126_);
  and (_11129_, _11128_, _11112_);
  or (_11130_, _11129_, _11119_);
  or (_11131_, _11130_, _11118_);
  nand (_11132_, _11119_, _05855_);
  and (_11133_, _11132_, _01317_);
  and (_11134_, _11133_, _11131_);
  or (_11135_, _11134_, _10261_);
  and (_40981_, _11135_, _43100_);
  not (_11136_, _06298_);
  not (_11137_, _07856_);
  and (_11138_, _11137_, \oc8051_golden_model_1.PCON [7]);
  and (_11139_, _07923_, _07856_);
  or (_11140_, _11139_, _11138_);
  or (_11141_, _11140_, _06132_);
  and (_11142_, _08548_, _07856_);
  or (_11143_, _11142_, _11138_);
  or (_11144_, _11143_, _06161_);
  and (_11145_, _07856_, \oc8051_golden_model_1.ACC [7]);
  or (_11146_, _11145_, _11138_);
  and (_11147_, _11146_, _07056_);
  and (_11148_, _07057_, \oc8051_golden_model_1.PCON [7]);
  or (_11149_, _11148_, _06160_);
  or (_11150_, _11149_, _11147_);
  and (_11151_, _11150_, _07075_);
  and (_11152_, _11151_, _11144_);
  and (_11153_, _11140_, _06217_);
  or (_11154_, _11153_, _11152_);
  and (_11155_, _11154_, _06229_);
  and (_11156_, _11146_, _06220_);
  or (_11157_, _11156_, _09842_);
  or (_11158_, _11157_, _11155_);
  and (_11159_, _11158_, _11141_);
  or (_11160_, _11159_, _06116_);
  and (_11161_, _08535_, _07856_);
  or (_11162_, _11138_, _06117_);
  or (_11163_, _11162_, _11161_);
  and (_11164_, _11163_, _06114_);
  and (_11165_, _11164_, _11160_);
  and (_11166_, _08782_, _07856_);
  or (_11167_, _11166_, _11138_);
  and (_11168_, _11167_, _05787_);
  or (_11169_, _11168_, _11165_);
  or (_11170_, _11169_, _11136_);
  and (_11171_, _08802_, _07856_);
  or (_11172_, _11138_, _07127_);
  or (_11173_, _11172_, _11171_);
  and (_11174_, _08607_, _07856_);
  or (_11175_, _11174_, _11138_);
  or (_11176_, _11175_, _06111_);
  and (_11177_, _11176_, _07125_);
  and (_11178_, _11177_, _11173_);
  and (_11179_, _11178_, _11170_);
  and (_11180_, _08810_, _07856_);
  or (_11181_, _11180_, _11138_);
  and (_11182_, _11181_, _06402_);
  or (_11183_, _11182_, _11179_);
  and (_11184_, _11183_, _07132_);
  or (_11185_, _11138_, _07926_);
  and (_11186_, _11175_, _06306_);
  and (_11187_, _11186_, _11185_);
  or (_11188_, _11187_, _11184_);
  and (_11189_, _11188_, _07130_);
  and (_11190_, _11146_, _06411_);
  and (_11191_, _11190_, _11185_);
  or (_11192_, _11191_, _06303_);
  or (_11193_, _11192_, _11189_);
  and (_11194_, _08801_, _07856_);
  or (_11195_, _11138_, _08819_);
  or (_11196_, _11195_, _11194_);
  and (_11197_, _11196_, _08824_);
  and (_11198_, _11197_, _11193_);
  nor (_11199_, _08809_, _11137_);
  or (_11200_, _11199_, _11138_);
  and (_11201_, _11200_, _06396_);
  or (_11202_, _11201_, _06433_);
  or (_11203_, _11202_, _11198_);
  or (_11204_, _11143_, _06829_);
  and (_11205_, _11204_, _06444_);
  and (_11206_, _11205_, _11203_);
  and (_11207_, _08345_, _07856_);
  or (_11208_, _11207_, _11138_);
  and (_11209_, _11208_, _06440_);
  or (_11210_, _11209_, _01321_);
  or (_11211_, _11210_, _11206_);
  or (_11212_, _01317_, \oc8051_golden_model_1.PCON [7]);
  and (_11213_, _11212_, _43100_);
  and (_40982_, _11213_, _11211_);
  not (_11214_, _07812_);
  and (_11215_, _11214_, \oc8051_golden_model_1.TMOD [7]);
  and (_11216_, _07923_, _07812_);
  or (_11217_, _11216_, _11215_);
  or (_11218_, _11217_, _06132_);
  and (_11219_, _08548_, _07812_);
  or (_11220_, _11219_, _11215_);
  or (_11221_, _11220_, _06161_);
  and (_11222_, _07812_, \oc8051_golden_model_1.ACC [7]);
  or (_11223_, _11222_, _11215_);
  and (_11224_, _11223_, _07056_);
  and (_11225_, _07057_, \oc8051_golden_model_1.TMOD [7]);
  or (_11226_, _11225_, _06160_);
  or (_11227_, _11226_, _11224_);
  and (_11228_, _11227_, _07075_);
  and (_11229_, _11228_, _11221_);
  and (_11230_, _11217_, _06217_);
  or (_11231_, _11230_, _11229_);
  and (_11232_, _11231_, _06229_);
  and (_11233_, _11223_, _06220_);
  or (_11234_, _11233_, _09842_);
  or (_11235_, _11234_, _11232_);
  and (_11236_, _11235_, _11218_);
  or (_11237_, _11236_, _06116_);
  and (_11238_, _08535_, _07812_);
  or (_11239_, _11215_, _06117_);
  or (_11240_, _11239_, _11238_);
  and (_11241_, _11240_, _06114_);
  and (_11242_, _11241_, _11237_);
  and (_11243_, _08782_, _07812_);
  or (_11244_, _11243_, _11215_);
  and (_11245_, _11244_, _05787_);
  or (_11246_, _11245_, _11242_);
  or (_11247_, _11246_, _11136_);
  and (_11248_, _08802_, _07812_);
  or (_11249_, _11215_, _07127_);
  or (_11250_, _11249_, _11248_);
  and (_11251_, _08607_, _07812_);
  or (_11252_, _11251_, _11215_);
  or (_11253_, _11252_, _06111_);
  and (_11254_, _11253_, _07125_);
  and (_11255_, _11254_, _11250_);
  and (_11256_, _11255_, _11247_);
  and (_11257_, _08810_, _07812_);
  or (_11258_, _11257_, _11215_);
  and (_11259_, _11258_, _06402_);
  or (_11260_, _11259_, _11256_);
  and (_11261_, _11260_, _07132_);
  or (_11262_, _11215_, _07926_);
  and (_11263_, _11252_, _06306_);
  and (_11264_, _11263_, _11262_);
  or (_11265_, _11264_, _11261_);
  and (_11266_, _11265_, _07130_);
  and (_11267_, _11223_, _06411_);
  and (_11268_, _11267_, _11262_);
  or (_11269_, _11268_, _06303_);
  or (_11270_, _11269_, _11266_);
  and (_11271_, _08801_, _07812_);
  or (_11272_, _11215_, _08819_);
  or (_11273_, _11272_, _11271_);
  and (_11274_, _11273_, _08824_);
  and (_11275_, _11274_, _11270_);
  nor (_11276_, _08809_, _11214_);
  or (_11277_, _11276_, _11215_);
  and (_11278_, _11277_, _06396_);
  or (_11279_, _11278_, _06433_);
  or (_11280_, _11279_, _11275_);
  or (_11281_, _11220_, _06829_);
  and (_11282_, _11281_, _06444_);
  and (_11283_, _11282_, _11280_);
  and (_11284_, _08345_, _07812_);
  or (_11285_, _11284_, _11215_);
  and (_11286_, _11285_, _06440_);
  or (_11287_, _11286_, _01321_);
  or (_11288_, _11287_, _11283_);
  or (_11289_, _01317_, \oc8051_golden_model_1.TMOD [7]);
  and (_11290_, _11289_, _43100_);
  and (_40983_, _11290_, _11288_);
  not (_11291_, \oc8051_golden_model_1.DPL [7]);
  nor (_11292_, _07849_, _11291_);
  and (_11293_, _07923_, _07849_);
  or (_11294_, _11293_, _11292_);
  or (_11295_, _11294_, _06132_);
  not (_11296_, _06293_);
  and (_11297_, _08548_, _07849_);
  or (_11298_, _11297_, _11292_);
  or (_11299_, _11298_, _06161_);
  and (_11300_, _07849_, \oc8051_golden_model_1.ACC [7]);
  or (_11301_, _11300_, _11292_);
  and (_11302_, _11301_, _07056_);
  nor (_11303_, _07056_, _11291_);
  or (_11304_, _11303_, _06160_);
  or (_11305_, _11304_, _11302_);
  and (_11306_, _11305_, _07075_);
  and (_11307_, _11306_, _11299_);
  and (_11308_, _11294_, _06217_);
  or (_11309_, _11308_, _06220_);
  or (_11310_, _11309_, _11307_);
  nor (_11311_, _05799_, _05774_);
  not (_11312_, _11311_);
  or (_11313_, _11301_, _06229_);
  and (_11314_, _11313_, _11312_);
  and (_11315_, _11314_, _11310_);
  and (_11316_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_11317_, _11316_, \oc8051_golden_model_1.DPL [2]);
  and (_11318_, _11317_, \oc8051_golden_model_1.DPL [3]);
  and (_11319_, _11318_, \oc8051_golden_model_1.DPL [4]);
  and (_11320_, _11319_, \oc8051_golden_model_1.DPL [5]);
  and (_11321_, _11320_, \oc8051_golden_model_1.DPL [6]);
  nor (_11322_, _11321_, \oc8051_golden_model_1.DPL [7]);
  and (_11323_, _11321_, \oc8051_golden_model_1.DPL [7]);
  nor (_11324_, _11323_, _11322_);
  and (_11325_, _11324_, _11311_);
  or (_11326_, _11325_, _11315_);
  and (_11327_, _11326_, _11296_);
  nor (_11328_, _08395_, _11296_);
  or (_11329_, _11328_, _09842_);
  or (_11330_, _11329_, _11327_);
  and (_11331_, _11330_, _11295_);
  or (_11332_, _11331_, _06116_);
  and (_11333_, _08535_, _07849_);
  or (_11334_, _11292_, _06117_);
  or (_11335_, _11334_, _11333_);
  and (_11336_, _11335_, _06114_);
  and (_11337_, _11336_, _11332_);
  and (_11338_, _08782_, _07849_);
  or (_11339_, _11338_, _11292_);
  and (_11340_, _11339_, _05787_);
  or (_11341_, _11340_, _11337_);
  or (_11342_, _11341_, _11136_);
  and (_11343_, _08802_, _07849_);
  or (_11344_, _11292_, _07127_);
  or (_11345_, _11344_, _11343_);
  and (_11346_, _08607_, _07849_);
  or (_11347_, _11346_, _11292_);
  or (_11348_, _11347_, _06111_);
  and (_11349_, _11348_, _07125_);
  and (_11350_, _11349_, _11345_);
  and (_11351_, _11350_, _11342_);
  and (_11352_, _08810_, _07849_);
  or (_11353_, _11352_, _11292_);
  and (_11354_, _11353_, _06402_);
  or (_11355_, _11354_, _11351_);
  and (_11356_, _11355_, _07132_);
  or (_11357_, _11292_, _07926_);
  and (_11358_, _11347_, _06306_);
  and (_11359_, _11358_, _11357_);
  or (_11360_, _11359_, _11356_);
  and (_11361_, _11360_, _07130_);
  and (_11362_, _11301_, _06411_);
  and (_11363_, _11362_, _11357_);
  or (_11364_, _11363_, _06303_);
  or (_11365_, _11364_, _11361_);
  and (_11366_, _08801_, _07849_);
  or (_11367_, _11292_, _08819_);
  or (_11368_, _11367_, _11366_);
  and (_11369_, _11368_, _08824_);
  and (_11370_, _11369_, _11365_);
  not (_11371_, _07849_);
  nor (_11372_, _08809_, _11371_);
  or (_11373_, _11372_, _11292_);
  and (_11374_, _11373_, _06396_);
  or (_11375_, _11374_, _06433_);
  or (_11376_, _11375_, _11370_);
  or (_11377_, _11298_, _06829_);
  and (_11378_, _11377_, _06444_);
  and (_11379_, _11378_, _11376_);
  and (_11380_, _08345_, _07849_);
  or (_11381_, _11380_, _11292_);
  and (_11382_, _11381_, _06440_);
  or (_11383_, _11382_, _01321_);
  or (_11384_, _11383_, _11379_);
  or (_11385_, _01317_, \oc8051_golden_model_1.DPL [7]);
  and (_11386_, _11385_, _43100_);
  and (_40985_, _11386_, _11384_);
  not (_11387_, \oc8051_golden_model_1.DPH [7]);
  nand (_11388_, _06625_, _06070_);
  nor (_11389_, _07835_, _11388_);
  and (_11390_, _11389_, _07787_);
  nor (_11391_, _11390_, _11387_);
  and (_11392_, _07923_, _07852_);
  or (_11393_, _11392_, _11391_);
  or (_11394_, _11393_, _06132_);
  and (_11395_, _08548_, _07852_);
  or (_11396_, _11395_, _11391_);
  or (_11397_, _11396_, _06161_);
  and (_11398_, _11390_, \oc8051_golden_model_1.ACC [7]);
  or (_11399_, _11398_, _11391_);
  and (_11400_, _11399_, _07056_);
  nor (_11401_, _07056_, _11387_);
  or (_11402_, _11401_, _06160_);
  or (_11403_, _11402_, _11400_);
  and (_11404_, _11403_, _07075_);
  and (_11405_, _11404_, _11397_);
  and (_11406_, _11393_, _06217_);
  or (_11407_, _11406_, _06220_);
  or (_11408_, _11407_, _11405_);
  or (_11409_, _11399_, _06229_);
  and (_11410_, _11409_, _11312_);
  and (_11411_, _11410_, _11408_);
  and (_11412_, _11323_, \oc8051_golden_model_1.DPH [0]);
  and (_11413_, _11412_, \oc8051_golden_model_1.DPH [1]);
  and (_11414_, _11413_, \oc8051_golden_model_1.DPH [2]);
  and (_11415_, _11414_, \oc8051_golden_model_1.DPH [3]);
  and (_11416_, _11415_, \oc8051_golden_model_1.DPH [4]);
  and (_11417_, _11416_, \oc8051_golden_model_1.DPH [5]);
  and (_11418_, _11417_, \oc8051_golden_model_1.DPH [6]);
  nand (_11419_, _11418_, \oc8051_golden_model_1.DPH [7]);
  or (_11420_, _11418_, \oc8051_golden_model_1.DPH [7]);
  and (_11421_, _11420_, _11311_);
  and (_11422_, _11421_, _11419_);
  or (_11423_, _11422_, _11411_);
  and (_11424_, _11423_, _11296_);
  and (_11425_, _06293_, _06039_);
  or (_11426_, _11425_, _09842_);
  or (_11427_, _11426_, _11424_);
  and (_11428_, _11427_, _11394_);
  or (_11429_, _11428_, _06116_);
  or (_11430_, _11391_, _06117_);
  and (_11431_, _08535_, _11390_);
  or (_11432_, _11431_, _11430_);
  and (_11433_, _11432_, _06114_);
  and (_11434_, _11433_, _11429_);
  and (_11435_, _08782_, _11390_);
  or (_11436_, _11435_, _11391_);
  and (_11437_, _11436_, _05787_);
  or (_11438_, _11437_, _11434_);
  or (_11439_, _11438_, _11136_);
  and (_11440_, _08802_, _07852_);
  or (_11441_, _11391_, _07127_);
  or (_11442_, _11441_, _11440_);
  and (_11443_, _08607_, _11390_);
  or (_11444_, _11443_, _11391_);
  or (_11445_, _11444_, _06111_);
  and (_11446_, _11445_, _07125_);
  and (_11447_, _11446_, _11442_);
  and (_11448_, _11447_, _11439_);
  and (_11449_, _08810_, _07852_);
  or (_11450_, _11449_, _11391_);
  and (_11451_, _11450_, _06402_);
  or (_11452_, _11451_, _11448_);
  and (_11453_, _11452_, _07132_);
  or (_11454_, _11391_, _07926_);
  and (_11455_, _11444_, _06306_);
  and (_11456_, _11455_, _11454_);
  or (_11457_, _11456_, _11453_);
  and (_11458_, _11457_, _07130_);
  and (_11459_, _11399_, _06411_);
  and (_11460_, _11459_, _11454_);
  or (_11461_, _11460_, _06303_);
  or (_11462_, _11461_, _11458_);
  and (_11463_, _08801_, _07852_);
  or (_11464_, _11391_, _08819_);
  or (_11465_, _11464_, _11463_);
  and (_11466_, _11465_, _08824_);
  and (_11467_, _11466_, _11462_);
  not (_11468_, _07852_);
  nor (_11469_, _08809_, _11468_);
  or (_11470_, _11469_, _11391_);
  and (_11471_, _11470_, _06396_);
  or (_11472_, _11471_, _06433_);
  or (_11473_, _11472_, _11467_);
  or (_11474_, _11396_, _06829_);
  and (_11475_, _11474_, _06444_);
  and (_11476_, _11475_, _11473_);
  and (_11477_, _08345_, _07852_);
  or (_11478_, _11477_, _11391_);
  and (_11479_, _11478_, _06440_);
  or (_11480_, _11479_, _01321_);
  or (_11481_, _11480_, _11476_);
  or (_11482_, _01317_, \oc8051_golden_model_1.DPH [7]);
  and (_11483_, _11482_, _43100_);
  and (_40986_, _11483_, _11481_);
  not (_11484_, _07837_);
  and (_11485_, _11484_, \oc8051_golden_model_1.TL1 [7]);
  and (_11486_, _07923_, _07837_);
  or (_11487_, _11486_, _11485_);
  or (_11488_, _11487_, _06132_);
  and (_11489_, _08548_, _07837_);
  or (_11490_, _11489_, _11485_);
  or (_11491_, _11490_, _06161_);
  and (_11492_, _07837_, \oc8051_golden_model_1.ACC [7]);
  or (_11493_, _11492_, _11485_);
  and (_11494_, _11493_, _07056_);
  and (_11495_, _07057_, \oc8051_golden_model_1.TL1 [7]);
  or (_11496_, _11495_, _06160_);
  or (_11497_, _11496_, _11494_);
  and (_11498_, _11497_, _07075_);
  and (_11499_, _11498_, _11491_);
  and (_11500_, _11487_, _06217_);
  or (_11501_, _11500_, _11499_);
  and (_11502_, _11501_, _06229_);
  and (_11503_, _11493_, _06220_);
  or (_11504_, _11503_, _09842_);
  or (_11505_, _11504_, _11502_);
  and (_11506_, _11505_, _11488_);
  or (_11507_, _11506_, _06116_);
  and (_11508_, _08535_, _07837_);
  or (_11509_, _11485_, _06117_);
  or (_11510_, _11509_, _11508_);
  and (_11511_, _11510_, _06114_);
  and (_11512_, _11511_, _11507_);
  and (_11513_, _08782_, _07837_);
  or (_11514_, _11513_, _11485_);
  and (_11515_, _11514_, _05787_);
  or (_11516_, _11515_, _11512_);
  or (_11517_, _11516_, _11136_);
  and (_11518_, _08802_, _07837_);
  or (_11519_, _11485_, _07127_);
  or (_11520_, _11519_, _11518_);
  and (_11521_, _08607_, _07837_);
  or (_11522_, _11521_, _11485_);
  or (_11523_, _11522_, _06111_);
  and (_11524_, _11523_, _07125_);
  and (_11525_, _11524_, _11520_);
  and (_11526_, _11525_, _11517_);
  and (_11527_, _08810_, _07837_);
  or (_11528_, _11527_, _11485_);
  and (_11529_, _11528_, _06402_);
  or (_11530_, _11529_, _11526_);
  and (_11531_, _11530_, _07132_);
  or (_11532_, _11485_, _07926_);
  and (_11533_, _11522_, _06306_);
  and (_11534_, _11533_, _11532_);
  or (_11535_, _11534_, _11531_);
  and (_11536_, _11535_, _07130_);
  and (_11537_, _11493_, _06411_);
  and (_11538_, _11537_, _11532_);
  or (_11539_, _11538_, _06303_);
  or (_11540_, _11539_, _11536_);
  and (_11541_, _08801_, _07837_);
  or (_11542_, _11485_, _08819_);
  or (_11543_, _11542_, _11541_);
  and (_11544_, _11543_, _08824_);
  and (_11545_, _11544_, _11540_);
  nor (_11546_, _08809_, _11484_);
  or (_11547_, _11546_, _11485_);
  and (_11548_, _11547_, _06396_);
  or (_11549_, _11548_, _06433_);
  or (_11550_, _11549_, _11545_);
  or (_11551_, _11490_, _06829_);
  and (_11552_, _11551_, _06444_);
  and (_11553_, _11552_, _11550_);
  and (_11554_, _08345_, _07837_);
  or (_11555_, _11554_, _11485_);
  and (_11556_, _11555_, _06440_);
  or (_11557_, _11556_, _01321_);
  or (_11558_, _11557_, _11553_);
  or (_11559_, _01317_, \oc8051_golden_model_1.TL1 [7]);
  and (_11560_, _11559_, _43100_);
  and (_40987_, _11560_, _11558_);
  not (_11561_, _07803_);
  and (_11562_, _11561_, \oc8051_golden_model_1.TL0 [7]);
  and (_11563_, _07923_, _07803_);
  or (_11564_, _11563_, _11562_);
  or (_11565_, _11564_, _06132_);
  and (_11566_, _08548_, _07803_);
  or (_11567_, _11566_, _11562_);
  or (_11568_, _11567_, _06161_);
  and (_11569_, _07803_, \oc8051_golden_model_1.ACC [7]);
  or (_11570_, _11569_, _11562_);
  and (_11571_, _11570_, _07056_);
  and (_11572_, _07057_, \oc8051_golden_model_1.TL0 [7]);
  or (_11573_, _11572_, _06160_);
  or (_11574_, _11573_, _11571_);
  and (_11575_, _11574_, _07075_);
  and (_11576_, _11575_, _11568_);
  and (_11577_, _11564_, _06217_);
  or (_11578_, _11577_, _11576_);
  and (_11579_, _11578_, _06229_);
  and (_11580_, _11570_, _06220_);
  or (_11581_, _11580_, _09842_);
  or (_11582_, _11581_, _11579_);
  and (_11583_, _11582_, _11565_);
  or (_11584_, _11583_, _06116_);
  and (_11585_, _08535_, _07803_);
  or (_11586_, _11562_, _06117_);
  or (_11587_, _11586_, _11585_);
  and (_11588_, _11587_, _06114_);
  and (_11589_, _11588_, _11584_);
  and (_11590_, _08782_, _07803_);
  or (_11591_, _11590_, _11562_);
  and (_11592_, _11591_, _05787_);
  or (_11593_, _11592_, _11589_);
  or (_11594_, _11593_, _11136_);
  and (_11595_, _08802_, _07803_);
  or (_11596_, _11562_, _07127_);
  or (_11597_, _11596_, _11595_);
  and (_11598_, _08607_, _07803_);
  or (_11599_, _11598_, _11562_);
  or (_11600_, _11599_, _06111_);
  and (_11601_, _11600_, _07125_);
  and (_11602_, _11601_, _11597_);
  and (_11603_, _11602_, _11594_);
  and (_11604_, _08810_, _07803_);
  or (_11605_, _11604_, _11562_);
  and (_11606_, _11605_, _06402_);
  or (_11607_, _11606_, _11603_);
  and (_11608_, _11607_, _07132_);
  or (_11609_, _11562_, _07926_);
  and (_11610_, _11599_, _06306_);
  and (_11611_, _11610_, _11609_);
  or (_11612_, _11611_, _11608_);
  and (_11613_, _11612_, _07130_);
  and (_11614_, _11570_, _06411_);
  and (_11615_, _11614_, _11609_);
  or (_11616_, _11615_, _06303_);
  or (_11617_, _11616_, _11613_);
  and (_11618_, _08801_, _07803_);
  or (_11619_, _11562_, _08819_);
  or (_11620_, _11619_, _11618_);
  and (_11621_, _11620_, _08824_);
  and (_11622_, _11621_, _11617_);
  nor (_11623_, _08809_, _11561_);
  or (_11624_, _11623_, _11562_);
  and (_11625_, _11624_, _06396_);
  or (_11626_, _11625_, _06433_);
  or (_11627_, _11626_, _11622_);
  or (_11628_, _11567_, _06829_);
  and (_11629_, _11628_, _06444_);
  and (_11630_, _11629_, _11627_);
  and (_11631_, _08345_, _07803_);
  or (_11632_, _11631_, _11562_);
  and (_11633_, _11632_, _06440_);
  or (_11634_, _11633_, _01321_);
  or (_11635_, _11634_, _11630_);
  or (_11636_, _01317_, \oc8051_golden_model_1.TL0 [7]);
  and (_11637_, _11636_, _43100_);
  and (_40988_, _11637_, _11635_);
  and (_11638_, _01321_, \oc8051_golden_model_1.TCON [7]);
  not (_11639_, _07788_);
  and (_11640_, _11639_, \oc8051_golden_model_1.TCON [7]);
  and (_11641_, _07923_, _07788_);
  or (_11642_, _11641_, _11640_);
  or (_11643_, _11642_, _06132_);
  not (_11644_, _08407_);
  and (_11645_, _11644_, \oc8051_golden_model_1.TCON [7]);
  and (_11646_, _08426_, _08407_);
  or (_11647_, _11646_, _11645_);
  and (_11648_, _11647_, _06152_);
  and (_11649_, _08548_, _07788_);
  or (_11650_, _11649_, _11640_);
  or (_11651_, _11650_, _06161_);
  and (_11652_, _07788_, \oc8051_golden_model_1.ACC [7]);
  or (_11653_, _11652_, _11640_);
  and (_11654_, _11653_, _07056_);
  and (_11655_, _07057_, \oc8051_golden_model_1.TCON [7]);
  or (_11656_, _11655_, _06160_);
  or (_11657_, _11656_, _11654_);
  and (_11658_, _11657_, _06157_);
  and (_11659_, _11658_, _11651_);
  and (_11660_, _08552_, _08407_);
  or (_11661_, _11660_, _11645_);
  and (_11662_, _11661_, _06156_);
  or (_11663_, _11662_, _06217_);
  or (_11664_, _11663_, _11659_);
  or (_11665_, _11642_, _07075_);
  and (_11666_, _11665_, _11664_);
  or (_11667_, _11666_, _06220_);
  or (_11668_, _11653_, _06229_);
  and (_11669_, _11668_, _06153_);
  and (_11670_, _11669_, _11667_);
  or (_11671_, _11670_, _11648_);
  and (_11672_, _11671_, _06146_);
  and (_11673_, _08569_, _08407_);
  or (_11674_, _11673_, _11645_);
  and (_11675_, _11674_, _06145_);
  or (_11676_, _11675_, _11672_);
  and (_11677_, _11676_, _06140_);
  and (_11678_, _08587_, _08407_);
  or (_11679_, _11678_, _11645_);
  and (_11680_, _11679_, _06139_);
  or (_11681_, _11680_, _09842_);
  or (_11682_, _11681_, _11677_);
  and (_11683_, _11682_, _11643_);
  or (_11684_, _11683_, _06116_);
  and (_11685_, _08535_, _07788_);
  or (_11686_, _11640_, _06117_);
  or (_11687_, _11686_, _11685_);
  and (_11688_, _11687_, _06114_);
  and (_11689_, _11688_, _11684_);
  and (_11690_, _08782_, _07788_);
  or (_11691_, _11690_, _11640_);
  and (_11692_, _11691_, _05787_);
  or (_11693_, _11692_, _11136_);
  or (_11694_, _11693_, _11689_);
  and (_11695_, _08802_, _07788_);
  or (_11696_, _11640_, _07127_);
  or (_11697_, _11696_, _11695_);
  and (_11698_, _08607_, _07788_);
  or (_11699_, _11698_, _11640_);
  or (_11700_, _11699_, _06111_);
  and (_11701_, _11700_, _07125_);
  and (_11702_, _11701_, _11697_);
  and (_11703_, _11702_, _11694_);
  and (_11704_, _08810_, _07788_);
  or (_11705_, _11704_, _11640_);
  and (_11706_, _11705_, _06402_);
  or (_11707_, _11706_, _11703_);
  and (_11708_, _11707_, _07132_);
  or (_11709_, _11640_, _07926_);
  and (_11710_, _11699_, _06306_);
  and (_11711_, _11710_, _11709_);
  or (_11712_, _11711_, _11708_);
  and (_11713_, _11712_, _07130_);
  and (_11714_, _11653_, _06411_);
  and (_11715_, _11714_, _11709_);
  or (_11716_, _11715_, _06303_);
  or (_11717_, _11716_, _11713_);
  and (_11718_, _08801_, _07788_);
  or (_11719_, _11640_, _08819_);
  or (_11720_, _11719_, _11718_);
  and (_11721_, _11720_, _08824_);
  and (_11722_, _11721_, _11717_);
  nor (_11723_, _08809_, _11639_);
  or (_11724_, _11723_, _11640_);
  and (_11725_, _11724_, _06396_);
  or (_11726_, _11725_, _06433_);
  or (_11727_, _11726_, _11722_);
  or (_11728_, _11650_, _06829_);
  and (_11729_, _11728_, _05749_);
  and (_11730_, _11729_, _11727_);
  and (_11731_, _11647_, _05748_);
  or (_11732_, _11731_, _06440_);
  or (_11733_, _11732_, _11730_);
  and (_11734_, _08345_, _07788_);
  or (_11735_, _11640_, _06444_);
  or (_11736_, _11735_, _11734_);
  and (_11737_, _11736_, _01317_);
  and (_11738_, _11737_, _11733_);
  or (_11739_, _11738_, _11638_);
  and (_40989_, _11739_, _43100_);
  not (_11740_, _07817_);
  and (_11741_, _11740_, \oc8051_golden_model_1.TH1 [7]);
  and (_11742_, _08548_, _07817_);
  or (_11743_, _11742_, _11741_);
  or (_11744_, _11743_, _06161_);
  and (_11745_, _07817_, \oc8051_golden_model_1.ACC [7]);
  or (_11746_, _11745_, _11741_);
  and (_11747_, _11746_, _07056_);
  and (_11748_, _07057_, \oc8051_golden_model_1.TH1 [7]);
  or (_11749_, _11748_, _06160_);
  or (_11750_, _11749_, _11747_);
  and (_11751_, _11750_, _07075_);
  and (_11752_, _11751_, _11744_);
  and (_11753_, _07923_, _07817_);
  or (_11754_, _11753_, _11741_);
  and (_11755_, _11754_, _06217_);
  or (_11756_, _11755_, _11752_);
  and (_11757_, _11756_, _06229_);
  and (_11758_, _11746_, _06220_);
  or (_11759_, _11758_, _09842_);
  or (_11760_, _11759_, _11757_);
  or (_11761_, _11754_, _06132_);
  and (_11762_, _11761_, _11760_);
  or (_11763_, _11762_, _06116_);
  and (_11764_, _08535_, _07817_);
  or (_11765_, _11741_, _06117_);
  or (_11766_, _11765_, _11764_);
  and (_11767_, _11766_, _06114_);
  and (_11768_, _11767_, _11763_);
  and (_11769_, _08782_, _07817_);
  or (_11770_, _11769_, _11741_);
  and (_11771_, _11770_, _05787_);
  or (_11772_, _11771_, _11768_);
  or (_11773_, _11772_, _11136_);
  and (_11774_, _08802_, _07817_);
  or (_11775_, _11741_, _07127_);
  or (_11776_, _11775_, _11774_);
  and (_11777_, _08607_, _07817_);
  or (_11778_, _11777_, _11741_);
  or (_11779_, _11778_, _06111_);
  and (_11780_, _11779_, _07125_);
  and (_11781_, _11780_, _11776_);
  and (_11782_, _11781_, _11773_);
  and (_11783_, _08810_, _07817_);
  or (_11784_, _11783_, _11741_);
  and (_11785_, _11784_, _06402_);
  or (_11786_, _11785_, _11782_);
  and (_11787_, _11786_, _07132_);
  or (_11788_, _11741_, _07926_);
  and (_11789_, _11778_, _06306_);
  and (_11790_, _11789_, _11788_);
  or (_11791_, _11790_, _11787_);
  and (_11792_, _11791_, _07130_);
  and (_11793_, _11746_, _06411_);
  and (_11794_, _11793_, _11788_);
  or (_11795_, _11794_, _06303_);
  or (_11796_, _11795_, _11792_);
  and (_11797_, _08801_, _07817_);
  or (_11798_, _11741_, _08819_);
  or (_11799_, _11798_, _11797_);
  and (_11800_, _11799_, _08824_);
  and (_11801_, _11800_, _11796_);
  nor (_11802_, _08809_, _11740_);
  or (_11803_, _11802_, _11741_);
  and (_11804_, _11803_, _06396_);
  or (_11805_, _11804_, _06433_);
  or (_11806_, _11805_, _11801_);
  or (_11807_, _11743_, _06829_);
  and (_11808_, _11807_, _06444_);
  and (_11809_, _11808_, _11806_);
  and (_11810_, _08345_, _07817_);
  or (_11811_, _11810_, _11741_);
  and (_11812_, _11811_, _06440_);
  or (_11813_, _11812_, _01321_);
  or (_11814_, _11813_, _11809_);
  or (_11815_, _01317_, \oc8051_golden_model_1.TH1 [7]);
  and (_11816_, _11815_, _43100_);
  and (_40991_, _11816_, _11814_);
  not (_11817_, _07823_);
  and (_11818_, _11817_, \oc8051_golden_model_1.TH0 [7]);
  and (_11819_, _08548_, _07823_);
  or (_11820_, _11819_, _11818_);
  or (_11821_, _11820_, _06161_);
  and (_11822_, _07823_, \oc8051_golden_model_1.ACC [7]);
  or (_11823_, _11822_, _11818_);
  and (_11824_, _11823_, _07056_);
  and (_11825_, _07057_, \oc8051_golden_model_1.TH0 [7]);
  or (_11826_, _11825_, _06160_);
  or (_11827_, _11826_, _11824_);
  and (_11828_, _11827_, _07075_);
  and (_11829_, _11828_, _11821_);
  and (_11830_, _07923_, _07823_);
  or (_11831_, _11830_, _11818_);
  and (_11832_, _11831_, _06217_);
  or (_11833_, _11832_, _11829_);
  and (_11834_, _11833_, _06229_);
  and (_11835_, _11823_, _06220_);
  or (_11836_, _11835_, _09842_);
  or (_11837_, _11836_, _11834_);
  or (_11838_, _11831_, _06132_);
  and (_11839_, _11838_, _11837_);
  or (_11840_, _11839_, _06116_);
  and (_11841_, _08535_, _07823_);
  or (_11842_, _11818_, _06117_);
  or (_11843_, _11842_, _11841_);
  and (_11844_, _11843_, _06114_);
  and (_11845_, _11844_, _11840_);
  and (_11846_, _08782_, _07823_);
  or (_11847_, _11846_, _11818_);
  and (_11848_, _11847_, _05787_);
  or (_11849_, _11848_, _11845_);
  or (_11850_, _11849_, _11136_);
  and (_11851_, _08802_, _07823_);
  or (_11852_, _11818_, _07127_);
  or (_11853_, _11852_, _11851_);
  and (_11854_, _08607_, _07823_);
  or (_11855_, _11854_, _11818_);
  or (_11856_, _11855_, _06111_);
  and (_11857_, _11856_, _07125_);
  and (_11858_, _11857_, _11853_);
  and (_11859_, _11858_, _11850_);
  and (_11860_, _08810_, _07823_);
  or (_11861_, _11860_, _11818_);
  and (_11862_, _11861_, _06402_);
  or (_11863_, _11862_, _11859_);
  and (_11864_, _11863_, _07132_);
  or (_11865_, _11818_, _07926_);
  and (_11866_, _11855_, _06306_);
  and (_11867_, _11866_, _11865_);
  or (_11868_, _11867_, _11864_);
  and (_11869_, _11868_, _07130_);
  and (_11870_, _11823_, _06411_);
  and (_11871_, _11870_, _11865_);
  or (_11872_, _11871_, _06303_);
  or (_11873_, _11872_, _11869_);
  and (_11874_, _08801_, _07823_);
  or (_11875_, _11818_, _08819_);
  or (_11876_, _11875_, _11874_);
  and (_11877_, _11876_, _08824_);
  and (_11878_, _11877_, _11873_);
  nor (_11879_, _08809_, _11817_);
  or (_11880_, _11879_, _11818_);
  and (_11881_, _11880_, _06396_);
  or (_11882_, _11881_, _06433_);
  or (_11883_, _11882_, _11878_);
  or (_11884_, _11820_, _06829_);
  and (_11885_, _11884_, _06444_);
  and (_11886_, _11885_, _11883_);
  and (_11887_, _08345_, _07823_);
  or (_11888_, _11887_, _11818_);
  and (_11889_, _11888_, _06440_);
  or (_11890_, _11889_, _01321_);
  or (_11891_, _11890_, _11886_);
  or (_11892_, _01317_, \oc8051_golden_model_1.TH0 [7]);
  and (_11893_, _11892_, _43100_);
  and (_40992_, _11893_, _11891_);
  and (_11894_, _08433_, _05426_);
  and (_11895_, _11894_, \oc8051_golden_model_1.PC [7]);
  and (_11896_, _11895_, _09231_);
  and (_11897_, _11896_, \oc8051_golden_model_1.PC [10]);
  and (_11898_, _11897_, \oc8051_golden_model_1.PC [11]);
  and (_11899_, _11898_, \oc8051_golden_model_1.PC [12]);
  and (_11900_, _11899_, \oc8051_golden_model_1.PC [13]);
  and (_11901_, _11900_, \oc8051_golden_model_1.PC [14]);
  or (_11902_, _11901_, \oc8051_golden_model_1.PC [15]);
  nand (_11903_, _11901_, \oc8051_golden_model_1.PC [15]);
  and (_11904_, _11903_, _11902_);
  and (_11905_, _11041_, _10963_);
  or (_11906_, _11905_, _11904_);
  and (_11907_, _10867_, _10380_);
  or (_11908_, _11907_, _11904_);
  nor (_11909_, _08441_, _06783_);
  not (_11910_, _11909_);
  nor (_11911_, _10841_, _10835_);
  and (_11912_, _11911_, _11910_);
  or (_11913_, _11912_, _11904_);
  and (_11914_, _10816_, _10808_);
  or (_11915_, _11914_, _11904_);
  nor (_11916_, _10787_, _06400_);
  not (_11917_, _11916_);
  nor (_11918_, _10778_, _10768_);
  and (_11919_, _11918_, _10762_);
  or (_11920_, _11919_, _11904_);
  or (_11921_, _09256_, _08787_);
  nor (_11922_, _09855_, _05801_);
  and (_11923_, _09239_, _05787_);
  nor (_11924_, _05799_, _05758_);
  not (_11925_, _11924_);
  or (_11926_, _09210_, _06070_);
  or (_11927_, _09025_, _06228_);
  and (_11928_, _11927_, _11926_);
  or (_11929_, _09211_, _06625_);
  or (_11930_, _09070_, _06626_);
  and (_11931_, _11930_, _11929_);
  and (_11932_, _11931_, _11928_);
  nand (_11933_, _09160_, _06107_);
  or (_11934_, _09115_, _06912_);
  nor (_11935_, _09114_, _09092_);
  or (_11936_, _11935_, _06913_);
  and (_11937_, _11936_, _11934_);
  and (_11938_, _11937_, _11933_);
  and (_11939_, _11938_, _11932_);
  or (_11940_, _09160_, _06107_);
  and (_11941_, _08838_, _06039_);
  nor (_11942_, _11941_, _08581_);
  or (_11943_, _09207_, _06203_);
  or (_11944_, _08883_, _07482_);
  and (_11945_, _11944_, _11943_);
  and (_11946_, _11945_, _11942_);
  or (_11947_, _08931_, _07805_);
  or (_11948_, _09208_, _06477_);
  and (_11949_, _11948_, _11947_);
  or (_11950_, _08980_, _07775_);
  or (_11951_, _09209_, _06876_);
  and (_11952_, _11951_, _11950_);
  and (_11953_, _11952_, _11949_);
  and (_11954_, _11953_, _11946_);
  and (_11955_, _11954_, _11940_);
  nand (_11956_, _11955_, _11939_);
  or (_11957_, _11956_, _09239_);
  and (_11958_, _11955_, _11939_);
  and (_11959_, _09242_, _09178_);
  and (_11960_, _11959_, \oc8051_golden_model_1.PC [11]);
  and (_11961_, _11960_, \oc8051_golden_model_1.PC [12]);
  and (_11962_, _11961_, \oc8051_golden_model_1.PC [13]);
  and (_11963_, _11962_, \oc8051_golden_model_1.PC [14]);
  nor (_11964_, _11962_, \oc8051_golden_model_1.PC [14]);
  nor (_11965_, _11964_, _11963_);
  not (_11966_, _11965_);
  nor (_11967_, _11966_, _08395_);
  and (_11968_, _11966_, _08395_);
  nor (_11969_, _11968_, _11967_);
  not (_11970_, _11969_);
  nor (_11971_, _11961_, \oc8051_golden_model_1.PC [13]);
  nor (_11972_, _11971_, _11962_);
  not (_11973_, _11972_);
  nor (_11974_, _11973_, _08395_);
  and (_11975_, _11973_, _08395_);
  nor (_11976_, _11960_, \oc8051_golden_model_1.PC [12]);
  nor (_11977_, _11976_, _11961_);
  not (_11978_, _11977_);
  nor (_11979_, _11978_, _08395_);
  nor (_11980_, _11959_, \oc8051_golden_model_1.PC [11]);
  nor (_11981_, _11980_, _11960_);
  not (_11982_, _11981_);
  nor (_11983_, _11982_, _08395_);
  and (_11984_, _11982_, _08395_);
  nor (_11985_, _11984_, _11983_);
  and (_11986_, _09231_, _09178_);
  nor (_11987_, _11986_, \oc8051_golden_model_1.PC [10]);
  nor (_11988_, _11987_, _11959_);
  not (_11989_, _11988_);
  nor (_11990_, _11989_, _08395_);
  and (_11991_, _11989_, _08395_);
  nor (_11992_, _11991_, _11990_);
  and (_11993_, _11992_, _11985_);
  and (_11994_, _09178_, \oc8051_golden_model_1.PC [8]);
  nor (_11995_, _11994_, \oc8051_golden_model_1.PC [9]);
  nor (_11996_, _11995_, _11986_);
  not (_11997_, _11996_);
  nor (_11998_, _11997_, _08395_);
  and (_11999_, _11997_, _08395_);
  nor (_12000_, _11999_, _11998_);
  nor (_12001_, _09181_, _08395_);
  and (_12002_, _09181_, _08395_);
  and (_12003_, _09176_, _08432_);
  nor (_12004_, _12003_, \oc8051_golden_model_1.PC [6]);
  nor (_12005_, _12004_, _09177_);
  not (_12006_, _12005_);
  nor (_12007_, _12006_, _08638_);
  and (_12008_, _12006_, _08638_);
  nor (_12009_, _12008_, _12007_);
  not (_12010_, _12009_);
  and (_12011_, _09176_, \oc8051_golden_model_1.PC [4]);
  nor (_12012_, _12011_, \oc8051_golden_model_1.PC [5]);
  nor (_12013_, _12012_, _12003_);
  not (_12014_, _12013_);
  nor (_12015_, _12014_, _08701_);
  and (_12016_, _12014_, _08701_);
  nor (_12017_, _09176_, \oc8051_golden_model_1.PC [4]);
  nor (_12018_, _12017_, _12011_);
  not (_12019_, _12018_);
  nor (_12020_, _12019_, _08670_);
  and (_12021_, _05449_, \oc8051_golden_model_1.PC [2]);
  nor (_12022_, _12021_, \oc8051_golden_model_1.PC [3]);
  nor (_12023_, _12022_, _09176_);
  not (_12024_, _12023_);
  nor (_12025_, _12024_, _06389_);
  and (_12026_, _12024_, _06389_);
  nor (_12027_, _05449_, \oc8051_golden_model_1.PC [2]);
  nor (_12028_, _12027_, _12021_);
  not (_12029_, _12028_);
  nor (_12030_, _12029_, _06521_);
  nor (_12031_, _06945_, _05879_);
  nor (_12032_, _06758_, \oc8051_golden_model_1.PC [0]);
  and (_12033_, _06945_, _05879_);
  nor (_12034_, _12033_, _12031_);
  and (_12035_, _12034_, _12032_);
  nor (_12036_, _12035_, _12031_);
  and (_12037_, _12029_, _06521_);
  nor (_12038_, _12037_, _12030_);
  not (_12039_, _12038_);
  nor (_12040_, _12039_, _12036_);
  nor (_12041_, _12040_, _12030_);
  nor (_12042_, _12041_, _12026_);
  nor (_12043_, _12042_, _12025_);
  and (_12044_, _12019_, _08670_);
  nor (_12045_, _12044_, _12020_);
  not (_12046_, _12045_);
  nor (_12047_, _12046_, _12043_);
  nor (_12048_, _12047_, _12020_);
  nor (_12049_, _12048_, _12016_);
  nor (_12050_, _12049_, _12015_);
  nor (_12051_, _12050_, _12010_);
  nor (_12052_, _12051_, _12007_);
  nor (_12053_, _12052_, _12002_);
  or (_12054_, _12053_, _12001_);
  nor (_12055_, _09178_, \oc8051_golden_model_1.PC [8]);
  nor (_12056_, _12055_, _11994_);
  not (_12057_, _12056_);
  nor (_12058_, _12057_, _08395_);
  and (_12059_, _12057_, _08395_);
  nor (_12060_, _12059_, _12058_);
  and (_12061_, _12060_, _12054_);
  and (_12062_, _12061_, _12000_);
  and (_12063_, _12062_, _11993_);
  nor (_12064_, _12058_, _11998_);
  not (_12065_, _12064_);
  and (_12066_, _12065_, _11993_);
  or (_12067_, _12066_, _11990_);
  or (_12068_, _12067_, _12063_);
  nor (_12069_, _12068_, _11983_);
  and (_12070_, _11978_, _08395_);
  nor (_12071_, _12070_, _11979_);
  not (_12072_, _12071_);
  nor (_12073_, _12072_, _12069_);
  nor (_12074_, _12073_, _11979_);
  nor (_12075_, _12074_, _11975_);
  nor (_12076_, _12075_, _11974_);
  nor (_12077_, _12076_, _11970_);
  nor (_12078_, _12077_, _11967_);
  and (_12079_, _09240_, _08395_);
  nor (_12080_, _09240_, _08395_);
  nor (_12081_, _12080_, _12079_);
  and (_12082_, _12081_, _12078_);
  nor (_12083_, _12081_, _12078_);
  nor (_12084_, _12083_, _12082_);
  not (_12085_, _12084_);
  or (_12086_, _12085_, _11958_);
  and (_12087_, _12086_, _06687_);
  and (_12088_, _12087_, _11957_);
  not (_12089_, _06687_);
  nor (_12090_, _07049_, _06107_);
  not (_12091_, _12090_);
  and (_12092_, _09194_, _06039_);
  and (_12093_, _08347_, _07482_);
  nor (_12094_, _12093_, _12092_);
  and (_12095_, _08012_, _06203_);
  and (_12096_, _08101_, _06477_);
  nor (_12097_, _12096_, _12095_);
  and (_12098_, _12097_, _12094_);
  and (_12099_, _08348_, _07805_);
  and (_12100_, _08349_, _07775_);
  nor (_12101_, _12100_, _12099_);
  and (_12102_, _08336_, _06876_);
  nor (_12103_, _12102_, _07924_);
  and (_12104_, _12103_, _12101_);
  and (_12105_, _12104_, _12098_);
  and (_12106_, _07474_, _06228_);
  and (_12107_, _07544_, _06070_);
  nor (_12108_, _12107_, _12106_);
  and (_12109_, _07657_, _06626_);
  and (_12110_, _07708_, _06625_);
  nor (_12111_, _12110_, _12109_);
  and (_12112_, _12111_, _12108_);
  and (_12113_, _07252_, _06913_);
  and (_12114_, _07306_, _06912_);
  and (_12115_, _07049_, _06107_);
  or (_12116_, _12115_, _12114_);
  nor (_12117_, _12116_, _12113_);
  and (_12118_, _12117_, _12112_);
  and (_12119_, _12118_, _12105_);
  and (_12120_, _12119_, _12091_);
  nand (_12121_, _12120_, _09240_);
  nand (_12122_, _06125_, _06144_);
  and (_12123_, _06119_, _06144_);
  nor (_12124_, _12123_, _06290_);
  and (_12125_, _12124_, _12122_);
  not (_12126_, _12125_);
  or (_12127_, _12120_, _12085_);
  and (_12128_, _12127_, _12126_);
  and (_12129_, _12128_, _12121_);
  and (_12130_, _09256_, _06220_);
  and (_12131_, _06221_, _05764_);
  or (_12132_, _12131_, _09256_);
  nor (_12133_, _05799_, _05762_);
  nor (_12134_, _12133_, _10490_);
  and (_12135_, _08211_, _08175_);
  and (_12136_, _08542_, _12135_);
  and (_12137_, _08014_, _07925_);
  and (_12138_, _12137_, _08539_);
  nand (_12139_, _12138_, _12136_);
  or (_12140_, _12139_, _09239_);
  and (_12141_, _12138_, _12136_);
  or (_12142_, _12141_, _12085_);
  and (_12143_, _12142_, _06160_);
  and (_12144_, _12143_, _12140_);
  nor (_12145_, _09246_, \oc8051_golden_model_1.PC [14]);
  nor (_12146_, _12145_, _09247_);
  and (_12147_, _12146_, _06039_);
  nor (_12148_, _12146_, _06039_);
  nor (_12149_, _12148_, _12147_);
  not (_12150_, _12149_);
  nor (_12151_, _09245_, \oc8051_golden_model_1.PC [13]);
  nor (_12152_, _12151_, _09246_);
  and (_12153_, _12152_, _06039_);
  nor (_12154_, _12152_, _06039_);
  nor (_12155_, _09244_, \oc8051_golden_model_1.PC [12]);
  nor (_12156_, _12155_, _09245_);
  and (_12157_, _12156_, _06039_);
  nor (_12158_, _09249_, \oc8051_golden_model_1.PC [10]);
  nor (_12159_, _12158_, _09250_);
  and (_12160_, _12159_, _06039_);
  not (_12161_, _12160_);
  nor (_12162_, _09250_, \oc8051_golden_model_1.PC [11]);
  nor (_12163_, _12162_, _09251_);
  and (_12164_, _12163_, _06039_);
  nor (_12165_, _12163_, _06039_);
  nor (_12166_, _12165_, _12164_);
  nor (_12167_, _12159_, _06039_);
  nor (_12168_, _12167_, _12160_);
  and (_12169_, _12168_, _12166_);
  and (_12170_, _08435_, \oc8051_golden_model_1.PC [8]);
  nor (_12171_, _12170_, \oc8051_golden_model_1.PC [9]);
  nor (_12172_, _12171_, _09249_);
  and (_12173_, _12172_, _06039_);
  nor (_12174_, _12172_, _06039_);
  nor (_12175_, _12174_, _12173_);
  and (_12176_, _08437_, _06039_);
  nor (_12177_, _08437_, _06039_);
  and (_12178_, _08432_, _05972_);
  nor (_12179_, _12178_, \oc8051_golden_model_1.PC [6]);
  nor (_12180_, _12179_, _08434_);
  not (_12181_, _12180_);
  nor (_12182_, _12181_, _06203_);
  and (_12183_, _12181_, _06203_);
  nor (_12184_, _12183_, _12182_);
  not (_12185_, _12184_);
  and (_12186_, _05972_, \oc8051_golden_model_1.PC [4]);
  nor (_12187_, _12186_, \oc8051_golden_model_1.PC [5]);
  nor (_12188_, _12187_, _12178_);
  not (_12189_, _12188_);
  nor (_12190_, _12189_, _06477_);
  and (_12191_, _12189_, _06477_);
  nor (_12192_, _05972_, \oc8051_golden_model_1.PC [4]);
  nor (_12193_, _12192_, _12186_);
  not (_12194_, _12193_);
  nor (_12195_, _12194_, _06876_);
  nor (_12196_, _06070_, _06322_);
  and (_12197_, _06070_, _06322_);
  nor (_12198_, _06625_, _05923_);
  nor (_12199_, _06912_, \oc8051_golden_model_1.PC [1]);
  nor (_12200_, _06107_, _05444_);
  and (_12201_, _06912_, \oc8051_golden_model_1.PC [1]);
  nor (_12202_, _12201_, _12199_);
  and (_12203_, _12202_, _12200_);
  nor (_12204_, _12203_, _12199_);
  and (_12205_, _06625_, _05923_);
  nor (_12206_, _12205_, _12198_);
  not (_12207_, _12206_);
  nor (_12208_, _12207_, _12204_);
  nor (_12209_, _12208_, _12198_);
  nor (_12210_, _12209_, _12197_);
  nor (_12211_, _12210_, _12196_);
  and (_12212_, _12194_, _06876_);
  nor (_12213_, _12212_, _12195_);
  not (_12214_, _12213_);
  nor (_12215_, _12214_, _12211_);
  nor (_12216_, _12215_, _12195_);
  nor (_12217_, _12216_, _12191_);
  nor (_12218_, _12217_, _12190_);
  nor (_12219_, _12218_, _12185_);
  nor (_12220_, _12219_, _12182_);
  nor (_12221_, _12220_, _12177_);
  or (_12222_, _12221_, _12176_);
  nor (_12223_, _08435_, \oc8051_golden_model_1.PC [8]);
  nor (_12224_, _12223_, _12170_);
  and (_12225_, _12224_, _06039_);
  nor (_12226_, _12224_, _06039_);
  nor (_12227_, _12226_, _12225_);
  and (_12228_, _12227_, _12222_);
  and (_12229_, _12228_, _12175_);
  and (_12230_, _12229_, _12169_);
  nor (_12231_, _12225_, _12173_);
  not (_12232_, _12231_);
  and (_12233_, _12232_, _12169_);
  or (_12234_, _12233_, _12164_);
  nor (_12235_, _12234_, _12230_);
  and (_12236_, _12235_, _12161_);
  nor (_12237_, _12156_, _06039_);
  nor (_12238_, _12237_, _12157_);
  not (_12239_, _12238_);
  nor (_12240_, _12239_, _12236_);
  nor (_12241_, _12240_, _12157_);
  nor (_12242_, _12241_, _12154_);
  nor (_12243_, _12242_, _12153_);
  nor (_12244_, _12243_, _12150_);
  nor (_12245_, _12244_, _12147_);
  nor (_12246_, _09256_, _06039_);
  and (_12247_, _09256_, _06039_);
  nor (_12248_, _12247_, _12246_);
  and (_12249_, _12248_, _12245_);
  nor (_12250_, _12248_, _12245_);
  or (_12251_, _12250_, _12249_);
  and (_12252_, _07252_, _07049_);
  and (_12253_, _08347_, _09194_);
  and (_12254_, _12253_, _12252_);
  and (_12255_, _08351_, _08350_);
  nand (_12256_, _12255_, _12254_);
  and (_12257_, _12256_, _12251_);
  and (_12258_, _12255_, _12254_);
  and (_12259_, _12258_, _09256_);
  or (_12260_, _12259_, _08443_);
  or (_12261_, _12260_, _12257_);
  nor (_12262_, _10473_, _10483_);
  and (_12263_, _12262_, _10471_);
  not (_12264_, _06653_);
  nor (_12265_, _07382_, _07372_);
  and (_12266_, _12265_, _12264_);
  and (_12267_, _12266_, _12263_);
  not (_12268_, _12267_);
  and (_12269_, _12268_, _11904_);
  and (_12270_, _09256_, _06581_);
  and (_12271_, _09256_, _07056_);
  nor (_12272_, _06581_, _09229_);
  and (_12273_, _12272_, _07057_);
  and (_12274_, _12273_, _12265_);
  or (_12275_, _12274_, _12271_);
  and (_12276_, _12275_, _12264_);
  or (_12277_, _12276_, _12270_);
  and (_12278_, _12277_, _12263_);
  or (_12279_, _12278_, _08445_);
  or (_12280_, _12279_, _12269_);
  nor (_12281_, _07064_, _06160_);
  and (_12282_, _12281_, _12280_);
  and (_12283_, _12282_, _12261_);
  or (_12284_, _12283_, _12144_);
  and (_12285_, _12284_, _12134_);
  not (_12286_, _12131_);
  nand (_12287_, _12134_, _07065_);
  and (_12288_, _12287_, _11904_);
  or (_12289_, _12288_, _12286_);
  or (_12290_, _12289_, _12285_);
  and (_12291_, _12290_, _12132_);
  and (_12292_, _10458_, _07082_);
  not (_12293_, _12292_);
  or (_12294_, _12293_, _12291_);
  or (_12295_, _12292_, _11904_);
  and (_12296_, _12295_, _06229_);
  and (_12297_, _12296_, _12294_);
  or (_12298_, _12297_, _12130_);
  nor (_12299_, _05799_, _05768_);
  nor (_12300_, _12299_, _10525_);
  and (_12301_, _12300_, _12298_);
  not (_12302_, _12300_);
  and (_12303_, _12302_, _11904_);
  not (_12304_, _05769_);
  nor (_12305_, _06151_, _12304_);
  and (_12306_, _12305_, _06153_);
  not (_12307_, _12306_);
  or (_12308_, _12307_, _12303_);
  or (_12309_, _12308_, _12301_);
  or (_12310_, _12306_, _09256_);
  and (_12311_, _12310_, _12125_);
  and (_12312_, _12311_, _12309_);
  or (_12313_, _12312_, _12129_);
  and (_12314_, _12313_, _12089_);
  or (_12315_, _12314_, _06236_);
  or (_12316_, _12315_, _12088_);
  not (_12317_, _06295_);
  nor (_12318_, _10273_, _10272_);
  nor (_12319_, _12318_, _10282_);
  not (_12320_, _10278_);
  nor (_12321_, _08211_, \oc8051_golden_model_1.ACC [0]);
  or (_12322_, _12321_, _10276_);
  and (_12323_, _12322_, _12320_);
  and (_12324_, _12323_, _12319_);
  nor (_12325_, _10268_, _10269_);
  nor (_12326_, _12325_, _10289_);
  nor (_12327_, _10295_, _08810_);
  and (_12328_, _12327_, _12326_);
  and (_12329_, _12328_, _12324_);
  and (_12330_, _12329_, _09239_);
  nor (_12331_, _12329_, _12084_);
  or (_12332_, _12331_, _06643_);
  or (_12333_, _12332_, _12330_);
  and (_12334_, _12333_, _12317_);
  and (_12335_, _12334_, _12316_);
  nor (_12336_, _11059_, _11060_);
  nor (_12337_, _12336_, _11063_);
  and (_12338_, _06107_, _05855_);
  nor (_12339_, _12338_, _11067_);
  nor (_12340_, _12339_, _11066_);
  and (_12341_, _12340_, _12337_);
  nor (_12342_, _11053_, _11054_);
  nor (_12343_, _12342_, _11058_);
  nor (_12344_, _11052_, _10794_);
  and (_12345_, _12344_, _12343_);
  and (_12346_, _12345_, _12341_);
  not (_12347_, _12346_);
  nand (_12348_, _12347_, _12084_);
  nand (_12349_, _12346_, _09240_);
  and (_12350_, _12349_, _06295_);
  and (_12351_, _12350_, _12348_);
  or (_12352_, _12351_, _12335_);
  and (_12353_, _12352_, _11925_);
  nand (_12354_, _11924_, _11904_);
  and (_12355_, _06124_, _06245_);
  nor (_12356_, _12355_, _06212_);
  nor (_12357_, _06701_, _07388_);
  and (_12358_, _06128_, _06245_);
  not (_12359_, _12358_);
  nor (_12360_, _07292_, _06145_);
  and (_12361_, _12360_, _12359_);
  and (_12362_, _12361_, _12357_);
  and (_12363_, _12362_, _12356_);
  nand (_12364_, _12363_, _12354_);
  or (_12365_, _12364_, _12353_);
  and (_12366_, _05786_, _06245_);
  not (_12367_, _12366_);
  nor (_12368_, _11311_, _09295_);
  and (_12369_, _12368_, _12367_);
  or (_12370_, _12363_, _09256_);
  and (_12371_, _12370_, _12369_);
  and (_12372_, _12371_, _12365_);
  not (_12373_, _12369_);
  and (_12374_, _12373_, _11904_);
  and (_12375_, _06256_, _05775_);
  not (_12376_, _12375_);
  or (_12377_, _12376_, _12374_);
  or (_12378_, _12377_, _12372_);
  and (_12379_, _06115_, _05790_);
  not (_12380_, _12379_);
  and (_12381_, _10554_, _12380_);
  or (_12382_, _12375_, _09256_);
  and (_12383_, _12382_, _12381_);
  and (_12384_, _12383_, _12378_);
  nor (_12385_, _10387_, _06260_);
  not (_12386_, _12385_);
  not (_12387_, _12381_);
  and (_12388_, _12387_, _11904_);
  or (_12389_, _12388_, _12386_);
  or (_12390_, _12389_, _12384_);
  or (_12391_, _12385_, _09256_);
  and (_12392_, _12391_, _05805_);
  and (_12393_, _12392_, _12390_);
  and (_12394_, _11904_, _05870_);
  nor (_12395_, _06139_, _05791_);
  not (_12396_, _12395_);
  or (_12397_, _12396_, _12394_);
  or (_12398_, _12397_, _12393_);
  or (_12399_, _12395_, _09256_);
  and (_12400_, _12399_, _11296_);
  and (_12401_, _12400_, _12398_);
  nand (_12402_, _09239_, _06293_);
  nand (_12403_, _12402_, _06133_);
  or (_12404_, _12403_, _12401_);
  or (_12405_, _09256_, _06133_);
  and (_12406_, _12405_, _06114_);
  and (_12407_, _12406_, _12404_);
  or (_12408_, _12407_, _11923_);
  and (_12409_, _12408_, _11922_);
  nor (_12410_, _06209_, _05829_);
  not (_12411_, _12410_);
  not (_12412_, _11922_);
  and (_12413_, _12412_, _11904_);
  or (_12414_, _12413_, _12411_);
  or (_12415_, _12414_, _12409_);
  and (_12416_, _05781_, _05746_);
  not (_12417_, _12416_);
  or (_12418_, _12410_, _09256_);
  and (_12419_, _12418_, _12417_);
  and (_12420_, _12419_, _12415_);
  and (_12421_, _12416_, _12251_);
  or (_12422_, _12421_, _08788_);
  or (_12423_, _12422_, _12420_);
  and (_12424_, _12423_, _11921_);
  or (_12425_, _12424_, _06110_);
  nand (_12426_, _09240_, _06110_);
  and (_12427_, _12426_, _10752_);
  and (_12428_, _12427_, _12425_);
  and (_12429_, _10751_, _09256_);
  or (_12430_, _12429_, _12428_);
  nor (_12431_, _05835_, _05799_);
  not (_12432_, _12431_);
  and (_12433_, _12432_, _12430_);
  not (_12434_, \oc8051_golden_model_1.DPH [0]);
  and (_12435_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_12436_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_12437_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_12438_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_12439_, _12438_, _12437_);
  not (_12440_, _12439_);
  and (_12441_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_12442_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_12443_, _12442_, _12441_);
  not (_12444_, _12443_);
  and (_12445_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_12446_, _05966_, _05962_);
  nor (_12447_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_12448_, _12447_, _12445_);
  not (_12449_, _12448_);
  nor (_12450_, _12449_, _12446_);
  nor (_12451_, _12450_, _12445_);
  nor (_12452_, _12451_, _12444_);
  nor (_12453_, _12452_, _12441_);
  nor (_12454_, _12453_, _12440_);
  nor (_12455_, _12454_, _12437_);
  nor (_12456_, _12455_, _12436_);
  nor (_12457_, _12456_, _12435_);
  nor (_12458_, _12457_, _12434_);
  and (_12459_, _12458_, \oc8051_golden_model_1.DPH [1]);
  and (_12460_, _12459_, \oc8051_golden_model_1.DPH [2]);
  and (_12461_, _12460_, \oc8051_golden_model_1.DPH [3]);
  and (_12462_, _12461_, \oc8051_golden_model_1.DPH [4]);
  and (_12463_, _12462_, \oc8051_golden_model_1.DPH [5]);
  and (_12464_, _12463_, \oc8051_golden_model_1.DPH [6]);
  nand (_12465_, _12464_, \oc8051_golden_model_1.DPH [7]);
  or (_12466_, _12464_, \oc8051_golden_model_1.DPH [7]);
  and (_12467_, _12466_, _12431_);
  and (_12468_, _12467_, _12465_);
  nor (_12469_, _06208_, _06076_);
  not (_12470_, _12469_);
  or (_12471_, _12470_, _12468_);
  or (_12472_, _12471_, _12433_);
  and (_12473_, _06109_, _05746_);
  not (_12474_, _12473_);
  or (_12475_, _12469_, _09256_);
  and (_12476_, _12475_, _12474_);
  and (_12477_, _12476_, _12472_);
  not (_12478_, _11919_);
  or (_12479_, _12251_, _11101_);
  not (_12480_, _11101_);
  or (_12481_, _12480_, _09256_);
  and (_12482_, _12481_, _12473_);
  and (_12483_, _12482_, _12479_);
  or (_12484_, _12483_, _12478_);
  or (_12485_, _12484_, _12477_);
  and (_12486_, _12485_, _11920_);
  or (_12487_, _12486_, _11917_);
  or (_12488_, _11916_, _09256_);
  and (_12489_, _12488_, _07127_);
  and (_12490_, _12489_, _12487_);
  nand (_12491_, _09239_, _06297_);
  not (_12492_, _05834_);
  nor (_12493_, _06402_, _12492_);
  nand (_12494_, _12493_, _12491_);
  or (_12495_, _12494_, _12490_);
  and (_12496_, _06399_, _05746_);
  not (_12497_, _12496_);
  or (_12498_, _12493_, _09256_);
  and (_12499_, _12498_, _12497_);
  and (_12500_, _12499_, _12495_);
  or (_12501_, _12251_, _12480_);
  or (_12502_, _11101_, _09256_);
  and (_12503_, _12502_, _12496_);
  and (_12504_, _12503_, _12501_);
  not (_12505_, _11914_);
  or (_12506_, _12505_, _12504_);
  or (_12507_, _12506_, _12500_);
  and (_12508_, _12507_, _11915_);
  or (_12509_, _12508_, _10822_);
  or (_12510_, _10821_, _09256_);
  and (_12511_, _12510_, _07132_);
  and (_12512_, _12511_, _12509_);
  nand (_12513_, _09239_, _06306_);
  nor (_12514_, _06411_, _07124_);
  nand (_12515_, _12514_, _12513_);
  or (_12516_, _12515_, _12512_);
  and (_12517_, _06408_, _05746_);
  not (_12518_, _12517_);
  or (_12519_, _12514_, _09256_);
  and (_12520_, _12519_, _12518_);
  and (_12521_, _12520_, _12516_);
  not (_12522_, _11912_);
  or (_12523_, _12251_, \oc8051_golden_model_1.PSW [7]);
  or (_12524_, _09256_, _10693_);
  and (_12525_, _12524_, _12517_);
  and (_12526_, _12525_, _12523_);
  or (_12527_, _12526_, _12522_);
  or (_12528_, _12527_, _12521_);
  and (_12529_, _12528_, _11913_);
  or (_12530_, _12529_, _10850_);
  or (_12531_, _10849_, _09256_);
  and (_12532_, _12531_, _08819_);
  and (_12533_, _12532_, _12530_);
  nand (_12534_, _09239_, _06303_);
  nor (_12535_, _06396_, _05842_);
  nand (_12536_, _12535_, _12534_);
  or (_12537_, _12536_, _12533_);
  and (_12538_, _05840_, _05746_);
  not (_12539_, _12538_);
  or (_12540_, _12535_, _09256_);
  and (_12541_, _12540_, _12539_);
  and (_12542_, _12541_, _12537_);
  or (_12543_, _12251_, _10693_);
  or (_12544_, _09256_, \oc8051_golden_model_1.PSW [7]);
  and (_12545_, _12544_, _12538_);
  and (_12546_, _12545_, _12543_);
  not (_12547_, _11907_);
  or (_12548_, _12547_, _12546_);
  or (_12549_, _12548_, _12542_);
  and (_12550_, _12549_, _11908_);
  or (_12551_, _12550_, _10897_);
  or (_12552_, _10896_, _09256_);
  and (_12553_, _12552_, _10926_);
  and (_12554_, _12553_, _12551_);
  and (_12555_, _11904_, _10925_);
  or (_12556_, _12555_, _06417_);
  or (_12557_, _12556_, _12554_);
  not (_12558_, _06417_);
  or (_12559_, _07923_, _12558_);
  and (_12560_, _12559_, _12557_);
  or (_12561_, _12560_, _07142_);
  nor (_12562_, _09256_, _05846_);
  nor (_12563_, _12562_, _06301_);
  and (_12564_, _12563_, _12561_);
  not (_12565_, _11905_);
  and (_12566_, _08415_, \oc8051_golden_model_1.IP [6]);
  and (_12567_, _08418_, \oc8051_golden_model_1.IE [6]);
  and (_12568_, _08409_, \oc8051_golden_model_1.ACC [6]);
  or (_12569_, _12568_, _12567_);
  or (_12570_, _12569_, _12566_);
  and (_12571_, _08413_, \oc8051_golden_model_1.SCON [6]);
  and (_12572_, _08404_, \oc8051_golden_model_1.PSW [6]);
  or (_12573_, _12572_, _12571_);
  and (_12574_, _08407_, \oc8051_golden_model_1.TCON [6]);
  and (_12575_, _08420_, \oc8051_golden_model_1.B [6]);
  or (_12576_, _12575_, _12574_);
  or (_12577_, _12576_, _12573_);
  or (_12578_, _12577_, _12570_);
  or (_12579_, _12578_, _08013_);
  and (_12580_, _07800_, _06626_);
  and (_12581_, _12580_, _12579_);
  and (_12582_, _08415_, \oc8051_golden_model_1.IP [3]);
  and (_12583_, _08420_, \oc8051_golden_model_1.B [3]);
  and (_12584_, _08409_, \oc8051_golden_model_1.ACC [3]);
  or (_12585_, _12584_, _12583_);
  or (_12586_, _12585_, _12582_);
  and (_12587_, _08407_, \oc8051_golden_model_1.TCON [3]);
  and (_12588_, _08413_, \oc8051_golden_model_1.SCON [3]);
  or (_12589_, _12588_, _12587_);
  and (_12590_, _08418_, \oc8051_golden_model_1.IE [3]);
  and (_12591_, _08404_, \oc8051_golden_model_1.PSW [3]);
  or (_12592_, _12591_, _12590_);
  or (_12593_, _12592_, _12589_);
  or (_12594_, _12593_, _12586_);
  or (_12595_, _12594_, _08138_);
  and (_12596_, _12595_, _07851_);
  nor (_12597_, _12596_, _12581_);
  and (_12598_, _08413_, \oc8051_golden_model_1.SCON [5]);
  and (_12599_, _08418_, \oc8051_golden_model_1.IE [5]);
  and (_12600_, _08409_, \oc8051_golden_model_1.ACC [5]);
  or (_12601_, _12600_, _12599_);
  or (_12602_, _12601_, _12598_);
  and (_12603_, _08404_, \oc8051_golden_model_1.PSW [5]);
  and (_12604_, _08420_, \oc8051_golden_model_1.B [5]);
  or (_12605_, _12604_, _12603_);
  and (_12606_, _08407_, \oc8051_golden_model_1.TCON [5]);
  and (_12607_, _08415_, \oc8051_golden_model_1.IP [5]);
  or (_12608_, _12607_, _12606_);
  or (_12609_, _12608_, _12605_);
  or (_12610_, _12609_, _12602_);
  or (_12611_, _12610_, _08102_);
  and (_12612_, _07780_, _06626_);
  and (_12613_, _12612_, _12611_);
  and (_12614_, _08409_, \oc8051_golden_model_1.ACC [1]);
  and (_12615_, _08415_, \oc8051_golden_model_1.IP [1]);
  and (_12616_, _08420_, \oc8051_golden_model_1.B [1]);
  or (_12617_, _12616_, _12615_);
  or (_12618_, _12617_, _12614_);
  and (_12619_, _08407_, \oc8051_golden_model_1.TCON [1]);
  and (_12620_, _08413_, \oc8051_golden_model_1.SCON [1]);
  or (_12621_, _12620_, _12619_);
  and (_12622_, _08418_, \oc8051_golden_model_1.IE [1]);
  and (_12623_, _08404_, \oc8051_golden_model_1.PSW [1]);
  or (_12624_, _12623_, _12622_);
  or (_12625_, _12624_, _12621_);
  or (_12626_, _12625_, _12618_);
  or (_12627_, _12626_, _08174_);
  and (_12628_, _12627_, _07781_);
  nor (_12629_, _12628_, _12613_);
  and (_12630_, _12629_, _12597_);
  and (_12631_, _08413_, \oc8051_golden_model_1.SCON [2]);
  and (_12632_, _08407_, \oc8051_golden_model_1.TCON [2]);
  and (_12633_, _08409_, \oc8051_golden_model_1.ACC [2]);
  or (_12634_, _12633_, _12632_);
  or (_12635_, _12634_, _12631_);
  and (_12636_, _08404_, \oc8051_golden_model_1.PSW [2]);
  and (_12637_, _08420_, \oc8051_golden_model_1.B [2]);
  or (_12638_, _12637_, _12636_);
  and (_12639_, _08418_, \oc8051_golden_model_1.IE [2]);
  and (_12640_, _08415_, \oc8051_golden_model_1.IP [2]);
  or (_12641_, _12640_, _12639_);
  or (_12642_, _12641_, _12638_);
  or (_12643_, _12642_, _12635_);
  or (_12644_, _12643_, _08246_);
  and (_12645_, _12644_, _07848_);
  nor (_12646_, _12645_, _08567_);
  and (_12647_, _08413_, \oc8051_golden_model_1.SCON [0]);
  and (_12648_, _08407_, \oc8051_golden_model_1.TCON [0]);
  and (_12649_, _08409_, \oc8051_golden_model_1.ACC [0]);
  or (_12650_, _12649_, _12648_);
  or (_12651_, _12650_, _12647_);
  and (_12652_, _08415_, \oc8051_golden_model_1.IP [0]);
  and (_12653_, _08420_, \oc8051_golden_model_1.B [0]);
  or (_12654_, _12653_, _12652_);
  and (_12655_, _08418_, \oc8051_golden_model_1.IE [0]);
  and (_12656_, _08404_, \oc8051_golden_model_1.PSW [0]);
  or (_12657_, _12656_, _12655_);
  or (_12658_, _12657_, _12654_);
  or (_12659_, _12658_, _12651_);
  or (_12660_, _12659_, _08210_);
  and (_12661_, _12660_, _07772_);
  and (_12662_, _08420_, \oc8051_golden_model_1.B [4]);
  and (_12663_, _08413_, \oc8051_golden_model_1.SCON [4]);
  and (_12664_, _08418_, \oc8051_golden_model_1.IE [4]);
  or (_12665_, _12664_, _12663_);
  or (_12666_, _12665_, _12662_);
  and (_12667_, _08415_, \oc8051_golden_model_1.IP [4]);
  and (_12668_, _08404_, \oc8051_golden_model_1.PSW [4]);
  or (_12669_, _12668_, _12667_);
  and (_12670_, _08407_, \oc8051_golden_model_1.TCON [4]);
  and (_12671_, _08409_, \oc8051_golden_model_1.ACC [4]);
  or (_12672_, _12671_, _12670_);
  or (_12673_, _12672_, _12669_);
  nor (_12674_, _12673_, _12666_);
  not (_12675_, _12674_);
  nor (_12676_, _12675_, _08337_);
  and (_12677_, _07771_, _06626_);
  not (_12678_, _12677_);
  nor (_12679_, _12678_, _12676_);
  nor (_12680_, _12679_, _12661_);
  and (_12681_, _12680_, _12646_);
  and (_12682_, _12681_, _12630_);
  nand (_12683_, _12084_, _12682_);
  or (_12684_, _09239_, _12682_);
  and (_12685_, _12684_, _06301_);
  and (_12686_, _12685_, _12683_);
  or (_12687_, _12686_, _12565_);
  or (_12688_, _12687_, _12564_);
  and (_12689_, _12688_, _11906_);
  nor (_12690_, _10264_, _06169_);
  not (_12691_, _12690_);
  or (_12692_, _12691_, _12689_);
  not (_12693_, _10262_);
  or (_12694_, _12690_, _09256_);
  and (_12695_, _12694_, _12693_);
  and (_12696_, _12695_, _12692_);
  and (_12697_, _11904_, _10262_);
  or (_12698_, _12697_, _06167_);
  or (_12699_, _12698_, _12696_);
  or (_12700_, _07923_, _06168_);
  and (_12701_, _12700_, _12699_);
  or (_12702_, _12701_, _05826_);
  not (_12703_, _05826_);
  or (_12704_, _09256_, _12703_);
  and (_12705_, _12704_, _06166_);
  and (_12706_, _12705_, _12702_);
  or (_12707_, _12085_, _12682_);
  nand (_12708_, _09240_, _12682_);
  and (_12709_, _12708_, _12707_);
  and (_12710_, _12709_, _06165_);
  and (_12711_, _08362_, _07154_);
  not (_12712_, _12711_);
  or (_12713_, _12712_, _12710_);
  or (_12714_, _12713_, _12706_);
  or (_12716_, _12711_, _11904_);
  and (_12717_, _12716_, _06829_);
  and (_12718_, _12717_, _12714_);
  nor (_12719_, _11094_, _11089_);
  nand (_12720_, _09256_, _06433_);
  nand (_12721_, _12720_, _12719_);
  or (_12722_, _12721_, _12718_);
  not (_12723_, _06310_);
  or (_12724_, _11904_, _12719_);
  and (_12725_, _12724_, _12723_);
  and (_12726_, _12725_, _12722_);
  and (_12727_, _06310_, _06039_);
  or (_12728_, _12727_, _05823_);
  or (_12729_, _12728_, _12726_);
  not (_12730_, _05823_);
  or (_12731_, _09256_, _12730_);
  and (_12732_, _12731_, _05749_);
  and (_12733_, _12732_, _12729_);
  and (_12734_, _12709_, _05748_);
  nor (_12735_, _09189_, _07168_);
  not (_12737_, _12735_);
  or (_12738_, _12737_, _12734_);
  or (_12739_, _12738_, _12733_);
  or (_12740_, _12735_, _11904_);
  and (_12741_, _12740_, _06444_);
  and (_12742_, _12741_, _12739_);
  nand (_12743_, _09256_, _06440_);
  nor (_12744_, _11119_, _11112_);
  nand (_12745_, _12744_, _12743_);
  or (_12746_, _12745_, _12742_);
  not (_12747_, _06305_);
  or (_12748_, _12744_, _11904_);
  and (_12749_, _12748_, _12747_);
  and (_12750_, _12749_, _12746_);
  and (_12751_, _06305_, _06039_);
  or (_12752_, _12751_, _05821_);
  or (_12753_, _12752_, _12750_);
  and (_12754_, _05820_, _05746_);
  not (_12755_, _12754_);
  or (_12756_, _09256_, _05822_);
  and (_12757_, _12756_, _12755_);
  and (_12758_, _12757_, _12753_);
  and (_12759_, _12754_, _11904_);
  or (_12760_, _12759_, _12758_);
  or (_12761_, _12760_, _01321_);
  or (_12762_, _01317_, \oc8051_golden_model_1.PC [15]);
  and (_12763_, _12762_, _43100_);
  and (_40993_, _12763_, _12761_);
  nor (_12764_, \oc8051_golden_model_1.P2 [7], rst);
  nor (_12765_, _12764_, _00000_);
  not (_12766_, \oc8051_golden_model_1.P2 [7]);
  not (_12767_, _07825_);
  nor (_12768_, _12767_, _07790_);
  nor (_12769_, _12768_, _12766_);
  and (_12770_, _12768_, _07923_);
  or (_12771_, _12770_, _12769_);
  or (_12772_, _12771_, _06132_);
  and (_12773_, _08403_, _07825_);
  nor (_12774_, _12773_, _12766_);
  and (_12775_, _07847_, \oc8051_golden_model_1.P0 [7]);
  and (_12776_, _12773_, \oc8051_golden_model_1.P2 [7]);
  or (_12777_, _12776_, _12775_);
  and (_12778_, _08403_, _07777_);
  and (_12779_, _12778_, \oc8051_golden_model_1.P1 [7]);
  and (_12780_, _08403_, _07829_);
  and (_12781_, _12780_, \oc8051_golden_model_1.P3 [7]);
  or (_12782_, _12781_, _12779_);
  or (_12783_, _12782_, _12777_);
  or (_12784_, _12783_, _08425_);
  and (_12785_, _12784_, _08399_);
  and (_12786_, _12785_, _12773_);
  or (_12787_, _12786_, _12774_);
  and (_12788_, _12787_, _06152_);
  and (_12789_, _07847_, _07772_);
  and (_12790_, _12789_, \oc8051_golden_model_1.P0 [7]);
  not (_12791_, _07777_);
  nor (_12792_, _07790_, _12791_);
  and (_12793_, _12792_, \oc8051_golden_model_1.P1 [7]);
  nor (_12794_, _12793_, _12790_);
  and (_12795_, _12768_, \oc8051_golden_model_1.P2 [7]);
  not (_12796_, _07829_);
  nor (_12797_, _12796_, _07790_);
  and (_12798_, _12797_, \oc8051_golden_model_1.P3 [7]);
  nor (_12799_, _12798_, _12795_);
  and (_12800_, _12799_, _12794_);
  and (_12801_, _12800_, _07925_);
  not (_12802_, _12801_);
  and (_12803_, _12797_, \oc8051_golden_model_1.P3 [6]);
  and (_12804_, _12792_, \oc8051_golden_model_1.P1 [6]);
  or (_12805_, _12804_, _12803_);
  and (_12806_, _12789_, \oc8051_golden_model_1.P0 [6]);
  and (_12807_, _12768_, \oc8051_golden_model_1.P2 [6]);
  or (_12808_, _12807_, _12806_);
  nor (_12809_, _12808_, _12805_);
  nand (_12810_, _12809_, _08014_);
  and (_12811_, _12797_, \oc8051_golden_model_1.P3 [5]);
  and (_12812_, _12792_, \oc8051_golden_model_1.P1 [5]);
  or (_12813_, _12812_, _12811_);
  and (_12814_, _12789_, \oc8051_golden_model_1.P0 [5]);
  and (_12815_, _12768_, \oc8051_golden_model_1.P2 [5]);
  or (_12816_, _12815_, _12814_);
  nor (_12817_, _12816_, _12813_);
  nand (_12818_, _12817_, _08103_);
  and (_12819_, _12797_, \oc8051_golden_model_1.P3 [4]);
  and (_12820_, _12792_, \oc8051_golden_model_1.P1 [4]);
  or (_12821_, _12820_, _12819_);
  and (_12822_, _12789_, \oc8051_golden_model_1.P0 [4]);
  and (_12823_, _12768_, \oc8051_golden_model_1.P2 [4]);
  or (_12824_, _12823_, _12822_);
  nor (_12825_, _12824_, _12821_);
  nand (_12826_, _12825_, _08338_);
  and (_12827_, _12797_, \oc8051_golden_model_1.P3 [3]);
  and (_12828_, _12792_, \oc8051_golden_model_1.P1 [3]);
  or (_12829_, _12828_, _12827_);
  and (_12830_, _12789_, \oc8051_golden_model_1.P0 [3]);
  and (_12831_, _12768_, \oc8051_golden_model_1.P2 [3]);
  or (_12832_, _12831_, _12830_);
  nor (_12833_, _12832_, _12829_);
  nand (_12834_, _12833_, _08139_);
  and (_12835_, _12797_, \oc8051_golden_model_1.P3 [2]);
  and (_12836_, _12792_, \oc8051_golden_model_1.P1 [2]);
  or (_12837_, _12836_, _12835_);
  and (_12838_, _12789_, \oc8051_golden_model_1.P0 [2]);
  and (_12839_, _12768_, \oc8051_golden_model_1.P2 [2]);
  or (_12840_, _12839_, _12838_);
  nor (_12841_, _12840_, _12837_);
  nand (_12842_, _12841_, _08247_);
  and (_12843_, _12789_, \oc8051_golden_model_1.P0 [1]);
  and (_12844_, _12792_, \oc8051_golden_model_1.P1 [1]);
  or (_12845_, _12844_, _12843_);
  and (_12846_, _12768_, \oc8051_golden_model_1.P2 [1]);
  and (_12847_, _12797_, \oc8051_golden_model_1.P3 [1]);
  or (_12848_, _12847_, _12846_);
  nor (_12849_, _12848_, _12845_);
  nand (_12850_, _12849_, _08175_);
  and (_12851_, _12789_, \oc8051_golden_model_1.P0 [0]);
  and (_12852_, _12792_, \oc8051_golden_model_1.P1 [0]);
  or (_12853_, _12852_, _12851_);
  and (_12854_, _12768_, \oc8051_golden_model_1.P2 [0]);
  and (_12855_, _12797_, \oc8051_golden_model_1.P3 [0]);
  or (_12856_, _12855_, _12854_);
  or (_12857_, _12856_, _12853_);
  or (_12858_, _12857_, _08211_);
  or (_12859_, _12858_, _12850_);
  nor (_12860_, _12859_, _12842_);
  not (_12861_, _12860_);
  nor (_12862_, _12861_, _12834_);
  not (_12863_, _12862_);
  nor (_12864_, _12863_, _12826_);
  not (_12865_, _12864_);
  nor (_12866_, _12865_, _12818_);
  not (_12867_, _12866_);
  nor (_12868_, _12867_, _12810_);
  or (_12869_, _12868_, _12802_);
  nand (_12870_, _12868_, _12802_);
  and (_12871_, _12870_, _12869_);
  and (_12872_, _12871_, _12768_);
  or (_12873_, _12872_, _12769_);
  or (_12874_, _12873_, _06161_);
  and (_12875_, _12768_, \oc8051_golden_model_1.ACC [7]);
  or (_12876_, _12875_, _12769_);
  and (_12877_, _12876_, _07056_);
  nor (_12878_, _07056_, _12766_);
  or (_12879_, _12878_, _06160_);
  or (_12880_, _12879_, _12877_);
  and (_12881_, _12880_, _06157_);
  and (_12882_, _12881_, _12874_);
  or (_12883_, _12783_, _08552_);
  and (_12884_, _12883_, _12773_);
  or (_12885_, _12884_, _12774_);
  and (_12886_, _12885_, _06156_);
  or (_12887_, _12886_, _06217_);
  or (_12888_, _12887_, _12882_);
  or (_12889_, _12771_, _07075_);
  and (_12890_, _12889_, _12888_);
  or (_12891_, _12890_, _06220_);
  or (_12892_, _12876_, _06229_);
  and (_12893_, _12892_, _06153_);
  and (_12894_, _12893_, _12891_);
  or (_12895_, _12894_, _12788_);
  and (_12896_, _12895_, _06146_);
  nand (_12897_, _12784_, _07855_);
  or (_12898_, _12897_, _12774_);
  and (_12899_, _12885_, _06145_);
  and (_12900_, _12899_, _12898_);
  or (_12901_, _12900_, _12896_);
  and (_12902_, _12901_, _06140_);
  or (_12903_, _12785_, _08586_);
  and (_12904_, _12903_, _12773_);
  or (_12905_, _12904_, _12774_);
  and (_12906_, _12905_, _06139_);
  or (_12907_, _12906_, _09842_);
  or (_12908_, _12907_, _12902_);
  and (_12909_, _12908_, _12772_);
  or (_12910_, _12909_, _06116_);
  and (_12911_, _12768_, _08535_);
  or (_12912_, _12769_, _06117_);
  or (_12913_, _12912_, _12911_);
  and (_12914_, _12913_, _06114_);
  and (_12915_, _12914_, _12910_);
  and (_12916_, _08731_, _08703_);
  and (_12917_, _12916_, \oc8051_golden_model_1.P0 [7]);
  and (_12918_, _08717_, _08731_);
  and (_12919_, _12918_, \oc8051_golden_model_1.P1 [7]);
  and (_12920_, _08748_, _08731_);
  and (_12921_, _12920_, \oc8051_golden_model_1.P2 [7]);
  and (_12922_, _08731_, _08745_);
  and (_12923_, _12922_, \oc8051_golden_model_1.P3 [7]);
  or (_12924_, _12923_, _12921_);
  or (_12925_, _12924_, _12919_);
  or (_12926_, _12925_, _12917_);
  or (_12927_, _12926_, _08782_);
  and (_12928_, _12927_, _12768_);
  or (_12929_, _12928_, _12769_);
  and (_12930_, _12929_, _05787_);
  or (_12931_, _12930_, _06110_);
  or (_12932_, _12931_, _12915_);
  and (_12933_, _12768_, _08607_);
  or (_12934_, _12933_, _12769_);
  or (_12935_, _12934_, _06111_);
  and (_12936_, _12935_, _07127_);
  and (_12937_, _12936_, _12932_);
  nand (_12938_, _12801_, _08395_);
  and (_12939_, _12938_, _12768_);
  or (_12940_, _12939_, _12769_);
  or (_12941_, _12801_, _08395_);
  or (_12942_, _12941_, _12769_);
  and (_12943_, _12942_, _06297_);
  and (_12944_, _12943_, _12940_);
  or (_12945_, _12944_, _12937_);
  and (_12946_, _12945_, _07125_);
  nand (_12947_, _12801_, _08430_);
  and (_12948_, _12947_, _12768_);
  or (_12949_, _12948_, _12769_);
  or (_12950_, _12801_, _08430_);
  or (_12951_, _12950_, _12769_);
  and (_12952_, _12951_, _06402_);
  and (_12953_, _12952_, _12949_);
  or (_12954_, _12953_, _12946_);
  and (_12955_, _12954_, _07132_);
  or (_12956_, _12802_, _12769_);
  and (_12957_, _12934_, _06306_);
  and (_12958_, _12957_, _12956_);
  or (_12959_, _12958_, _12955_);
  and (_12960_, _12959_, _07130_);
  and (_12961_, _12876_, _06411_);
  and (_12962_, _12961_, _12956_);
  or (_12963_, _12962_, _06303_);
  or (_12964_, _12963_, _12960_);
  or (_12965_, _12940_, _08819_);
  and (_12966_, _12965_, _08824_);
  and (_12967_, _12966_, _12964_);
  and (_12968_, _12949_, _06396_);
  or (_12969_, _12968_, _06433_);
  or (_12970_, _12969_, _12967_);
  or (_12971_, _12873_, _06829_);
  and (_12972_, _12971_, _05749_);
  and (_12973_, _12972_, _12970_);
  and (_12974_, _12787_, _05748_);
  or (_12975_, _12974_, _06440_);
  or (_12976_, _12975_, _12973_);
  and (_12977_, _12858_, _12850_);
  and (_12978_, _12977_, _12842_);
  and (_12979_, _12978_, _12834_);
  and (_12980_, _12979_, _12826_);
  and (_12981_, _12980_, _12818_);
  nand (_12982_, _12981_, _12810_);
  nand (_12983_, _12982_, _12801_);
  or (_12984_, _12982_, _12801_);
  and (_12985_, _12984_, _12983_);
  and (_12986_, _12985_, _12768_);
  or (_12987_, _12769_, _06444_);
  or (_12988_, _12987_, _12986_);
  and (_12989_, _12988_, _01317_);
  and (_12990_, _12989_, _12976_);
  or (_40994_, _12990_, _12765_);
  not (_12991_, _12797_);
  and (_12992_, _12991_, \oc8051_golden_model_1.P3 [7]);
  and (_12993_, _12797_, _07923_);
  or (_12994_, _12993_, _12992_);
  or (_12995_, _12994_, _06132_);
  not (_12996_, _12780_);
  and (_12997_, _12996_, \oc8051_golden_model_1.P3 [7]);
  and (_12998_, _12785_, _12780_);
  or (_12999_, _12998_, _12997_);
  and (_13000_, _12999_, _06152_);
  and (_13001_, _12871_, _12797_);
  or (_13002_, _13001_, _12992_);
  or (_13003_, _13002_, _06161_);
  and (_13004_, _12797_, \oc8051_golden_model_1.ACC [7]);
  or (_13005_, _13004_, _12992_);
  and (_13006_, _13005_, _07056_);
  and (_13007_, _07057_, \oc8051_golden_model_1.P3 [7]);
  or (_13008_, _13007_, _06160_);
  or (_13009_, _13008_, _13006_);
  and (_13010_, _13009_, _06157_);
  and (_13011_, _13010_, _13003_);
  and (_13012_, _12883_, _12780_);
  or (_13013_, _13012_, _12997_);
  and (_13014_, _13013_, _06156_);
  or (_13015_, _13014_, _06217_);
  or (_13016_, _13015_, _13011_);
  or (_13017_, _12994_, _07075_);
  and (_13018_, _13017_, _13016_);
  or (_13019_, _13018_, _06220_);
  or (_13020_, _13005_, _06229_);
  and (_13021_, _13020_, _06153_);
  and (_13022_, _13021_, _13019_);
  or (_13023_, _13022_, _13000_);
  and (_13024_, _13023_, _06146_);
  or (_13025_, _12997_, _12897_);
  and (_13026_, _13013_, _06145_);
  and (_13027_, _13026_, _13025_);
  or (_13028_, _13027_, _13024_);
  and (_13029_, _13028_, _06140_);
  and (_13030_, _12903_, _12780_);
  or (_13031_, _13030_, _12997_);
  and (_13032_, _13031_, _06139_);
  or (_13033_, _13032_, _09842_);
  or (_13034_, _13033_, _13029_);
  and (_13035_, _13034_, _12995_);
  or (_13036_, _13035_, _06116_);
  and (_13037_, _12797_, _08535_);
  or (_13038_, _12992_, _06117_);
  or (_13039_, _13038_, _13037_);
  and (_13040_, _13039_, _06114_);
  and (_13041_, _13040_, _13036_);
  and (_13042_, _12927_, _12797_);
  or (_13043_, _13042_, _12992_);
  and (_13044_, _13043_, _05787_);
  or (_13045_, _13044_, _06110_);
  or (_13046_, _13045_, _13041_);
  and (_13047_, _12797_, _08607_);
  or (_13048_, _13047_, _12992_);
  or (_13049_, _13048_, _06111_);
  and (_13050_, _13049_, _07127_);
  and (_13051_, _13050_, _13046_);
  and (_13052_, _12938_, _12797_);
  or (_13053_, _13052_, _12992_);
  or (_13054_, _12992_, _12941_);
  and (_13055_, _13054_, _06297_);
  and (_13056_, _13055_, _13053_);
  or (_13057_, _13056_, _13051_);
  and (_13058_, _13057_, _07125_);
  and (_13059_, _12947_, _12797_);
  or (_13060_, _13059_, _12992_);
  or (_13061_, _12992_, _12950_);
  and (_13062_, _13061_, _06402_);
  and (_13063_, _13062_, _13060_);
  or (_13064_, _13063_, _13058_);
  and (_13065_, _13064_, _07132_);
  or (_13066_, _12992_, _12802_);
  and (_13067_, _13048_, _06306_);
  and (_13068_, _13067_, _13066_);
  or (_13069_, _13068_, _13065_);
  and (_13070_, _13069_, _07130_);
  and (_13071_, _13005_, _06411_);
  and (_13072_, _13071_, _13066_);
  or (_13073_, _13072_, _06303_);
  or (_13074_, _13073_, _13070_);
  or (_13075_, _13053_, _08819_);
  and (_13076_, _13075_, _08824_);
  and (_13077_, _13076_, _13074_);
  and (_13078_, _13060_, _06396_);
  or (_13079_, _13078_, _06433_);
  or (_13080_, _13079_, _13077_);
  or (_13081_, _13002_, _06829_);
  and (_13082_, _13081_, _05749_);
  and (_13083_, _13082_, _13080_);
  and (_13084_, _12999_, _05748_);
  or (_13085_, _13084_, _06440_);
  or (_13086_, _13085_, _13083_);
  and (_13087_, _12985_, _12797_);
  or (_13088_, _12992_, _06444_);
  or (_13089_, _13088_, _13087_);
  and (_13090_, _13089_, _01317_);
  and (_13091_, _13090_, _13086_);
  nor (_13092_, \oc8051_golden_model_1.P3 [7], rst);
  nor (_13093_, _13092_, _00000_);
  or (_40995_, _13093_, _13091_);
  nor (_13094_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_13095_, _13094_, _00000_);
  not (_13096_, _12789_);
  and (_13097_, _13096_, \oc8051_golden_model_1.P0 [7]);
  and (_13098_, _12789_, _07923_);
  or (_13099_, _13098_, _13097_);
  or (_13100_, _13099_, _06132_);
  not (_13101_, _07847_);
  and (_13102_, _13101_, \oc8051_golden_model_1.P0 [7]);
  and (_13103_, _12785_, _07847_);
  or (_13104_, _13103_, _13102_);
  and (_13105_, _13104_, _06152_);
  and (_13106_, _12871_, _12789_);
  or (_13107_, _13106_, _13097_);
  or (_13108_, _13107_, _06161_);
  and (_13109_, _12789_, \oc8051_golden_model_1.ACC [7]);
  or (_13110_, _13109_, _13097_);
  and (_13111_, _13110_, _07056_);
  and (_13112_, _07057_, \oc8051_golden_model_1.P0 [7]);
  or (_13113_, _13112_, _06160_);
  or (_13114_, _13113_, _13111_);
  and (_13115_, _13114_, _06157_);
  and (_13116_, _13115_, _13108_);
  and (_13117_, _12883_, _07847_);
  or (_13118_, _13117_, _13102_);
  and (_13119_, _13118_, _06156_);
  or (_13120_, _13119_, _06217_);
  or (_13121_, _13120_, _13116_);
  or (_13122_, _13099_, _07075_);
  and (_13123_, _13122_, _13121_);
  or (_13124_, _13123_, _06220_);
  or (_13125_, _13110_, _06229_);
  and (_13126_, _13125_, _06153_);
  and (_13127_, _13126_, _13124_);
  or (_13128_, _13127_, _13105_);
  and (_13129_, _13128_, _06146_);
  or (_13130_, _13102_, _12897_);
  and (_13131_, _13118_, _06145_);
  and (_13132_, _13131_, _13130_);
  or (_13133_, _13132_, _13129_);
  and (_13134_, _13133_, _06140_);
  and (_13135_, _12903_, _07847_);
  or (_13136_, _13135_, _13102_);
  and (_13137_, _13136_, _06139_);
  or (_13138_, _13137_, _09842_);
  or (_13139_, _13138_, _13134_);
  and (_13140_, _13139_, _13100_);
  or (_13141_, _13140_, _06116_);
  and (_13142_, _12789_, _08535_);
  or (_13143_, _13097_, _06117_);
  or (_13144_, _13143_, _13142_);
  and (_13145_, _13144_, _06114_);
  and (_13146_, _13145_, _13141_);
  and (_13147_, _12927_, _12789_);
  or (_13148_, _13147_, _13097_);
  and (_13149_, _13148_, _05787_);
  or (_13150_, _13149_, _11136_);
  or (_13151_, _13150_, _13146_);
  and (_13152_, _12938_, _12789_);
  and (_13153_, _13152_, _12941_);
  or (_13154_, _13097_, _07127_);
  or (_13155_, _13154_, _13153_);
  and (_13156_, _12789_, _08607_);
  or (_13157_, _13156_, _13097_);
  or (_13158_, _13157_, _06111_);
  and (_13159_, _13158_, _07125_);
  and (_13160_, _13159_, _13155_);
  and (_13161_, _13160_, _13151_);
  and (_13162_, _12947_, _12789_);
  and (_13163_, _13162_, _12950_);
  or (_13164_, _13163_, _13097_);
  and (_13165_, _13164_, _06402_);
  or (_13166_, _13165_, _13161_);
  and (_13167_, _13166_, _07132_);
  or (_13168_, _13097_, _12802_);
  and (_13169_, _13157_, _06306_);
  and (_13170_, _13169_, _13168_);
  or (_13171_, _13170_, _13167_);
  and (_13172_, _13171_, _07130_);
  and (_13173_, _13110_, _06411_);
  and (_13174_, _13173_, _13168_);
  or (_13175_, _13174_, _06303_);
  or (_13176_, _13175_, _13172_);
  or (_13177_, _13097_, _08819_);
  or (_13178_, _13177_, _13152_);
  and (_13179_, _13178_, _08824_);
  and (_13180_, _13179_, _13176_);
  or (_13181_, _13162_, _13097_);
  and (_13182_, _13181_, _06396_);
  or (_13183_, _13182_, _06433_);
  or (_13184_, _13183_, _13180_);
  or (_13185_, _13107_, _06829_);
  and (_13186_, _13185_, _05749_);
  and (_13187_, _13186_, _13184_);
  and (_13188_, _13104_, _05748_);
  or (_13189_, _13188_, _06440_);
  or (_13190_, _13189_, _13187_);
  and (_13191_, _12985_, _12789_);
  or (_13192_, _13097_, _06444_);
  or (_13193_, _13192_, _13191_);
  and (_13194_, _13193_, _01317_);
  and (_13195_, _13194_, _13190_);
  or (_40997_, _13195_, _13095_);
  not (_13196_, _12792_);
  and (_13197_, _13196_, \oc8051_golden_model_1.P1 [7]);
  and (_13198_, _12792_, _07923_);
  or (_13199_, _13198_, _13197_);
  or (_13200_, _13199_, _06132_);
  not (_13201_, _12778_);
  and (_13202_, _13201_, \oc8051_golden_model_1.P1 [7]);
  and (_13203_, _12785_, _12778_);
  or (_13204_, _13203_, _13202_);
  and (_13205_, _13204_, _06152_);
  and (_13206_, _12871_, _12792_);
  or (_13207_, _13206_, _13197_);
  or (_13208_, _13207_, _06161_);
  and (_13209_, _12792_, \oc8051_golden_model_1.ACC [7]);
  or (_13210_, _13209_, _13197_);
  and (_13211_, _13210_, _07056_);
  and (_13212_, _07057_, \oc8051_golden_model_1.P1 [7]);
  or (_13213_, _13212_, _06160_);
  or (_13214_, _13213_, _13211_);
  and (_13215_, _13214_, _06157_);
  and (_13216_, _13215_, _13208_);
  and (_13217_, _12883_, _12778_);
  or (_13218_, _13217_, _13202_);
  and (_13219_, _13218_, _06156_);
  or (_13220_, _13219_, _06217_);
  or (_13221_, _13220_, _13216_);
  or (_13222_, _13199_, _07075_);
  and (_13223_, _13222_, _13221_);
  or (_13224_, _13223_, _06220_);
  or (_13225_, _13210_, _06229_);
  and (_13226_, _13225_, _06153_);
  and (_13227_, _13226_, _13224_);
  or (_13228_, _13227_, _13205_);
  and (_13229_, _13228_, _06146_);
  or (_13230_, _13202_, _12897_);
  and (_13231_, _13218_, _06145_);
  and (_13232_, _13231_, _13230_);
  or (_13233_, _13232_, _13229_);
  and (_13234_, _13233_, _06140_);
  and (_13235_, _12903_, _12778_);
  or (_13236_, _13235_, _13202_);
  and (_13237_, _13236_, _06139_);
  or (_13238_, _13237_, _09842_);
  or (_13239_, _13238_, _13234_);
  and (_13240_, _13239_, _13200_);
  or (_13241_, _13240_, _06116_);
  and (_13242_, _12792_, _08535_);
  or (_13243_, _13197_, _06117_);
  or (_13244_, _13243_, _13242_);
  and (_13245_, _13244_, _06114_);
  and (_13246_, _13245_, _13241_);
  and (_13247_, _12927_, _12792_);
  or (_13248_, _13247_, _13197_);
  and (_13249_, _13248_, _05787_);
  or (_13250_, _13249_, _06110_);
  or (_13251_, _13250_, _13246_);
  and (_13252_, _12792_, _08607_);
  or (_13253_, _13252_, _13197_);
  or (_13254_, _13253_, _06111_);
  and (_13255_, _13254_, _07127_);
  and (_13256_, _13255_, _13251_);
  and (_13257_, _12938_, _12792_);
  or (_13258_, _13257_, _13197_);
  or (_13259_, _13197_, _12941_);
  and (_13260_, _13259_, _06297_);
  and (_13261_, _13260_, _13258_);
  or (_13262_, _13261_, _13256_);
  and (_13263_, _13262_, _07125_);
  and (_13264_, _12947_, _12792_);
  or (_13265_, _13264_, _13197_);
  or (_13266_, _13197_, _12950_);
  and (_13267_, _13266_, _06402_);
  and (_13268_, _13267_, _13265_);
  or (_13269_, _13268_, _13263_);
  and (_13270_, _13269_, _07132_);
  or (_13271_, _13197_, _12802_);
  and (_13272_, _13253_, _06306_);
  and (_13273_, _13272_, _13271_);
  or (_13274_, _13273_, _13270_);
  and (_13275_, _13274_, _07130_);
  and (_13276_, _13210_, _06411_);
  and (_13277_, _13276_, _13271_);
  or (_13278_, _13277_, _06303_);
  or (_13279_, _13278_, _13275_);
  or (_13280_, _13258_, _08819_);
  and (_13281_, _13280_, _08824_);
  and (_13282_, _13281_, _13279_);
  and (_13283_, _13265_, _06396_);
  or (_13284_, _13283_, _06433_);
  or (_13285_, _13284_, _13282_);
  or (_13286_, _13207_, _06829_);
  and (_13287_, _13286_, _05749_);
  and (_13288_, _13287_, _13285_);
  and (_13289_, _13204_, _05748_);
  or (_13290_, _13289_, _06440_);
  or (_13291_, _13290_, _13288_);
  and (_13292_, _12985_, _12792_);
  or (_13293_, _13197_, _06444_);
  or (_13294_, _13293_, _13292_);
  and (_13295_, _13294_, _01317_);
  and (_13296_, _13295_, _13291_);
  nor (_13297_, \oc8051_golden_model_1.P1 [7], rst);
  nor (_13298_, _13297_, _00000_);
  or (_40998_, _13298_, _13296_);
  and (_13299_, _01321_, \oc8051_golden_model_1.IP [7]);
  not (_13300_, _07830_);
  and (_13301_, _13300_, \oc8051_golden_model_1.IP [7]);
  and (_13302_, _07923_, _07830_);
  or (_13303_, _13302_, _13301_);
  or (_13304_, _13303_, _06132_);
  not (_13305_, _08415_);
  and (_13306_, _13305_, \oc8051_golden_model_1.IP [7]);
  and (_13307_, _08426_, _08415_);
  or (_13308_, _13307_, _13306_);
  and (_13309_, _13308_, _06152_);
  and (_13310_, _08548_, _07830_);
  or (_13311_, _13310_, _13301_);
  or (_13312_, _13311_, _06161_);
  and (_13313_, _07830_, \oc8051_golden_model_1.ACC [7]);
  or (_13314_, _13313_, _13301_);
  and (_13315_, _13314_, _07056_);
  and (_13316_, _07057_, \oc8051_golden_model_1.IP [7]);
  or (_13317_, _13316_, _06160_);
  or (_13318_, _13317_, _13315_);
  and (_13319_, _13318_, _06157_);
  and (_13320_, _13319_, _13312_);
  and (_13321_, _08552_, _08415_);
  or (_13322_, _13321_, _13306_);
  and (_13323_, _13322_, _06156_);
  or (_13324_, _13323_, _06217_);
  or (_13325_, _13324_, _13320_);
  or (_13326_, _13303_, _07075_);
  and (_13327_, _13326_, _13325_);
  or (_13328_, _13327_, _06220_);
  or (_13329_, _13314_, _06229_);
  and (_13330_, _13329_, _06153_);
  and (_13331_, _13330_, _13328_);
  or (_13332_, _13331_, _13309_);
  and (_13333_, _13332_, _06146_);
  and (_13334_, _08569_, _08415_);
  or (_13335_, _13334_, _13306_);
  and (_13336_, _13335_, _06145_);
  or (_13337_, _13336_, _13333_);
  and (_13338_, _13337_, _06140_);
  and (_13339_, _08587_, _08415_);
  or (_13340_, _13339_, _13306_);
  and (_13341_, _13340_, _06139_);
  or (_13342_, _13341_, _09842_);
  or (_13343_, _13342_, _13338_);
  and (_13344_, _13343_, _13304_);
  or (_13345_, _13344_, _06116_);
  and (_13346_, _08535_, _07830_);
  or (_13347_, _13301_, _06117_);
  or (_13348_, _13347_, _13346_);
  and (_13349_, _13348_, _06114_);
  and (_13350_, _13349_, _13345_);
  and (_13351_, _08782_, _07830_);
  or (_13352_, _13351_, _13301_);
  and (_13353_, _13352_, _05787_);
  or (_13354_, _13353_, _11136_);
  or (_13355_, _13354_, _13350_);
  and (_13356_, _08802_, _07830_);
  or (_13357_, _13301_, _07127_);
  or (_13358_, _13357_, _13356_);
  and (_13359_, _08607_, _07830_);
  or (_13360_, _13359_, _13301_);
  or (_13361_, _13360_, _06111_);
  and (_13362_, _13361_, _07125_);
  and (_13363_, _13362_, _13358_);
  and (_13364_, _13363_, _13355_);
  and (_13365_, _08810_, _07830_);
  or (_13366_, _13365_, _13301_);
  and (_13367_, _13366_, _06402_);
  or (_13368_, _13367_, _13364_);
  and (_13369_, _13368_, _07132_);
  or (_13370_, _13301_, _07926_);
  and (_13371_, _13360_, _06306_);
  and (_13372_, _13371_, _13370_);
  or (_13373_, _13372_, _13369_);
  and (_13374_, _13373_, _07130_);
  and (_13375_, _13314_, _06411_);
  and (_13376_, _13375_, _13370_);
  or (_13377_, _13376_, _06303_);
  or (_13378_, _13377_, _13374_);
  and (_13379_, _08801_, _07830_);
  or (_13380_, _13301_, _08819_);
  or (_13381_, _13380_, _13379_);
  and (_13382_, _13381_, _08824_);
  and (_13383_, _13382_, _13378_);
  nor (_13384_, _08809_, _13300_);
  or (_13385_, _13384_, _13301_);
  and (_13386_, _13385_, _06396_);
  or (_13387_, _13386_, _06433_);
  or (_13388_, _13387_, _13383_);
  or (_13389_, _13311_, _06829_);
  and (_13390_, _13389_, _05749_);
  and (_13391_, _13390_, _13388_);
  and (_13392_, _13308_, _05748_);
  or (_13393_, _13392_, _06440_);
  or (_13394_, _13393_, _13391_);
  and (_13395_, _08345_, _07830_);
  or (_13396_, _13301_, _06444_);
  or (_13397_, _13396_, _13395_);
  and (_13398_, _13397_, _01317_);
  and (_13399_, _13398_, _13394_);
  or (_13400_, _13399_, _13299_);
  and (_40999_, _13400_, _43100_);
  and (_13401_, _01321_, \oc8051_golden_model_1.IE [7]);
  not (_13402_, _07826_);
  and (_13403_, _13402_, \oc8051_golden_model_1.IE [7]);
  and (_13404_, _07923_, _07826_);
  or (_13405_, _13404_, _13403_);
  or (_13406_, _13405_, _06132_);
  not (_13407_, _08418_);
  and (_13408_, _13407_, \oc8051_golden_model_1.IE [7]);
  and (_13409_, _08426_, _08418_);
  or (_13410_, _13409_, _13408_);
  and (_13411_, _13410_, _06152_);
  and (_13412_, _08548_, _07826_);
  or (_13413_, _13412_, _13403_);
  or (_13414_, _13413_, _06161_);
  and (_13415_, _07826_, \oc8051_golden_model_1.ACC [7]);
  or (_13416_, _13415_, _13403_);
  and (_13417_, _13416_, _07056_);
  and (_13418_, _07057_, \oc8051_golden_model_1.IE [7]);
  or (_13419_, _13418_, _06160_);
  or (_13420_, _13419_, _13417_);
  and (_13421_, _13420_, _06157_);
  and (_13422_, _13421_, _13414_);
  and (_13423_, _08552_, _08418_);
  or (_13424_, _13423_, _13408_);
  and (_13425_, _13424_, _06156_);
  or (_13426_, _13425_, _06217_);
  or (_13427_, _13426_, _13422_);
  or (_13428_, _13405_, _07075_);
  and (_13429_, _13428_, _13427_);
  or (_13430_, _13429_, _06220_);
  or (_13431_, _13416_, _06229_);
  and (_13432_, _13431_, _06153_);
  and (_13433_, _13432_, _13430_);
  or (_13434_, _13433_, _13411_);
  and (_13435_, _13434_, _06146_);
  and (_13436_, _08569_, _08418_);
  or (_13437_, _13436_, _13408_);
  and (_13438_, _13437_, _06145_);
  or (_13439_, _13438_, _13435_);
  and (_13440_, _13439_, _06140_);
  and (_13441_, _08587_, _08418_);
  or (_13442_, _13441_, _13408_);
  and (_13443_, _13442_, _06139_);
  or (_13444_, _13443_, _09842_);
  or (_13445_, _13444_, _13440_);
  and (_13446_, _13445_, _13406_);
  or (_13447_, _13446_, _06116_);
  and (_13448_, _08535_, _07826_);
  or (_13449_, _13403_, _06117_);
  or (_13450_, _13449_, _13448_);
  and (_13451_, _13450_, _06114_);
  and (_13452_, _13451_, _13447_);
  and (_13453_, _08782_, _07826_);
  or (_13454_, _13453_, _13403_);
  and (_13455_, _13454_, _05787_);
  or (_13456_, _13455_, _11136_);
  or (_13457_, _13456_, _13452_);
  and (_13458_, _08802_, _07826_);
  or (_13459_, _13403_, _07127_);
  or (_13460_, _13459_, _13458_);
  and (_13461_, _08607_, _07826_);
  or (_13462_, _13461_, _13403_);
  or (_13463_, _13462_, _06111_);
  and (_13464_, _13463_, _07125_);
  and (_13465_, _13464_, _13460_);
  and (_13466_, _13465_, _13457_);
  and (_13467_, _08810_, _07826_);
  or (_13468_, _13467_, _13403_);
  and (_13469_, _13468_, _06402_);
  or (_13470_, _13469_, _13466_);
  and (_13471_, _13470_, _07132_);
  or (_13472_, _13403_, _07926_);
  and (_13473_, _13462_, _06306_);
  and (_13474_, _13473_, _13472_);
  or (_13475_, _13474_, _13471_);
  and (_13476_, _13475_, _07130_);
  and (_13477_, _13416_, _06411_);
  and (_13478_, _13477_, _13472_);
  or (_13479_, _13478_, _06303_);
  or (_13480_, _13479_, _13476_);
  and (_13481_, _08801_, _07826_);
  or (_13482_, _13403_, _08819_);
  or (_13483_, _13482_, _13481_);
  and (_13484_, _13483_, _08824_);
  and (_13485_, _13484_, _13480_);
  nor (_13486_, _08809_, _13402_);
  or (_13487_, _13486_, _13403_);
  and (_13488_, _13487_, _06396_);
  or (_13489_, _13488_, _06433_);
  or (_13490_, _13489_, _13485_);
  or (_13491_, _13413_, _06829_);
  and (_13492_, _13491_, _05749_);
  and (_13493_, _13492_, _13490_);
  and (_13494_, _13410_, _05748_);
  or (_13495_, _13494_, _06440_);
  or (_13496_, _13495_, _13493_);
  and (_13497_, _08345_, _07826_);
  or (_13498_, _13403_, _06444_);
  or (_13499_, _13498_, _13497_);
  and (_13500_, _13499_, _01317_);
  and (_13501_, _13500_, _13496_);
  or (_13502_, _13501_, _13401_);
  and (_41000_, _13502_, _43100_);
  and (_13503_, _01321_, \oc8051_golden_model_1.SCON [7]);
  not (_13504_, _07778_);
  and (_13505_, _13504_, \oc8051_golden_model_1.SCON [7]);
  and (_13506_, _07923_, _07778_);
  or (_13507_, _13506_, _13505_);
  or (_13508_, _13507_, _06132_);
  not (_13509_, _08413_);
  and (_13510_, _13509_, \oc8051_golden_model_1.SCON [7]);
  and (_13511_, _08426_, _08413_);
  or (_13512_, _13511_, _13510_);
  and (_13513_, _13512_, _06152_);
  and (_13514_, _08548_, _07778_);
  or (_13515_, _13514_, _13505_);
  or (_13516_, _13515_, _06161_);
  and (_13517_, _07778_, \oc8051_golden_model_1.ACC [7]);
  or (_13518_, _13517_, _13505_);
  and (_13519_, _13518_, _07056_);
  and (_13520_, _07057_, \oc8051_golden_model_1.SCON [7]);
  or (_13521_, _13520_, _06160_);
  or (_13522_, _13521_, _13519_);
  and (_13523_, _13522_, _06157_);
  and (_13524_, _13523_, _13516_);
  and (_13525_, _08552_, _08413_);
  or (_13526_, _13525_, _13510_);
  and (_13527_, _13526_, _06156_);
  or (_13528_, _13527_, _06217_);
  or (_13529_, _13528_, _13524_);
  or (_13530_, _13507_, _07075_);
  and (_13531_, _13530_, _13529_);
  or (_13532_, _13531_, _06220_);
  or (_13533_, _13518_, _06229_);
  and (_13534_, _13533_, _06153_);
  and (_13535_, _13534_, _13532_);
  or (_13536_, _13535_, _13513_);
  and (_13537_, _13536_, _06146_);
  and (_13538_, _08569_, _08413_);
  or (_13539_, _13538_, _13510_);
  and (_13540_, _13539_, _06145_);
  or (_13541_, _13540_, _13537_);
  and (_13542_, _13541_, _06140_);
  and (_13543_, _08587_, _08413_);
  or (_13544_, _13543_, _13510_);
  and (_13545_, _13544_, _06139_);
  or (_13546_, _13545_, _09842_);
  or (_13547_, _13546_, _13542_);
  and (_13548_, _13547_, _13508_);
  or (_13549_, _13548_, _06116_);
  and (_13550_, _08535_, _07778_);
  or (_13551_, _13505_, _06117_);
  or (_13552_, _13551_, _13550_);
  and (_13553_, _13552_, _06114_);
  and (_13554_, _13553_, _13549_);
  and (_13555_, _08782_, _07778_);
  or (_13556_, _13555_, _13505_);
  and (_13557_, _13556_, _05787_);
  or (_13558_, _13557_, _11136_);
  or (_13559_, _13558_, _13554_);
  and (_13560_, _08802_, _07778_);
  or (_13561_, _13505_, _07127_);
  or (_13562_, _13561_, _13560_);
  and (_13563_, _08607_, _07778_);
  or (_13564_, _13563_, _13505_);
  or (_13565_, _13564_, _06111_);
  and (_13566_, _13565_, _07125_);
  and (_13567_, _13566_, _13562_);
  and (_13568_, _13567_, _13559_);
  and (_13569_, _08810_, _07778_);
  or (_13570_, _13569_, _13505_);
  and (_13571_, _13570_, _06402_);
  or (_13572_, _13571_, _13568_);
  and (_13573_, _13572_, _07132_);
  or (_13574_, _13505_, _07926_);
  and (_13575_, _13564_, _06306_);
  and (_13576_, _13575_, _13574_);
  or (_13577_, _13576_, _13573_);
  and (_13578_, _13577_, _07130_);
  and (_13579_, _13518_, _06411_);
  and (_13580_, _13579_, _13574_);
  or (_13581_, _13580_, _06303_);
  or (_13582_, _13581_, _13578_);
  and (_13583_, _08801_, _07778_);
  or (_13584_, _13505_, _08819_);
  or (_13585_, _13584_, _13583_);
  and (_13586_, _13585_, _08824_);
  and (_13587_, _13586_, _13582_);
  nor (_13588_, _08809_, _13504_);
  or (_13589_, _13588_, _13505_);
  and (_13590_, _13589_, _06396_);
  or (_13591_, _13590_, _06433_);
  or (_13592_, _13591_, _13587_);
  or (_13593_, _13515_, _06829_);
  and (_13594_, _13593_, _05749_);
  and (_13595_, _13594_, _13592_);
  and (_13596_, _13512_, _05748_);
  or (_13597_, _13596_, _06440_);
  or (_13598_, _13597_, _13595_);
  and (_13599_, _08345_, _07778_);
  or (_13600_, _13505_, _06444_);
  or (_13601_, _13600_, _13599_);
  and (_13602_, _13601_, _01317_);
  and (_13603_, _13602_, _13598_);
  or (_13604_, _13603_, _13503_);
  and (_41001_, _13604_, _43100_);
  not (_13605_, \oc8051_golden_model_1.SP [7]);
  nor (_13606_, _01317_, _13605_);
  and (_13607_, _07756_, \oc8051_golden_model_1.SP [4]);
  and (_13608_, _13607_, \oc8051_golden_model_1.SP [5]);
  and (_13609_, _13608_, \oc8051_golden_model_1.SP [6]);
  or (_13610_, _13609_, \oc8051_golden_model_1.SP [7]);
  nand (_13611_, _13609_, \oc8051_golden_model_1.SP [7]);
  and (_13612_, _13611_, _13610_);
  or (_13613_, _13612_, _07160_);
  nor (_13614_, _11388_, _07814_);
  and (_13615_, _13614_, _07787_);
  nor (_13616_, _13615_, _13605_);
  and (_13617_, _08810_, _07858_);
  or (_13618_, _13617_, _13616_);
  and (_13619_, _13618_, _06402_);
  not (_13620_, _06133_);
  and (_13621_, _07923_, _07858_);
  or (_13622_, _13616_, _06116_);
  or (_13623_, _13622_, _13621_);
  and (_13624_, _13623_, _13620_);
  and (_13625_, _08548_, _07858_);
  or (_13626_, _13625_, _13616_);
  or (_13627_, _13626_, _06161_);
  and (_13628_, _13615_, \oc8051_golden_model_1.ACC [7]);
  or (_13629_, _13628_, _13616_);
  or (_13630_, _13629_, _07057_);
  or (_13631_, _07056_, \oc8051_golden_model_1.SP [7]);
  and (_13632_, _13631_, _06582_);
  and (_13633_, _13632_, _13630_);
  and (_13634_, _13612_, _06581_);
  or (_13635_, _13634_, _06160_);
  or (_13636_, _13635_, _13633_);
  and (_13637_, _13636_, _05764_);
  and (_13638_, _13637_, _13627_);
  and (_13639_, _13612_, _07485_);
  or (_13640_, _13639_, _06217_);
  or (_13641_, _13640_, _13638_);
  not (_13642_, \oc8051_golden_model_1.SP [6]);
  not (_13643_, \oc8051_golden_model_1.SP [5]);
  not (_13644_, \oc8051_golden_model_1.SP [4]);
  and (_13645_, _08453_, _13644_);
  and (_13646_, _13645_, _13643_);
  and (_13647_, _13646_, _13642_);
  and (_13648_, _13647_, _06142_);
  nor (_13650_, _13648_, _13605_);
  and (_13651_, _13648_, _13605_);
  nor (_13652_, _13651_, _13650_);
  nand (_13653_, _13652_, _06217_);
  and (_13654_, _13653_, _13641_);
  or (_13655_, _13654_, _06220_);
  or (_13656_, _13629_, _06229_);
  and (_13657_, _13656_, _07191_);
  and (_13658_, _13657_, _13655_);
  and (_13659_, _13608_, \oc8051_golden_model_1.SP [0]);
  and (_13661_, _13659_, \oc8051_golden_model_1.SP [6]);
  nor (_13662_, _13661_, _13605_);
  and (_13663_, _13661_, _13605_);
  or (_13664_, _13663_, _13662_);
  nand (_13665_, _13664_, _06151_);
  nand (_13666_, _13665_, _07389_);
  or (_13667_, _13666_, _13658_);
  or (_13668_, _13612_, _07389_);
  and (_13669_, _13668_, _06132_);
  and (_13670_, _13669_, _13667_);
  or (_13672_, _13670_, _13624_);
  or (_13673_, _13616_, _06117_);
  and (_13674_, _08535_, _13615_);
  or (_13675_, _13674_, _13673_);
  and (_13676_, _13675_, _06114_);
  and (_13677_, _13676_, _13672_);
  and (_13678_, _08782_, _07858_);
  or (_13679_, _13678_, _13616_);
  and (_13680_, _13679_, _05787_);
  or (_13681_, _13680_, _06110_);
  or (_13683_, _13681_, _13677_);
  and (_13684_, _08607_, _13615_);
  or (_13685_, _13684_, _13616_);
  or (_13686_, _13685_, _06111_);
  and (_13687_, _13686_, _13683_);
  or (_13688_, _13687_, _06076_);
  or (_13689_, _13612_, _05836_);
  and (_13690_, _13689_, _13688_);
  or (_13691_, _13690_, _06297_);
  and (_13692_, _08802_, _13615_);
  or (_13694_, _13692_, _13616_);
  or (_13695_, _13694_, _07127_);
  and (_13696_, _13695_, _07125_);
  and (_13697_, _13696_, _13691_);
  or (_13698_, _13697_, _13619_);
  and (_13699_, _13698_, _07132_);
  or (_13700_, _13616_, _07926_);
  and (_13701_, _13685_, _06306_);
  and (_13702_, _13701_, _13700_);
  or (_13703_, _13702_, _13699_);
  and (_13705_, _13703_, _12514_);
  and (_13706_, _13629_, _06411_);
  and (_13707_, _13706_, _13700_);
  and (_13708_, _13612_, _07124_);
  or (_13709_, _13708_, _06303_);
  or (_13710_, _13709_, _13707_);
  or (_13711_, _13710_, _13705_);
  and (_13712_, _08801_, _07858_);
  or (_13713_, _13616_, _08819_);
  or (_13714_, _13713_, _13712_);
  and (_13716_, _13714_, _13711_);
  or (_13717_, _13716_, _06396_);
  not (_13718_, _07858_);
  nor (_13719_, _08809_, _13718_);
  or (_13720_, _13616_, _08824_);
  or (_13721_, _13720_, _13719_);
  and (_13722_, _13721_, _12558_);
  and (_13723_, _13722_, _13717_);
  or (_13724_, _13647_, \oc8051_golden_model_1.SP [7]);
  nand (_13725_, _13647_, \oc8051_golden_model_1.SP [7]);
  and (_13727_, _13725_, _13724_);
  and (_13728_, _13727_, _06417_);
  or (_13729_, _13728_, _07142_);
  or (_13730_, _13729_, _13723_);
  or (_13731_, _13612_, _05846_);
  and (_13732_, _13731_, _13730_);
  or (_13733_, _13732_, _06167_);
  or (_13734_, _13727_, _06168_);
  and (_13735_, _13734_, _06829_);
  and (_13736_, _13735_, _13733_);
  and (_13738_, _13626_, _06433_);
  or (_13739_, _13738_, _07577_);
  or (_13740_, _13739_, _13736_);
  and (_13741_, _13740_, _13613_);
  or (_13742_, _13741_, _06440_);
  and (_13743_, _08345_, _07858_);
  or (_13744_, _13616_, _06444_);
  or (_13745_, _13744_, _13743_);
  and (_13746_, _13745_, _01317_);
  and (_13747_, _13746_, _13742_);
  or (_13749_, _13747_, _13606_);
  and (_41003_, _13749_, _43100_);
  not (_13750_, _07783_);
  and (_13751_, _13750_, \oc8051_golden_model_1.SBUF [7]);
  and (_13752_, _08548_, _07783_);
  or (_13753_, _13752_, _13751_);
  or (_13754_, _13753_, _06161_);
  and (_13755_, _07783_, \oc8051_golden_model_1.ACC [7]);
  or (_13756_, _13755_, _13751_);
  and (_13757_, _13756_, _07056_);
  and (_13759_, _07057_, \oc8051_golden_model_1.SBUF [7]);
  or (_13760_, _13759_, _06160_);
  or (_13761_, _13760_, _13757_);
  and (_13762_, _13761_, _07075_);
  and (_13763_, _13762_, _13754_);
  and (_13764_, _07923_, _07783_);
  or (_13765_, _13764_, _13751_);
  and (_13766_, _13765_, _06217_);
  or (_13767_, _13766_, _13763_);
  and (_13768_, _13767_, _06229_);
  and (_13770_, _13756_, _06220_);
  or (_13771_, _13770_, _09842_);
  or (_13772_, _13771_, _13768_);
  or (_13773_, _13765_, _06132_);
  and (_13774_, _13773_, _13772_);
  or (_13775_, _13774_, _06116_);
  and (_13776_, _08535_, _07783_);
  or (_13777_, _13751_, _06117_);
  or (_13778_, _13777_, _13776_);
  and (_13779_, _13778_, _06114_);
  and (_13781_, _13779_, _13775_);
  and (_13782_, _08782_, _07783_);
  or (_13783_, _13782_, _13751_);
  and (_13784_, _13783_, _05787_);
  or (_13785_, _13784_, _13781_);
  or (_13786_, _13785_, _11136_);
  and (_13787_, _08802_, _07783_);
  or (_13788_, _13751_, _07127_);
  or (_13789_, _13788_, _13787_);
  and (_13790_, _08607_, _07783_);
  or (_13792_, _13790_, _13751_);
  or (_13793_, _13792_, _06111_);
  and (_13794_, _13793_, _07125_);
  and (_13795_, _13794_, _13789_);
  and (_13796_, _13795_, _13786_);
  and (_13797_, _08810_, _07783_);
  or (_13798_, _13797_, _13751_);
  and (_13799_, _13798_, _06402_);
  or (_13800_, _13799_, _13796_);
  and (_13801_, _13800_, _07132_);
  or (_13802_, _13751_, _07926_);
  and (_13803_, _13792_, _06306_);
  and (_13804_, _13803_, _13802_);
  or (_13805_, _13804_, _13801_);
  and (_13806_, _13805_, _07130_);
  and (_13807_, _13756_, _06411_);
  and (_13808_, _13807_, _13802_);
  or (_13809_, _13808_, _06303_);
  or (_13810_, _13809_, _13806_);
  and (_13811_, _08801_, _07783_);
  or (_13812_, _13751_, _08819_);
  or (_13813_, _13812_, _13811_);
  and (_13814_, _13813_, _08824_);
  and (_13815_, _13814_, _13810_);
  nor (_13816_, _08809_, _13750_);
  or (_13817_, _13816_, _13751_);
  and (_13818_, _13817_, _06396_);
  or (_13819_, _13818_, _06433_);
  or (_13820_, _13819_, _13815_);
  or (_13821_, _13753_, _06829_);
  and (_13822_, _13821_, _06444_);
  and (_13823_, _13822_, _13820_);
  and (_13824_, _08345_, _07783_);
  or (_13825_, _13824_, _13751_);
  and (_13826_, _13825_, _06440_);
  or (_13827_, _13826_, _01321_);
  or (_13828_, _13827_, _13823_);
  or (_13829_, _01317_, \oc8051_golden_model_1.SBUF [7]);
  and (_13830_, _13829_, _43100_);
  and (_41004_, _13830_, _13828_);
  nor (_13831_, _01317_, _10693_);
  and (_13832_, _11094_, \oc8051_golden_model_1.ACC [0]);
  nor (_13833_, _07794_, _10693_);
  and (_13834_, _08810_, _07794_);
  or (_13835_, _13834_, _13833_);
  and (_13836_, _13835_, _06402_);
  and (_13837_, _08782_, _07794_);
  or (_13838_, _13837_, _13833_);
  and (_13839_, _13838_, _05787_);
  and (_13840_, _07923_, _07794_);
  or (_13841_, _13840_, _13833_);
  or (_13842_, _13841_, _06132_);
  not (_13843_, _06254_);
  not (_13844_, _06255_);
  nor (_13845_, _12682_, _13844_);
  nor (_13846_, _09295_, _06255_);
  and (_13847_, _08548_, _07794_);
  or (_13848_, _13847_, _13833_);
  or (_13849_, _13848_, _06161_);
  and (_13850_, _07794_, \oc8051_golden_model_1.ACC [7]);
  or (_13851_, _13850_, _13833_);
  and (_13852_, _13851_, _07056_);
  nor (_13853_, _07056_, _10693_);
  or (_13854_, _13853_, _06160_);
  or (_13855_, _13854_, _13852_);
  and (_13856_, _13855_, _10491_);
  and (_13857_, _13856_, _13849_);
  nor (_13858_, _10508_, _10507_);
  nor (_13859_, _13858_, _10491_);
  not (_13860_, _06221_);
  or (_13861_, _12133_, _13860_);
  or (_13862_, _13861_, _13859_);
  or (_13863_, _13862_, _13857_);
  nor (_13864_, _08404_, _10693_);
  and (_13865_, _08552_, _08404_);
  or (_13866_, _13865_, _13864_);
  or (_13867_, _13866_, _06157_);
  or (_13868_, _13841_, _07075_);
  and (_13869_, _13868_, _13867_);
  and (_13870_, _13869_, _13863_);
  or (_13871_, _13870_, _06220_);
  or (_13872_, _13851_, _06229_);
  nor (_13873_, _12299_, _06152_);
  and (_13874_, _13873_, _13872_);
  and (_13875_, _13874_, _13871_);
  and (_13876_, _08426_, _08404_);
  or (_13877_, _13876_, _13864_);
  and (_13878_, _13877_, _06152_);
  or (_13879_, _13878_, _12126_);
  or (_13880_, _13879_, _13875_);
  and (_13881_, _12108_, _12109_);
  or (_13882_, _13881_, _12106_);
  and (_13883_, _12113_, _12112_);
  or (_13884_, _13883_, _13882_);
  and (_13885_, _13884_, _12105_);
  not (_13886_, _12101_);
  nand (_13887_, _13886_, _12098_);
  and (_13888_, _13887_, _12094_);
  nor (_13889_, _13888_, _07924_);
  or (_13890_, _13889_, _12119_);
  nor (_13891_, _13890_, _13885_);
  nor (_13892_, _13891_, _12120_);
  or (_13893_, _13892_, _12125_);
  and (_13894_, _13893_, _12089_);
  and (_13895_, _13894_, _13880_);
  not (_13896_, _11929_);
  nand (_13897_, _11927_, _13896_);
  nand (_13898_, _13897_, _11926_);
  not (_13899_, _11934_);
  or (_13900_, _11938_, _13899_);
  and (_13901_, _13900_, _11932_);
  or (_13902_, _13901_, _13898_);
  and (_13903_, _13902_, _11954_);
  nor (_13904_, _11943_, _08581_);
  nand (_13905_, _11951_, _11948_);
  and (_13906_, _11946_, _13905_);
  and (_13907_, _13906_, _11947_);
  or (_13908_, _13907_, _11941_);
  or (_13909_, _13908_, _13904_);
  or (_13910_, _13909_, _13903_);
  and (_13911_, _11956_, _06687_);
  and (_13912_, _13911_, _13910_);
  or (_13913_, _13912_, _13895_);
  and (_13914_, _13913_, _06643_);
  nand (_13915_, _08139_, \oc8051_golden_model_1.ACC [3]);
  nor (_13916_, _08247_, \oc8051_golden_model_1.ACC [2]);
  nor (_13917_, _08139_, \oc8051_golden_model_1.ACC [3]);
  or (_13918_, _13917_, _13916_);
  and (_13919_, _13918_, _13915_);
  nor (_13920_, _08175_, \oc8051_golden_model_1.ACC [1]);
  nor (_13921_, _08211_, _05855_);
  nor (_13922_, _13921_, _10278_);
  or (_13923_, _13922_, _13920_);
  and (_13924_, _13923_, _12319_);
  or (_13925_, _13924_, _13919_);
  and (_13926_, _13925_, _12328_);
  nand (_13927_, _08103_, \oc8051_golden_model_1.ACC [5]);
  nor (_13928_, _08338_, \oc8051_golden_model_1.ACC [4]);
  nor (_13929_, _08103_, \oc8051_golden_model_1.ACC [5]);
  or (_13930_, _13929_, _13928_);
  and (_13931_, _13930_, _13927_);
  and (_13932_, _13931_, _12327_);
  nor (_13933_, _07925_, \oc8051_golden_model_1.ACC [7]);
  or (_13934_, _08014_, \oc8051_golden_model_1.ACC [6]);
  nor (_13935_, _13934_, _08810_);
  or (_13936_, _13935_, _13933_);
  or (_13937_, _13936_, _13932_);
  or (_13938_, _13937_, _13926_);
  nor (_13939_, _12329_, _06643_);
  and (_13940_, _13939_, _13938_);
  or (_13941_, _13940_, _13914_);
  and (_13942_, _13941_, _12317_);
  nor (_13943_, _06912_, \oc8051_golden_model_1.ACC [1]);
  and (_13944_, _06912_, \oc8051_golden_model_1.ACC [1]);
  and (_13945_, _06107_, \oc8051_golden_model_1.ACC [0]);
  nor (_13946_, _13945_, _13944_);
  or (_13947_, _13946_, _13943_);
  and (_13948_, _13947_, _12337_);
  nand (_13949_, _06070_, \oc8051_golden_model_1.ACC [3]);
  nor (_13950_, _06070_, \oc8051_golden_model_1.ACC [3]);
  nor (_13951_, _06625_, \oc8051_golden_model_1.ACC [2]);
  or (_13952_, _13951_, _13950_);
  and (_13953_, _13952_, _13949_);
  or (_13954_, _13953_, _13948_);
  and (_13955_, _13954_, _12345_);
  nand (_13956_, _06477_, \oc8051_golden_model_1.ACC [5]);
  nor (_13957_, _06477_, \oc8051_golden_model_1.ACC [5]);
  nor (_13958_, _06876_, \oc8051_golden_model_1.ACC [4]);
  or (_13959_, _13958_, _13957_);
  and (_13960_, _13959_, _13956_);
  and (_13961_, _13960_, _12344_);
  and (_13962_, _06039_, _08430_);
  or (_13963_, _06203_, \oc8051_golden_model_1.ACC [6]);
  nor (_13964_, _13963_, _10794_);
  or (_13965_, _13964_, _13962_);
  or (_13966_, _13965_, _13961_);
  or (_13967_, _13966_, _13955_);
  nor (_13968_, _12346_, _12317_);
  and (_13969_, _13968_, _13967_);
  or (_13970_, _13969_, _11924_);
  or (_13971_, _13970_, _13942_);
  nand (_13972_, _11924_, \oc8051_golden_model_1.PSW [7]);
  and (_13973_, _13972_, _06146_);
  and (_13974_, _13973_, _13971_);
  or (_13975_, _13864_, _08568_);
  and (_13976_, _13975_, _06145_);
  and (_13977_, _13976_, _13866_);
  nor (_13978_, _13977_, _13974_);
  nor (_13979_, _13978_, _06212_);
  and (_13980_, _12682_, \oc8051_golden_model_1.PSW [7]);
  and (_13981_, _13980_, _06212_);
  or (_13982_, _13981_, _13979_);
  and (_13983_, _13982_, _13846_);
  or (_13984_, _13983_, _13845_);
  and (_13985_, _13984_, _13843_);
  or (_13986_, _12682_, \oc8051_golden_model_1.PSW [7]);
  nand (_13987_, _13986_, _06254_);
  nand (_13988_, _13987_, _10553_);
  or (_13989_, _13988_, _13985_);
  and (_13990_, _10302_, _07923_);
  and (_13991_, _10313_, _10308_);
  nor (_13992_, _13991_, _10306_);
  nand (_13993_, _10315_, _10308_);
  or (_13994_, _13993_, _10572_);
  and (_13995_, _13994_, _13992_);
  or (_13996_, _13995_, _13990_);
  and (_13997_, _13996_, _10546_);
  or (_13998_, _13997_, _10554_);
  and (_13999_, _13998_, _13989_);
  and (_14000_, _13996_, _10545_);
  or (_14001_, _14000_, _12379_);
  or (_14002_, _14001_, _13999_);
  and (_14003_, _10593_, _10589_);
  nor (_14004_, _14003_, _10587_);
  nand (_14005_, _10640_, _10589_);
  or (_14006_, _14005_, _10638_);
  and (_14007_, _14006_, _14004_);
  and (_14008_, _10583_, _08535_);
  or (_14009_, _14008_, _12380_);
  or (_14010_, _14009_, _14007_);
  and (_14011_, _14010_, _14002_);
  or (_14012_, _14011_, _06260_);
  and (_14013_, _10405_, _10401_);
  nor (_14014_, _14013_, _10399_);
  nand (_14015_, _10447_, _10401_);
  or (_14016_, _14015_, _10445_);
  and (_14017_, _14016_, _14014_);
  and (_14018_, _10395_, _07926_);
  or (_14019_, _14018_, _06265_);
  or (_14020_, _14019_, _14017_);
  and (_14021_, _14020_, _10388_);
  and (_14022_, _14021_, _14012_);
  and (_14023_, _10665_, _10662_);
  nor (_14024_, _14023_, _10660_);
  nand (_14025_, _10713_, _10662_);
  or (_14026_, _14025_, _10711_);
  and (_14027_, _14026_, _14024_);
  or (_14028_, _14027_, _10655_);
  and (_14029_, _14028_, _10387_);
  or (_14030_, _14029_, _09842_);
  or (_14031_, _14030_, _14022_);
  and (_14032_, _14031_, _13842_);
  or (_14033_, _14032_, _06116_);
  and (_14034_, _08535_, _07794_);
  or (_14035_, _13833_, _06117_);
  or (_14036_, _14035_, _14034_);
  and (_14037_, _14036_, _06114_);
  and (_14038_, _14037_, _14033_);
  or (_14039_, _14038_, _13839_);
  nor (_14040_, _09855_, _06209_);
  and (_14041_, _14040_, _14039_);
  nor (_14042_, _12682_, _10693_);
  and (_14043_, _14042_, _06209_);
  or (_14044_, _14043_, _06110_);
  or (_14045_, _14044_, _14041_);
  and (_14046_, _08607_, _07794_);
  or (_14047_, _14046_, _13833_);
  or (_14048_, _14047_, _06111_);
  and (_14049_, _14048_, _14045_);
  or (_14050_, _14049_, _06208_);
  nand (_14051_, _12682_, _10693_);
  or (_14052_, _14051_, _06768_);
  and (_14053_, _14052_, _14050_);
  or (_14054_, _14053_, _06297_);
  and (_14055_, _08802_, _07794_);
  or (_14056_, _14055_, _13833_);
  or (_14057_, _14056_, _07127_);
  and (_14058_, _14057_, _07125_);
  and (_14059_, _14058_, _14054_);
  or (_14060_, _14059_, _13836_);
  and (_14061_, _14060_, _07132_);
  or (_14062_, _13833_, _07926_);
  and (_14063_, _14047_, _06306_);
  and (_14064_, _14063_, _14062_);
  or (_14065_, _14064_, _14061_);
  and (_14066_, _14065_, _07130_);
  and (_14067_, _13851_, _06411_);
  and (_14068_, _14067_, _14062_);
  or (_14069_, _14068_, _06303_);
  or (_14070_, _14069_, _14066_);
  and (_14071_, _08801_, _07794_);
  or (_14072_, _13833_, _08819_);
  or (_14073_, _14072_, _14071_);
  and (_14074_, _14073_, _08824_);
  and (_14075_, _14074_, _14070_);
  not (_14076_, _07794_);
  nor (_14077_, _08809_, _14076_);
  or (_14078_, _14077_, _13833_);
  and (_14079_, _14078_, _06396_);
  or (_14080_, _14079_, _12547_);
  or (_14081_, _14080_, _14075_);
  nor (_14082_, _10586_, _08430_);
  or (_14083_, _14082_, _10889_);
  or (_14084_, _10867_, _14008_);
  or (_14085_, _14084_, _14083_);
  nor (_14086_, _10305_, _08430_);
  or (_14087_, _14086_, _10368_);
  or (_14088_, _10380_, _13990_);
  or (_14089_, _14088_, _14087_);
  and (_14090_, _14089_, _06407_);
  and (_14091_, _14090_, _14085_);
  and (_14092_, _14091_, _14081_);
  nor (_14093_, _10398_, _08430_);
  or (_14094_, _14093_, _10919_);
  or (_14095_, _10895_, _14018_);
  or (_14096_, _14095_, _14094_);
  and (_14097_, _14096_, _10897_);
  or (_14098_, _14097_, _14092_);
  and (_14099_, _10659_, \oc8051_golden_model_1.ACC [7]);
  or (_14100_, _14099_, _10949_);
  or (_14101_, _10927_, _10655_);
  or (_14102_, _14101_, _14100_);
  and (_14103_, _14102_, _10926_);
  and (_14104_, _14103_, _14098_);
  nand (_14105_, _10925_, \oc8051_golden_model_1.ACC [7]);
  nand (_14106_, _14105_, _10962_);
  or (_14107_, _14106_, _14104_);
  nor (_14108_, _10997_, _10763_);
  or (_14109_, _14108_, _10765_);
  and (_14110_, _14109_, _10957_);
  or (_14111_, _14110_, _10963_);
  and (_14112_, _14111_, _14107_);
  and (_14113_, _14109_, _10956_);
  or (_14114_, _14113_, _11003_);
  or (_14115_, _14114_, _14112_);
  and (_14116_, _11038_, _10783_);
  not (_14117_, _10781_);
  or (_14118_, _11005_, _10782_);
  and (_14119_, _14118_, _14117_);
  or (_14120_, _14119_, _11041_);
  or (_14121_, _14120_, _14116_);
  and (_14122_, _14121_, _06171_);
  and (_14123_, _14122_, _14115_);
  not (_14124_, _08809_);
  not (_14125_, _08808_);
  nand (_14126_, _10297_, _14125_);
  and (_14127_, _14126_, _06169_);
  and (_14128_, _14127_, _14124_);
  or (_14129_, _14128_, _10264_);
  or (_14130_, _14129_, _14123_);
  not (_14131_, _10793_);
  or (_14132_, _11080_, _10792_);
  and (_14133_, _14132_, _10264_);
  nand (_14134_, _14133_, _14131_);
  and (_14135_, _14134_, _06829_);
  and (_14136_, _14135_, _14130_);
  and (_14137_, _13848_, _06433_);
  nor (_14138_, _14137_, _14136_);
  nor (_14139_, _14138_, _11094_);
  or (_14140_, _14139_, _13832_);
  and (_14141_, _14140_, _05749_);
  and (_14142_, _13877_, _05748_);
  or (_14143_, _14142_, _06440_);
  or (_14144_, _14143_, _14141_);
  and (_14145_, _08345_, _07794_);
  or (_14146_, _13833_, _06444_);
  or (_14147_, _14146_, _14145_);
  and (_14148_, _14147_, _01317_);
  and (_14149_, _14148_, _14144_);
  or (_14150_, _14149_, _13831_);
  and (_41005_, _14150_, _43100_);
  nor (_14151_, _07593_, _07418_);
  nor (_14152_, _14151_, _07747_);
  nor (_14153_, _07418_, _07174_);
  nor (_14154_, _14153_, _07419_);
  and (_14155_, _14154_, _07417_);
  and (_14156_, _14155_, _14152_);
  or (_14157_, _14156_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_14158_, _07764_, _07755_);
  nor (_14159_, _07765_, _14158_);
  and (_14160_, _14159_, _07178_);
  and (_14161_, _14160_, _07764_);
  not (_14162_, _14161_);
  and (_14163_, _14162_, _14157_);
  not (_14164_, _14156_);
  nand (_14165_, _05823_, _05444_);
  not (_14166_, _08825_);
  or (_14167_, _08211_, _08708_);
  and (_14168_, _14167_, _08820_);
  or (_14169_, _12660_, _07772_);
  nand (_14170_, _07772_, _10693_);
  and (_14171_, _14170_, _14169_);
  and (_14172_, _14171_, _07103_);
  or (_14173_, _08211_, _06251_);
  not (_14174_, _07772_);
  and (_14175_, _12660_, _14174_);
  or (_14176_, _14175_, _08398_);
  nor (_14177_, _08443_, _07049_);
  and (_14178_, _06581_, \oc8051_golden_model_1.PC [0]);
  nor (_14179_, _06581_, _05855_);
  or (_14180_, _14179_, _14178_);
  and (_14181_, _14180_, _08443_);
  or (_14182_, _14181_, _14177_);
  and (_14183_, _14182_, _08429_);
  nor (_14184_, _08211_, _08429_);
  or (_14185_, _14184_, _14183_);
  and (_14186_, _14185_, _08428_);
  and (_14187_, _14169_, _06159_);
  or (_14188_, _14187_, _07485_);
  or (_14189_, _14188_, _14186_);
  nor (_14190_, _05764_, \oc8051_golden_model_1.PC [0]);
  nor (_14191_, _14190_, _07076_);
  and (_14192_, _14191_, _14189_);
  and (_14193_, _07076_, _07049_);
  or (_14194_, _14193_, _07086_);
  or (_14195_, _14194_, _14192_);
  and (_14196_, _14195_, _14176_);
  or (_14197_, _14196_, _06151_);
  or (_14198_, _08211_, _07191_);
  and (_14199_, _14198_, _06149_);
  and (_14200_, _14199_, _14197_);
  nor (_14201_, _12661_, _06149_);
  and (_14202_, _14201_, _14169_);
  or (_14203_, _14202_, _14200_);
  and (_14204_, _14203_, _05760_);
  or (_14205_, _05760_, _05444_);
  nand (_14206_, _06251_, _14205_);
  or (_14207_, _14206_, _14204_);
  and (_14208_, _14207_, _14173_);
  or (_14209_, _14208_, _06701_);
  and (_14210_, _09160_, _06172_);
  or (_14211_, _08209_, _07104_);
  or (_14212_, _14211_, _14210_);
  and (_14213_, _14212_, _08580_);
  and (_14214_, _14213_, _14209_);
  or (_14215_, _14214_, _14172_);
  or (_14216_, _14215_, _05791_);
  and (_14217_, _05791_, _05444_);
  nor (_14218_, _14217_, _08591_);
  and (_14219_, _14218_, _14216_);
  and (_14220_, _08591_, _07049_);
  or (_14221_, _14220_, _08595_);
  or (_14222_, _14221_, _14219_);
  or (_14223_, _09160_, _08601_);
  and (_14224_, _14223_, _08600_);
  and (_14225_, _14224_, _14222_);
  and (_14226_, _08395_, _07049_);
  and (_14227_, _08765_, \oc8051_golden_model_1.DPL [0]);
  and (_14228_, _08760_, \oc8051_golden_model_1.DPH [0]);
  and (_14229_, _08758_, \oc8051_golden_model_1.SP [0]);
  or (_14230_, _14229_, _14228_);
  or (_14231_, _14230_, _14227_);
  and (_14232_, _08726_, \oc8051_golden_model_1.TCON [0]);
  and (_14233_, _08775_, \oc8051_golden_model_1.TMOD [0]);
  and (_14234_, _08773_, \oc8051_golden_model_1.TL0 [0]);
  or (_14235_, _14234_, _14233_);
  or (_14236_, _14235_, _14232_);
  or (_14237_, _14236_, _14231_);
  and (_14238_, _08734_, \oc8051_golden_model_1.PSW [0]);
  and (_14239_, _08738_, \oc8051_golden_model_1.ACC [0]);
  and (_14240_, _08741_, \oc8051_golden_model_1.B [0]);
  or (_14241_, _14240_, _14239_);
  or (_14242_, _14241_, _14238_);
  and (_14243_, _08746_, \oc8051_golden_model_1.IP [0]);
  and (_14244_, _08749_, \oc8051_golden_model_1.IE [0]);
  and (_14245_, _08752_, \oc8051_golden_model_1.SBUF [0]);
  or (_14246_, _14245_, _14244_);
  or (_14247_, _14246_, _14243_);
  or (_14248_, _14247_, _14242_);
  and (_14249_, _08724_, \oc8051_golden_model_1.TL1 [0]);
  and (_14250_, _08710_, \oc8051_golden_model_1.TH1 [0]);
  and (_14251_, _08718_, \oc8051_golden_model_1.SCON [0]);
  or (_14252_, _14251_, _14250_);
  or (_14253_, _14252_, _14249_);
  and (_14254_, _08706_, \oc8051_golden_model_1.TH0 [0]);
  and (_14255_, _08770_, \oc8051_golden_model_1.PCON [0]);
  or (_14256_, _14255_, _14254_);
  or (_14257_, _14256_, _14253_);
  or (_14258_, _14257_, _14248_);
  or (_14259_, _14258_, _14237_);
  or (_14260_, _14259_, _14226_);
  and (_14261_, _14260_, _08599_);
  or (_14262_, _14261_, _08788_);
  or (_14263_, _14262_, _14225_);
  and (_14264_, _08788_, _06107_);
  nor (_14265_, _14264_, _06112_);
  and (_14266_, _14265_, _14263_);
  and (_14267_, _08708_, _06112_);
  or (_14268_, _14267_, _06076_);
  or (_14269_, _14268_, _14266_);
  nor (_14270_, _05836_, \oc8051_golden_model_1.PC [0]);
  nor (_14271_, _14270_, _07128_);
  and (_14272_, _14271_, _14269_);
  and (_14273_, _08211_, _08708_);
  not (_14274_, _14273_);
  and (_14275_, _14274_, _14167_);
  and (_14276_, _14275_, _07128_);
  or (_14277_, _14276_, _14272_);
  and (_14278_, _14277_, _08807_);
  nor (_14279_, _12322_, _08807_);
  or (_14280_, _14279_, _07133_);
  or (_14281_, _14280_, _14278_);
  or (_14282_, _14273_, _08806_);
  and (_14283_, _14282_, _08364_);
  and (_14284_, _14283_, _14281_);
  and (_14285_, _10276_, _07131_);
  or (_14286_, _14285_, _07124_);
  or (_14287_, _14286_, _14284_);
  nor (_14288_, _05848_, \oc8051_golden_model_1.PC [0]);
  nor (_14289_, _14288_, _08820_);
  and (_14290_, _14289_, _14287_);
  or (_14291_, _14290_, _14168_);
  and (_14292_, _14291_, _14166_);
  nor (_14293_, _12321_, _14166_);
  or (_14294_, _14293_, _07142_);
  or (_14295_, _14294_, _14292_);
  or (_14296_, _05846_, \oc8051_golden_model_1.PC [0]);
  and (_14297_, _14296_, _08362_);
  and (_14298_, _14297_, _14295_);
  nor (_14299_, _08362_, _07049_);
  or (_14300_, _14299_, _14298_);
  and (_14301_, _14300_, _07154_);
  nor (_14302_, _09160_, _07154_);
  or (_14303_, _14302_, _07152_);
  or (_14304_, _14303_, _14301_);
  nand (_14305_, _08211_, _07152_);
  and (_14306_, _14305_, _12723_);
  and (_14307_, _14306_, _14304_);
  and (_14308_, _06310_, _05444_);
  or (_14309_, _14308_, _05823_);
  or (_14310_, _14309_, _14307_);
  and (_14311_, _14310_, _14165_);
  or (_14312_, _14311_, _06073_);
  or (_14313_, _14175_, _06074_);
  and (_14314_, _14313_, _09193_);
  and (_14315_, _14314_, _14312_);
  nor (_14316_, _09193_, _07049_);
  or (_14317_, _14316_, _14315_);
  and (_14318_, _14317_, _07169_);
  nor (_14319_, _09160_, _07169_);
  or (_14320_, _14319_, _07167_);
  or (_14321_, _14320_, _14318_);
  nand (_14322_, _08211_, _07167_);
  and (_14323_, _14322_, _07417_);
  and (_14324_, _14323_, _14321_);
  or (_14325_, _14324_, _14164_);
  and (_14326_, _14325_, _14163_);
  and (_14327_, _07764_, _07178_);
  and (_14328_, _14327_, _14159_);
  nand (_14329_, _12057_, _06310_);
  or (_14330_, _12224_, _06310_);
  and (_14331_, _14330_, _14329_);
  and (_14332_, _14331_, _07764_);
  and (_14333_, _14332_, _14328_);
  or (_41013_, _14333_, _14326_);
  or (_14334_, _14156_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_14335_, _14334_, _14162_);
  and (_14336_, _06284_, _05820_);
  nor (_14337_, _09212_, _09161_);
  and (_14338_, _14337_, _14336_);
  not (_14339_, _14336_);
  or (_14340_, _09195_, _08352_);
  nor (_14341_, _14340_, _09193_);
  nor (_14342_, _05846_, \oc8051_golden_model_1.PC [1]);
  nand (_14343_, _08175_, _06945_);
  nor (_14344_, _08175_, _06945_);
  not (_14345_, _14344_);
  and (_14346_, _14345_, _14343_);
  and (_14347_, _14346_, _07128_);
  not (_14348_, _07781_);
  and (_14349_, _12627_, _14348_);
  and (_14350_, _07781_, \oc8051_golden_model_1.PSW [7]);
  or (_14351_, _14350_, _14349_);
  and (_14352_, _14351_, _07103_);
  nand (_14353_, _08175_, _06252_);
  or (_14354_, _14349_, _08398_);
  or (_14355_, _14340_, _08443_);
  nor (_14356_, _06581_, _05887_);
  and (_14357_, _06581_, _05407_);
  or (_14358_, _14357_, _14356_);
  nor (_14359_, _14358_, _07377_);
  nand (_14360_, _14359_, _07667_);
  and (_14361_, _14360_, _14355_);
  and (_14362_, _14361_, _08429_);
  nor (_14363_, _08541_, _08212_);
  nor (_14364_, _14363_, _08429_);
  or (_14365_, _14364_, _14362_);
  or (_14366_, _14365_, _06159_);
  or (_14367_, _12627_, _07781_);
  or (_14368_, _14367_, _08428_);
  and (_14369_, _14368_, _14366_);
  or (_14370_, _14369_, _07485_);
  nor (_14371_, _05764_, _05407_);
  nor (_14372_, _14371_, _07076_);
  and (_14373_, _14372_, _14370_);
  and (_14374_, _07306_, _07076_);
  or (_14375_, _14374_, _07086_);
  or (_14376_, _14375_, _14373_);
  and (_14377_, _14376_, _14354_);
  or (_14378_, _14377_, _06151_);
  nand (_14379_, _08175_, _06151_);
  and (_14380_, _14379_, _06149_);
  and (_14381_, _14380_, _14378_);
  not (_14382_, _12628_);
  and (_14383_, _14367_, _14382_);
  and (_14384_, _14383_, _06148_);
  or (_14385_, _14384_, _14381_);
  and (_14386_, _14385_, _05760_);
  or (_14387_, _05760_, \oc8051_golden_model_1.PC [1]);
  nand (_14388_, _06251_, _14387_);
  or (_14389_, _14388_, _14386_);
  and (_14390_, _14389_, _14353_);
  or (_14391_, _14390_, _06701_);
  and (_14392_, _09115_, _06172_);
  or (_14393_, _08173_, _07104_);
  or (_14394_, _14393_, _14392_);
  and (_14395_, _14394_, _08580_);
  and (_14396_, _14395_, _14391_);
  or (_14397_, _14396_, _14352_);
  or (_14398_, _14397_, _05791_);
  and (_14399_, _05791_, \oc8051_golden_model_1.PC [1]);
  nor (_14400_, _14399_, _08591_);
  and (_14401_, _14400_, _14398_);
  and (_14402_, _07306_, _08591_);
  or (_14403_, _14402_, _08595_);
  or (_14404_, _14403_, _14401_);
  or (_14405_, _09115_, _08601_);
  and (_14406_, _14405_, _08600_);
  and (_14407_, _14406_, _14404_);
  and (_14408_, _08395_, _07306_);
  and (_14409_, _08773_, \oc8051_golden_model_1.TL0 [1]);
  and (_14410_, _08775_, \oc8051_golden_model_1.TMOD [1]);
  and (_14411_, _08710_, \oc8051_golden_model_1.TH1 [1]);
  or (_14412_, _14411_, _14410_);
  or (_14413_, _14412_, _14409_);
  and (_14414_, _08724_, \oc8051_golden_model_1.TL1 [1]);
  and (_14415_, _08770_, \oc8051_golden_model_1.PCON [1]);
  and (_14416_, _08760_, \oc8051_golden_model_1.DPH [1]);
  or (_14417_, _14416_, _14415_);
  or (_14418_, _14417_, _14414_);
  and (_14419_, _08738_, \oc8051_golden_model_1.ACC [1]);
  and (_14420_, _08741_, \oc8051_golden_model_1.B [1]);
  or (_14421_, _14420_, _14419_);
  and (_14422_, _08749_, \oc8051_golden_model_1.IE [1]);
  and (_14423_, _08746_, \oc8051_golden_model_1.IP [1]);
  or (_14424_, _14423_, _14422_);
  or (_14425_, _14424_, _14421_);
  and (_14426_, _08765_, \oc8051_golden_model_1.DPL [1]);
  and (_14427_, _08758_, \oc8051_golden_model_1.SP [1]);
  or (_14428_, _14427_, _14426_);
  or (_14429_, _14428_, _14425_);
  and (_14430_, _08706_, \oc8051_golden_model_1.TH0 [1]);
  and (_14431_, _08726_, \oc8051_golden_model_1.TCON [1]);
  and (_14432_, _08734_, \oc8051_golden_model_1.PSW [1]);
  or (_14433_, _14432_, _14431_);
  and (_14434_, _08718_, \oc8051_golden_model_1.SCON [1]);
  and (_14435_, _08752_, \oc8051_golden_model_1.SBUF [1]);
  or (_14436_, _14435_, _14434_);
  or (_14437_, _14436_, _14433_);
  or (_14438_, _14437_, _14430_);
  or (_14439_, _14438_, _14429_);
  or (_14440_, _14439_, _14418_);
  or (_14441_, _14440_, _14413_);
  or (_14442_, _14441_, _14408_);
  and (_14443_, _14442_, _08599_);
  or (_14444_, _14443_, _08788_);
  or (_14445_, _14444_, _14407_);
  and (_14446_, _08788_, _06912_);
  nor (_14447_, _14446_, _06112_);
  and (_14448_, _14447_, _14445_);
  and (_14449_, _08763_, _06112_);
  or (_14450_, _14449_, _06076_);
  or (_14451_, _14450_, _14448_);
  nor (_14452_, _05836_, _05407_);
  nor (_14453_, _14452_, _07128_);
  and (_14454_, _14453_, _14451_);
  or (_14455_, _14454_, _14347_);
  and (_14456_, _14455_, _08807_);
  and (_14457_, _10278_, _07126_);
  or (_14458_, _14457_, _07133_);
  or (_14459_, _14458_, _14456_);
  or (_14460_, _14344_, _08806_);
  and (_14461_, _14460_, _08364_);
  and (_14462_, _14461_, _14459_);
  and (_14463_, _10275_, _07131_);
  or (_14464_, _14463_, _07124_);
  or (_14465_, _14464_, _14462_);
  nor (_14466_, _05848_, _05407_);
  nor (_14467_, _14466_, _08820_);
  and (_14468_, _14467_, _14465_);
  and (_14469_, _14343_, _08820_);
  or (_14470_, _14469_, _08825_);
  or (_14471_, _14470_, _14468_);
  nand (_14472_, _10277_, _08825_);
  and (_14473_, _14472_, _05846_);
  and (_14474_, _14473_, _14471_);
  nor (_14475_, _14474_, _14342_);
  nor (_14476_, _14475_, _06530_);
  and (_14477_, _14340_, _06530_);
  or (_14478_, _14477_, _06565_);
  or (_14479_, _14478_, _14476_);
  not (_14480_, _06972_);
  or (_14481_, _14340_, _06564_);
  and (_14482_, _14481_, _14480_);
  and (_14483_, _14482_, _14479_);
  and (_14484_, _14340_, _06972_);
  or (_14485_, _14484_, _07325_);
  or (_14486_, _14485_, _14483_);
  and (_14487_, _06284_, _05591_);
  not (_14488_, _14487_);
  or (_14489_, _14340_, _07326_);
  and (_14490_, _14489_, _14488_);
  and (_14491_, _14490_, _14486_);
  nand (_14492_, _14337_, _06276_);
  and (_14493_, _14492_, _07153_);
  or (_14494_, _14493_, _14491_);
  and (_14495_, _06281_, _05591_);
  nand (_14496_, _14337_, _14495_);
  and (_14497_, _14496_, _08837_);
  and (_14498_, _14497_, _14494_);
  nor (_14499_, _14363_, _08837_);
  or (_14500_, _14499_, _06310_);
  or (_14501_, _14500_, _14498_);
  nand (_14502_, _06310_, _05879_);
  and (_14503_, _14502_, _12730_);
  and (_14504_, _14503_, _14501_);
  and (_14505_, _05823_, _05407_);
  or (_14506_, _06073_, _14505_);
  or (_14507_, _14506_, _14504_);
  or (_14508_, _14349_, _06074_);
  and (_14509_, _14508_, _09193_);
  and (_14510_, _14509_, _14507_);
  or (_14511_, _14510_, _14341_);
  and (_14512_, _14511_, _14339_);
  or (_14513_, _14512_, _14338_);
  and (_14514_, _14513_, _06835_);
  and (_14515_, _14337_, _06834_);
  or (_14516_, _14515_, _07167_);
  or (_14517_, _14516_, _14514_);
  not (_14518_, _07167_);
  or (_14519_, _14363_, _14518_);
  and (_14520_, _14519_, _07417_);
  and (_14521_, _14520_, _14517_);
  or (_14522_, _14521_, _14164_);
  and (_14523_, _14522_, _14335_);
  nand (_14524_, _11997_, _06310_);
  or (_14525_, _12172_, _06310_);
  and (_14526_, _14525_, _14524_);
  and (_14527_, _14526_, _07764_);
  and (_14528_, _14527_, _14328_);
  or (_41014_, _14528_, _14523_);
  or (_14529_, _14156_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_14530_, _14529_, _14162_);
  nor (_14531_, _05923_, _05846_);
  and (_14532_, _09211_, _06172_);
  or (_14533_, _14532_, _08245_);
  and (_14534_, _14533_, _06701_);
  not (_14535_, _07848_);
  and (_14536_, _12644_, _14535_);
  or (_14537_, _14536_, _08398_);
  or (_14538_, _12644_, _07848_);
  or (_14539_, _14538_, _08428_);
  nand (_14540_, _08541_, _08247_);
  or (_14541_, _08541_, _08247_);
  nand (_14542_, _14541_, _14540_);
  and (_14543_, _14542_, _06162_);
  and (_14544_, _08352_, _07657_);
  nor (_14545_, _08352_, _07657_);
  nor (_14546_, _14545_, _14544_);
  nand (_14547_, _14546_, _08445_);
  and (_14548_, _06581_, _05921_);
  nor (_14549_, _06581_, _09981_);
  nor (_14550_, _14549_, _14548_);
  and (_14551_, _14550_, _08443_);
  nor (_14552_, _14551_, _06162_);
  and (_14553_, _14552_, _14547_);
  or (_14554_, _14553_, _06159_);
  or (_14555_, _14554_, _14543_);
  and (_14556_, _14555_, _14539_);
  or (_14557_, _14556_, _07485_);
  nor (_14558_, _05921_, _05764_);
  nor (_14559_, _14558_, _07076_);
  and (_14560_, _14559_, _14557_);
  and (_14561_, _07708_, _07076_);
  or (_14562_, _14561_, _07086_);
  or (_14563_, _14562_, _14560_);
  and (_14564_, _14563_, _14537_);
  or (_14565_, _14564_, _06151_);
  nand (_14566_, _08247_, _06151_);
  and (_14567_, _14566_, _06149_);
  and (_14568_, _14567_, _14565_);
  not (_14569_, _12645_);
  and (_14570_, _14538_, _14569_);
  and (_14571_, _14570_, _06148_);
  or (_14572_, _14571_, _14568_);
  and (_14573_, _14572_, _05760_);
  or (_14574_, _05923_, _05760_);
  nand (_14575_, _06251_, _14574_);
  or (_14576_, _14575_, _14573_);
  nand (_14577_, _08247_, _06252_);
  and (_14578_, _14577_, _07104_);
  and (_14579_, _14578_, _14576_);
  or (_14580_, _14579_, _14534_);
  and (_14581_, _14580_, _08580_);
  and (_14582_, _07848_, \oc8051_golden_model_1.PSW [7]);
  or (_14583_, _14582_, _14536_);
  and (_14584_, _14583_, _07103_);
  or (_14585_, _14584_, _05791_);
  or (_14586_, _14585_, _14581_);
  and (_14587_, _05923_, _05791_);
  nor (_14588_, _14587_, _08591_);
  and (_14589_, _14588_, _14586_);
  and (_14590_, _07708_, _08591_);
  or (_14591_, _14590_, _08595_);
  or (_14592_, _14591_, _14589_);
  or (_14593_, _09211_, _08601_);
  and (_14594_, _14593_, _08600_);
  and (_14595_, _14594_, _14592_);
  and (_14596_, _08395_, _07708_);
  and (_14597_, _08724_, \oc8051_golden_model_1.TL1 [2]);
  and (_14598_, _08710_, \oc8051_golden_model_1.TH1 [2]);
  and (_14599_, _08718_, \oc8051_golden_model_1.SCON [2]);
  or (_14600_, _14599_, _14598_);
  or (_14601_, _14600_, _14597_);
  and (_14602_, _08706_, \oc8051_golden_model_1.TH0 [2]);
  and (_14603_, _08726_, \oc8051_golden_model_1.TCON [2]);
  or (_14604_, _14603_, _14602_);
  or (_14605_, _14604_, _14601_);
  and (_14606_, _08734_, \oc8051_golden_model_1.PSW [2]);
  and (_14607_, _08741_, \oc8051_golden_model_1.B [2]);
  and (_14608_, _08738_, \oc8051_golden_model_1.ACC [2]);
  or (_14609_, _14608_, _14607_);
  or (_14610_, _14609_, _14606_);
  and (_14611_, _08746_, \oc8051_golden_model_1.IP [2]);
  and (_14612_, _08749_, \oc8051_golden_model_1.IE [2]);
  and (_14613_, _08752_, \oc8051_golden_model_1.SBUF [2]);
  or (_14614_, _14613_, _14612_);
  or (_14615_, _14614_, _14611_);
  or (_14616_, _14615_, _14610_);
  and (_14617_, _08760_, \oc8051_golden_model_1.DPH [2]);
  and (_14618_, _08758_, \oc8051_golden_model_1.SP [2]);
  or (_14619_, _14618_, _14617_);
  and (_14620_, _08765_, \oc8051_golden_model_1.DPL [2]);
  or (_14621_, _14620_, _14619_);
  and (_14622_, _08770_, \oc8051_golden_model_1.PCON [2]);
  and (_14623_, _08775_, \oc8051_golden_model_1.TMOD [2]);
  and (_14624_, _08773_, \oc8051_golden_model_1.TL0 [2]);
  or (_14625_, _14624_, _14623_);
  or (_14626_, _14625_, _14622_);
  or (_14627_, _14626_, _14621_);
  or (_14628_, _14627_, _14616_);
  or (_14629_, _14628_, _14605_);
  or (_14630_, _14629_, _14596_);
  and (_14631_, _14630_, _08599_);
  or (_14632_, _14631_, _08788_);
  or (_14633_, _14632_, _14595_);
  and (_14634_, _08788_, _06625_);
  nor (_14635_, _14634_, _06112_);
  and (_14636_, _14635_, _14633_);
  and (_14637_, _08768_, _06112_);
  or (_14638_, _14637_, _06076_);
  or (_14639_, _14638_, _14636_);
  nor (_14640_, _05921_, _05836_);
  nor (_14641_, _14640_, _07128_);
  and (_14642_, _14641_, _14639_);
  nand (_14643_, _08247_, _06521_);
  nor (_14644_, _08247_, _06521_);
  not (_14645_, _14644_);
  and (_14646_, _14645_, _14643_);
  and (_14647_, _14646_, _07128_);
  or (_14648_, _14647_, _14642_);
  and (_14649_, _14648_, _08807_);
  and (_14650_, _10282_, _07126_);
  or (_14651_, _14650_, _14649_);
  and (_14652_, _14651_, _08806_);
  and (_14653_, _14644_, _07133_);
  or (_14654_, _14653_, _14652_);
  and (_14655_, _14654_, _08364_);
  and (_14656_, _10274_, _07131_);
  or (_14657_, _14656_, _07124_);
  or (_14658_, _14657_, _14655_);
  nor (_14659_, _05921_, _05848_);
  nor (_14660_, _14659_, _08820_);
  and (_14661_, _14660_, _14658_);
  and (_14662_, _14643_, _08820_);
  or (_14663_, _14662_, _08825_);
  or (_14664_, _14663_, _14661_);
  nand (_14665_, _10281_, _08825_);
  and (_14666_, _14665_, _05846_);
  and (_14667_, _14666_, _14664_);
  or (_14668_, _14667_, _14531_);
  and (_14669_, _14668_, _08361_);
  nor (_14670_, _14546_, _08361_);
  or (_14671_, _14670_, _07325_);
  nor (_14672_, _14671_, _14669_);
  and (_14673_, _14546_, _07325_);
  or (_14674_, _14673_, _14487_);
  nor (_14675_, _14674_, _14672_);
  nor (_14676_, _09161_, _09070_);
  nor (_14677_, _14676_, _09162_);
  nand (_14678_, _14677_, _06276_);
  and (_14679_, _14678_, _07153_);
  or (_14680_, _14679_, _14675_);
  nand (_14681_, _14677_, _14495_);
  and (_14682_, _14681_, _08837_);
  and (_14683_, _14682_, _14680_);
  and (_14684_, _14542_, _07152_);
  or (_14685_, _14684_, _06310_);
  or (_14686_, _14685_, _14683_);
  nand (_14687_, _12029_, _06310_);
  and (_14688_, _14687_, _12730_);
  and (_14689_, _14688_, _14686_);
  and (_14690_, _05921_, _05823_);
  or (_14691_, _06073_, _14690_);
  or (_14692_, _14691_, _14689_);
  or (_14693_, _14536_, _06074_);
  and (_14694_, _14693_, _09193_);
  and (_14695_, _14694_, _14692_);
  nor (_14696_, _09195_, _07708_);
  nor (_14697_, _14696_, _09196_);
  and (_14698_, _14697_, _09189_);
  or (_14699_, _14698_, _14336_);
  or (_14700_, _14699_, _14695_);
  nor (_14701_, _09212_, _09211_);
  nor (_14702_, _14701_, _09213_);
  or (_14703_, _14702_, _14339_);
  and (_14704_, _14703_, _14700_);
  and (_14705_, _14704_, _06835_);
  and (_14706_, _14702_, _06834_);
  or (_14707_, _14706_, _07167_);
  or (_14708_, _14707_, _14705_);
  nor (_14709_, _08248_, _08212_);
  nor (_14710_, _14709_, _08249_);
  or (_14711_, _14710_, _14518_);
  and (_14712_, _14711_, _07417_);
  and (_14713_, _14712_, _14708_);
  or (_14714_, _14713_, _14164_);
  and (_14715_, _14714_, _14530_);
  nand (_14716_, _11989_, _06310_);
  or (_14717_, _12159_, _06310_);
  and (_14718_, _14717_, _14716_);
  and (_14719_, _14718_, _07764_);
  and (_14720_, _14719_, _14328_);
  or (_41016_, _14720_, _14715_);
  or (_14721_, _14156_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_14722_, _14721_, _14162_);
  nor (_14723_, _06322_, _05846_);
  nand (_14724_, _08139_, _06389_);
  nor (_14725_, _08139_, _06389_);
  not (_14726_, _14725_);
  and (_14727_, _14726_, _14724_);
  and (_14728_, _14727_, _07128_);
  and (_14729_, _07851_, \oc8051_golden_model_1.PSW [7]);
  not (_14730_, _07851_);
  and (_14731_, _12595_, _14730_);
  or (_14732_, _14731_, _14729_);
  and (_14733_, _14732_, _07103_);
  or (_14734_, _14731_, _08398_);
  or (_14735_, _12595_, _07851_);
  or (_14736_, _14735_, _08428_);
  and (_14737_, _14540_, _08140_);
  or (_14738_, _14737_, _08543_);
  and (_14739_, _14738_, _06162_);
  nor (_14740_, _14544_, _07474_);
  nor (_14741_, _14740_, _08353_);
  nand (_14742_, _14741_, _08445_);
  and (_14743_, _06581_, _05974_);
  nor (_14744_, _06581_, _10028_);
  nor (_14745_, _14744_, _14743_);
  and (_14746_, _14745_, _08443_);
  nor (_14747_, _14746_, _06162_);
  and (_14748_, _14747_, _14742_);
  or (_14749_, _14748_, _06159_);
  or (_14750_, _14749_, _14739_);
  and (_14751_, _14750_, _14736_);
  or (_14752_, _14751_, _07485_);
  nor (_14753_, _05974_, _05764_);
  nor (_14754_, _14753_, _07076_);
  and (_14755_, _14754_, _14752_);
  and (_14756_, _07544_, _07076_);
  or (_14757_, _14756_, _07086_);
  or (_14758_, _14757_, _14755_);
  and (_14759_, _14758_, _14734_);
  or (_14760_, _14759_, _06151_);
  nand (_14761_, _08139_, _06151_);
  and (_14762_, _14761_, _06149_);
  and (_14763_, _14762_, _14760_);
  not (_14764_, _12596_);
  and (_14765_, _14735_, _14764_);
  and (_14766_, _14765_, _06148_);
  or (_14767_, _14766_, _14763_);
  and (_14768_, _14767_, _05760_);
  or (_14769_, _06322_, _05760_);
  nand (_14770_, _06251_, _14769_);
  or (_14771_, _14770_, _14768_);
  nand (_14772_, _08139_, _06252_);
  and (_14773_, _14772_, _14771_);
  or (_14774_, _14773_, _06701_);
  and (_14775_, _09210_, _06172_);
  or (_14776_, _08137_, _07104_);
  or (_14777_, _14776_, _14775_);
  and (_14778_, _14777_, _08580_);
  and (_14779_, _14778_, _14774_);
  or (_14780_, _14779_, _14733_);
  or (_14781_, _14780_, _05791_);
  and (_14782_, _06322_, _05791_);
  nor (_14783_, _14782_, _08591_);
  and (_14784_, _14783_, _14781_);
  and (_14785_, _07544_, _08591_);
  or (_14786_, _14785_, _08595_);
  or (_14787_, _14786_, _14784_);
  or (_14788_, _09210_, _08601_);
  and (_14789_, _14788_, _08600_);
  and (_14790_, _14789_, _14787_);
  and (_14791_, _08395_, _07544_);
  and (_14792_, _08724_, \oc8051_golden_model_1.TL1 [3]);
  and (_14793_, _08710_, \oc8051_golden_model_1.TH1 [3]);
  and (_14794_, _08718_, \oc8051_golden_model_1.SCON [3]);
  or (_14795_, _14794_, _14793_);
  or (_14796_, _14795_, _14792_);
  and (_14797_, _08770_, \oc8051_golden_model_1.PCON [3]);
  and (_14798_, _08706_, \oc8051_golden_model_1.TH0 [3]);
  or (_14799_, _14798_, _14797_);
  or (_14800_, _14799_, _14796_);
  and (_14801_, _08734_, \oc8051_golden_model_1.PSW [3]);
  and (_14802_, _08741_, \oc8051_golden_model_1.B [3]);
  and (_14803_, _08738_, \oc8051_golden_model_1.ACC [3]);
  or (_14804_, _14803_, _14802_);
  or (_14805_, _14804_, _14801_);
  and (_14806_, _08746_, \oc8051_golden_model_1.IP [3]);
  and (_14807_, _08749_, \oc8051_golden_model_1.IE [3]);
  and (_14808_, _08752_, \oc8051_golden_model_1.SBUF [3]);
  or (_14809_, _14808_, _14807_);
  or (_14810_, _14809_, _14806_);
  or (_14811_, _14810_, _14805_);
  and (_14812_, _08765_, \oc8051_golden_model_1.DPL [3]);
  and (_14813_, _08758_, \oc8051_golden_model_1.SP [3]);
  and (_14814_, _08760_, \oc8051_golden_model_1.DPH [3]);
  or (_14815_, _14814_, _14813_);
  or (_14816_, _14815_, _14812_);
  and (_14817_, _08775_, \oc8051_golden_model_1.TMOD [3]);
  and (_14818_, _08773_, \oc8051_golden_model_1.TL0 [3]);
  or (_14819_, _14818_, _14817_);
  and (_14820_, _08726_, \oc8051_golden_model_1.TCON [3]);
  or (_14821_, _14820_, _14819_);
  or (_14822_, _14821_, _14816_);
  or (_14823_, _14822_, _14811_);
  or (_14824_, _14823_, _14800_);
  or (_14825_, _14824_, _14791_);
  and (_14826_, _14825_, _08599_);
  or (_14827_, _14826_, _08788_);
  or (_14828_, _14827_, _14790_);
  and (_14829_, _08788_, _06070_);
  nor (_14830_, _14829_, _06112_);
  and (_14831_, _14830_, _14828_);
  and (_14832_, _08712_, _06112_);
  or (_14833_, _14832_, _06076_);
  or (_14834_, _14833_, _14831_);
  nor (_14835_, _05974_, _05836_);
  nor (_14836_, _14835_, _07128_);
  and (_14837_, _14836_, _14834_);
  or (_14838_, _14837_, _14728_);
  and (_14839_, _14838_, _08807_);
  and (_14840_, _12318_, _07126_);
  or (_14841_, _14840_, _07133_);
  or (_14842_, _14841_, _14839_);
  or (_14843_, _14725_, _08806_);
  and (_14844_, _14843_, _08364_);
  and (_14845_, _14844_, _14842_);
  and (_14846_, _10272_, _07131_);
  or (_14847_, _14846_, _07124_);
  or (_14848_, _14847_, _14845_);
  nor (_14849_, _05974_, _05848_);
  nor (_14850_, _14849_, _08820_);
  and (_14851_, _14850_, _14848_);
  and (_14852_, _14724_, _08820_);
  or (_14853_, _14852_, _08825_);
  or (_14854_, _14853_, _14851_);
  nand (_14855_, _10273_, _08825_);
  and (_14856_, _14855_, _05846_);
  and (_14857_, _14856_, _14854_);
  or (_14858_, _14857_, _14723_);
  and (_14859_, _14858_, _08361_);
  nor (_14860_, _14741_, _08361_);
  or (_14861_, _14860_, _07325_);
  nor (_14862_, _14861_, _14859_);
  and (_14863_, _14741_, _07325_);
  or (_14864_, _14863_, _14487_);
  nor (_14865_, _14864_, _14862_);
  nor (_14866_, _09162_, _09025_);
  nor (_14867_, _14866_, _09163_);
  nand (_14868_, _14867_, _06276_);
  and (_14869_, _14868_, _07153_);
  or (_14870_, _14869_, _14865_);
  nand (_14871_, _14867_, _14495_);
  and (_14872_, _14871_, _08837_);
  and (_14873_, _14872_, _14870_);
  and (_14874_, _14738_, _07152_);
  or (_14875_, _14874_, _06310_);
  or (_14876_, _14875_, _14873_);
  nand (_14877_, _12024_, _06310_);
  and (_14878_, _14877_, _12730_);
  and (_14879_, _14878_, _14876_);
  and (_14880_, _05974_, _05823_);
  or (_14881_, _06073_, _14880_);
  or (_14882_, _14881_, _14879_);
  or (_14883_, _14731_, _06074_);
  and (_14884_, _14883_, _09193_);
  and (_14885_, _14884_, _14882_);
  nor (_14886_, _09196_, _07544_);
  nor (_14887_, _14886_, _09197_);
  or (_14888_, _14887_, _07168_);
  and (_14889_, _14888_, _12737_);
  or (_14890_, _14889_, _14885_);
  nor (_14891_, _09213_, _09210_);
  nor (_14892_, _14891_, _09214_);
  or (_14893_, _14892_, _07169_);
  and (_14894_, _14893_, _14890_);
  or (_14895_, _14894_, _07167_);
  nor (_14896_, _08249_, _08140_);
  nor (_14897_, _14896_, _08250_);
  or (_14898_, _14897_, _14518_);
  and (_14899_, _14898_, _07417_);
  and (_14900_, _14899_, _14895_);
  or (_14901_, _14900_, _14164_);
  and (_14902_, _14901_, _14722_);
  nand (_14903_, _11982_, _06310_);
  or (_14904_, _12163_, _06310_);
  and (_14905_, _14904_, _14903_);
  and (_14906_, _14905_, _07764_);
  and (_14907_, _14906_, _14328_);
  or (_41017_, _14907_, _14902_);
  nor (_14908_, _14156_, _08284_);
  nor (_14909_, _09214_, _09209_);
  nor (_14910_, _14909_, _09215_);
  or (_14911_, _14910_, _07169_);
  nor (_14912_, _12194_, _05846_);
  and (_14913_, _08353_, _08349_);
  nor (_14914_, _08353_, _08349_);
  nor (_14915_, _14914_, _14913_);
  nand (_14916_, _14915_, _08445_);
  nor (_14917_, _06581_, _09902_);
  and (_14918_, _12193_, _06581_);
  nor (_14919_, _14918_, _14917_);
  nand (_14920_, _14919_, _08443_);
  and (_14921_, _14920_, _14916_);
  or (_14922_, _14921_, _07064_);
  or (_14923_, _09209_, _07065_);
  and (_14924_, _14923_, _14922_);
  and (_14925_, _14924_, _08429_);
  nand (_14926_, _08543_, _08338_);
  or (_14927_, _08543_, _08338_);
  nand (_14928_, _14927_, _14926_);
  and (_14929_, _14928_, _06162_);
  or (_14930_, _14929_, _14925_);
  and (_14931_, _14930_, _08428_);
  nand (_14932_, _12678_, _12676_);
  and (_14933_, _14932_, _06159_);
  or (_14934_, _14933_, _07485_);
  or (_14935_, _14934_, _14931_);
  nor (_14936_, _12193_, _05764_);
  nor (_14937_, _14936_, _07076_);
  and (_14938_, _14937_, _14935_);
  and (_14939_, _08336_, _07076_);
  or (_14940_, _14939_, _07086_);
  or (_14941_, _14940_, _14938_);
  nor (_14942_, _12677_, _12676_);
  or (_14943_, _14942_, _08398_);
  and (_14944_, _14943_, _14941_);
  or (_14945_, _14944_, _06151_);
  nand (_14946_, _08338_, _06151_);
  and (_14947_, _14946_, _06149_);
  and (_14948_, _14947_, _14945_);
  not (_14949_, _12679_);
  and (_14950_, _14932_, _14949_);
  and (_14951_, _14950_, _06148_);
  or (_14952_, _14951_, _14948_);
  and (_14953_, _14952_, _05760_);
  or (_14954_, _12194_, _05760_);
  nand (_14955_, _14954_, _06251_);
  or (_14956_, _14955_, _14953_);
  nand (_14957_, _08338_, _06252_);
  and (_14958_, _14957_, _14956_);
  or (_14959_, _14958_, _06701_);
  and (_14960_, _09209_, _06172_);
  or (_14961_, _08283_, _07104_);
  or (_14962_, _14961_, _14960_);
  and (_14963_, _14962_, _08580_);
  and (_14964_, _14963_, _14959_);
  and (_14965_, _12677_, \oc8051_golden_model_1.PSW [7]);
  or (_14966_, _14965_, _14942_);
  and (_14967_, _14966_, _07103_);
  or (_14968_, _14967_, _05791_);
  or (_14969_, _14968_, _14964_);
  and (_14970_, _12194_, _05791_);
  nor (_14971_, _14970_, _08591_);
  and (_14972_, _14971_, _14969_);
  and (_14973_, _08336_, _08591_);
  or (_14974_, _14973_, _08595_);
  or (_14975_, _14974_, _14972_);
  or (_14976_, _09209_, _08601_);
  and (_14977_, _14976_, _08600_);
  and (_14978_, _14977_, _14975_);
  and (_14979_, _08395_, _08336_);
  and (_14980_, _08710_, \oc8051_golden_model_1.TH1 [4]);
  and (_14981_, _08775_, \oc8051_golden_model_1.TMOD [4]);
  and (_14982_, _08706_, \oc8051_golden_model_1.TH0 [4]);
  or (_14983_, _14982_, _14981_);
  or (_14984_, _14983_, _14980_);
  and (_14985_, _08760_, \oc8051_golden_model_1.DPH [4]);
  and (_14986_, _08724_, \oc8051_golden_model_1.TL1 [4]);
  and (_14987_, _08758_, \oc8051_golden_model_1.SP [4]);
  or (_14988_, _14987_, _14986_);
  or (_14989_, _14988_, _14985_);
  and (_14990_, _08752_, \oc8051_golden_model_1.SBUF [4]);
  and (_14991_, _08746_, \oc8051_golden_model_1.IP [4]);
  or (_14992_, _14991_, _14990_);
  and (_14993_, _08718_, \oc8051_golden_model_1.SCON [4]);
  and (_14994_, _08741_, \oc8051_golden_model_1.B [4]);
  or (_14995_, _14994_, _14993_);
  or (_14996_, _14995_, _14992_);
  and (_14997_, _08765_, \oc8051_golden_model_1.DPL [4]);
  and (_14998_, _08770_, \oc8051_golden_model_1.PCON [4]);
  or (_14999_, _14998_, _14997_);
  or (_15000_, _14999_, _14996_);
  and (_15001_, _08773_, \oc8051_golden_model_1.TL0 [4]);
  and (_15002_, _08726_, \oc8051_golden_model_1.TCON [4]);
  and (_15003_, _08749_, \oc8051_golden_model_1.IE [4]);
  or (_15004_, _15003_, _15002_);
  and (_15005_, _08738_, \oc8051_golden_model_1.ACC [4]);
  and (_15006_, _08734_, \oc8051_golden_model_1.PSW [4]);
  or (_15007_, _15006_, _15005_);
  or (_15008_, _15007_, _15004_);
  or (_15009_, _15008_, _15001_);
  or (_15010_, _15009_, _15000_);
  or (_15011_, _15010_, _14989_);
  or (_15012_, _15011_, _14984_);
  or (_15013_, _15012_, _14979_);
  and (_15014_, _15013_, _08599_);
  or (_15015_, _15014_, _08788_);
  or (_15016_, _15015_, _14978_);
  and (_15017_, _08788_, _06876_);
  nor (_15018_, _15017_, _06112_);
  and (_15019_, _15018_, _15016_);
  and (_15020_, _08715_, _06112_);
  or (_15021_, _15020_, _06076_);
  or (_15022_, _15021_, _15019_);
  nor (_15023_, _12193_, _05836_);
  nor (_15024_, _15023_, _07128_);
  and (_15025_, _15024_, _15022_);
  nand (_15026_, _08670_, _08338_);
  nor (_15027_, _08670_, _08338_);
  not (_15028_, _15027_);
  and (_15029_, _15028_, _15026_);
  and (_15030_, _15029_, _07128_);
  or (_15031_, _15030_, _15025_);
  and (_15032_, _15031_, _08807_);
  and (_15033_, _10289_, _07126_);
  or (_15034_, _15033_, _07133_);
  or (_15035_, _15034_, _15032_);
  or (_15036_, _15027_, _08806_);
  and (_15037_, _15036_, _08364_);
  and (_15038_, _15037_, _15035_);
  and (_15039_, _10270_, _07131_);
  or (_15040_, _15039_, _07124_);
  or (_15041_, _15040_, _15038_);
  nor (_15042_, _12193_, _05848_);
  nor (_15043_, _15042_, _08820_);
  and (_15044_, _15043_, _15041_);
  and (_15045_, _15026_, _08820_);
  or (_15046_, _15045_, _08825_);
  or (_15047_, _15046_, _15044_);
  nand (_15048_, _10288_, _08825_);
  and (_15049_, _15048_, _05846_);
  and (_15050_, _15049_, _15047_);
  or (_15051_, _15050_, _14912_);
  and (_15052_, _15051_, _08361_);
  nor (_15053_, _14915_, _08361_);
  or (_15054_, _15053_, _07325_);
  nor (_15055_, _15054_, _15052_);
  and (_15056_, _14915_, _07325_);
  or (_15057_, _15056_, _14487_);
  nor (_15058_, _15057_, _15055_);
  nor (_15059_, _09163_, _08980_);
  nor (_15060_, _15059_, _09164_);
  nand (_15061_, _15060_, _06276_);
  and (_15062_, _15061_, _07153_);
  or (_15063_, _15062_, _15058_);
  nand (_15064_, _15060_, _14495_);
  and (_15065_, _15064_, _08837_);
  and (_15066_, _15065_, _15063_);
  and (_15067_, _14928_, _07152_);
  or (_15068_, _15067_, _06310_);
  or (_15069_, _15068_, _15066_);
  nand (_15070_, _12019_, _06310_);
  and (_15071_, _15070_, _12730_);
  and (_15072_, _15071_, _15069_);
  and (_15073_, _12193_, _05823_);
  or (_15074_, _15073_, _06073_);
  or (_15075_, _15074_, _15072_);
  or (_15076_, _14942_, _06074_);
  and (_15077_, _15076_, _09193_);
  and (_15078_, _15077_, _15075_);
  nor (_15079_, _09197_, _08336_);
  nor (_15080_, _15079_, _09198_);
  and (_15081_, _15080_, _09189_);
  or (_15082_, _15081_, _07168_);
  or (_15083_, _15082_, _15078_);
  and (_15084_, _15083_, _14911_);
  or (_15085_, _15084_, _07167_);
  nor (_15086_, _08339_, _08250_);
  nor (_15087_, _15086_, _08340_);
  or (_15088_, _15087_, _14518_);
  and (_15089_, _15088_, _07417_);
  and (_15090_, _15089_, _15085_);
  and (_15091_, _15090_, _14156_);
  or (_15092_, _15091_, _14908_);
  and (_15093_, _15092_, _14162_);
  nand (_15094_, _11978_, _06310_);
  or (_15095_, _12156_, _06310_);
  and (_15096_, _15095_, _15094_);
  and (_15097_, _15096_, _07764_);
  and (_15098_, _15097_, _14328_);
  or (_41018_, _15098_, _15093_);
  nor (_15099_, _14156_, _08049_);
  nor (_15100_, _09164_, _08931_);
  or (_15101_, _15100_, _09165_);
  and (_15102_, _15101_, _14495_);
  not (_15103_, _12612_);
  and (_15104_, _15103_, _12611_);
  or (_15105_, _15104_, _08398_);
  nor (_15106_, _06581_, _09930_);
  and (_15107_, _12188_, _06581_);
  or (_15108_, _15107_, _15106_);
  and (_15109_, _15108_, _08443_);
  nor (_15110_, _14913_, _08348_);
  or (_15111_, _15110_, _08354_);
  and (_15112_, _15111_, _08445_);
  or (_15113_, _15112_, _15109_);
  and (_15114_, _15113_, _07065_);
  and (_15115_, _09208_, _07064_);
  or (_15116_, _15115_, _15114_);
  and (_15117_, _15116_, _08429_);
  and (_15118_, _14926_, _08104_);
  or (_15119_, _15118_, _08544_);
  and (_15120_, _15119_, _06162_);
  or (_15121_, _15120_, _15117_);
  and (_15122_, _15121_, _08428_);
  or (_15123_, _12612_, _12611_);
  and (_15124_, _15123_, _06159_);
  or (_15125_, _15124_, _07485_);
  or (_15126_, _15125_, _15122_);
  nor (_15127_, _12188_, _05764_);
  nor (_15128_, _15127_, _07076_);
  and (_15129_, _15128_, _15126_);
  and (_15130_, _08101_, _07076_);
  or (_15131_, _15130_, _07086_);
  or (_15132_, _15131_, _15129_);
  and (_15133_, _15132_, _15105_);
  or (_15134_, _15133_, _06151_);
  nand (_15135_, _08103_, _06151_);
  and (_15136_, _15135_, _06149_);
  and (_15137_, _15136_, _15134_);
  not (_15138_, _12613_);
  and (_15139_, _15123_, _15138_);
  and (_15140_, _15139_, _06148_);
  or (_15141_, _15140_, _15137_);
  and (_15142_, _15141_, _05760_);
  or (_15143_, _12189_, _05760_);
  nand (_15144_, _15143_, _06251_);
  or (_15145_, _15144_, _15142_);
  nand (_15146_, _08103_, _06252_);
  and (_15147_, _15146_, _15145_);
  or (_15148_, _15147_, _06701_);
  and (_15149_, _09208_, _06172_);
  or (_15150_, _08048_, _07104_);
  or (_15151_, _15150_, _15149_);
  and (_15152_, _15151_, _08580_);
  and (_15153_, _15152_, _15148_);
  and (_15154_, _12612_, \oc8051_golden_model_1.PSW [7]);
  or (_15155_, _15154_, _15104_);
  and (_15156_, _15155_, _07103_);
  or (_15157_, _15156_, _05791_);
  or (_15158_, _15157_, _15153_);
  and (_15159_, _12189_, _05791_);
  nor (_15160_, _15159_, _08591_);
  and (_15161_, _15160_, _15158_);
  and (_15162_, _08101_, _08591_);
  or (_15163_, _15162_, _08595_);
  or (_15164_, _15163_, _15161_);
  or (_15165_, _09208_, _08601_);
  and (_15166_, _15165_, _08600_);
  and (_15167_, _15166_, _15164_);
  and (_15168_, _08395_, _08101_);
  and (_15169_, _08775_, \oc8051_golden_model_1.TMOD [5]);
  and (_15170_, _08706_, \oc8051_golden_model_1.TH0 [5]);
  and (_15171_, _08710_, \oc8051_golden_model_1.TH1 [5]);
  or (_15172_, _15171_, _15170_);
  or (_15173_, _15172_, _15169_);
  and (_15174_, _08770_, \oc8051_golden_model_1.PCON [5]);
  and (_15175_, _08724_, \oc8051_golden_model_1.TL1 [5]);
  and (_15176_, _08758_, \oc8051_golden_model_1.SP [5]);
  or (_15177_, _15176_, _15175_);
  or (_15178_, _15177_, _15174_);
  and (_15179_, _08741_, \oc8051_golden_model_1.B [5]);
  and (_15180_, _08738_, \oc8051_golden_model_1.ACC [5]);
  or (_15181_, _15180_, _15179_);
  and (_15182_, _08718_, \oc8051_golden_model_1.SCON [5]);
  and (_15183_, _08734_, \oc8051_golden_model_1.PSW [5]);
  or (_15184_, _15183_, _15182_);
  or (_15185_, _15184_, _15181_);
  and (_15186_, _08765_, \oc8051_golden_model_1.DPL [5]);
  and (_15187_, _08760_, \oc8051_golden_model_1.DPH [5]);
  or (_15188_, _15187_, _15186_);
  or (_15189_, _15188_, _15185_);
  and (_15190_, _08773_, \oc8051_golden_model_1.TL0 [5]);
  and (_15191_, _08752_, \oc8051_golden_model_1.SBUF [5]);
  and (_15192_, _08749_, \oc8051_golden_model_1.IE [5]);
  or (_15193_, _15192_, _15191_);
  and (_15194_, _08726_, \oc8051_golden_model_1.TCON [5]);
  and (_15196_, _08746_, \oc8051_golden_model_1.IP [5]);
  or (_15197_, _15196_, _15194_);
  or (_15198_, _15197_, _15193_);
  or (_15199_, _15198_, _15190_);
  or (_15200_, _15199_, _15189_);
  or (_15201_, _15200_, _15178_);
  or (_15202_, _15201_, _15173_);
  or (_15203_, _15202_, _15168_);
  and (_15204_, _15203_, _08599_);
  or (_15205_, _15204_, _08788_);
  or (_15206_, _15205_, _15167_);
  and (_15207_, _08788_, _06477_);
  nor (_15208_, _15207_, _06112_);
  and (_15209_, _15208_, _15206_);
  and (_15210_, _08736_, _06112_);
  or (_15211_, _15210_, _06076_);
  or (_15212_, _15211_, _15209_);
  nor (_15213_, _12188_, _05836_);
  nor (_15214_, _15213_, _07128_);
  and (_15215_, _15214_, _15212_);
  nand (_15216_, _08701_, _08103_);
  nor (_15217_, _08701_, _08103_);
  not (_15218_, _15217_);
  and (_15219_, _15218_, _15216_);
  and (_15220_, _15219_, _07128_);
  or (_15221_, _15220_, _15215_);
  and (_15222_, _15221_, _08807_);
  and (_15223_, _12325_, _07126_);
  or (_15224_, _15223_, _07133_);
  or (_15225_, _15224_, _15222_);
  or (_15226_, _15217_, _08806_);
  and (_15227_, _15226_, _08364_);
  and (_15228_, _15227_, _15225_);
  and (_15229_, _10268_, _07131_);
  or (_15230_, _15229_, _07124_);
  or (_15231_, _15230_, _15228_);
  nor (_15232_, _12188_, _05848_);
  nor (_15233_, _15232_, _08820_);
  and (_15234_, _15233_, _15231_);
  and (_15235_, _15216_, _08820_);
  or (_15236_, _15235_, _08825_);
  or (_15237_, _15236_, _15234_);
  nand (_15238_, _10269_, _08825_);
  and (_15239_, _15238_, _05846_);
  and (_15240_, _15239_, _15237_);
  or (_15241_, _12189_, _05846_);
  nand (_15242_, _15241_, _08362_);
  or (_15243_, _15242_, _15240_);
  or (_15244_, _15111_, _08362_);
  and (_15245_, _15244_, _14488_);
  and (_15246_, _15245_, _15243_);
  and (_15247_, _15101_, _14487_);
  nor (_15248_, _15247_, _15246_);
  nor (_15249_, _15248_, _14495_);
  or (_15250_, _15249_, _15102_);
  and (_15251_, _15250_, _08837_);
  and (_15252_, _15119_, _07152_);
  or (_15253_, _15252_, _06310_);
  or (_15254_, _15253_, _15251_);
  nand (_15255_, _12014_, _06310_);
  and (_15256_, _15255_, _12730_);
  and (_15257_, _15256_, _15254_);
  and (_15258_, _12188_, _05823_);
  or (_15259_, _15258_, _06073_);
  or (_15260_, _15259_, _15257_);
  or (_15261_, _15104_, _06074_);
  and (_15262_, _15261_, _09193_);
  and (_15263_, _15262_, _15260_);
  nor (_15264_, _09198_, _08101_);
  nor (_15265_, _15264_, _09199_);
  or (_15266_, _15265_, _07168_);
  and (_15267_, _15266_, _12737_);
  or (_15268_, _15267_, _15263_);
  nor (_15269_, _09215_, _09208_);
  nor (_15270_, _15269_, _09216_);
  or (_15271_, _15270_, _07169_);
  and (_15272_, _15271_, _15268_);
  or (_15273_, _15272_, _07167_);
  nor (_15274_, _08340_, _08104_);
  nor (_15275_, _15274_, _08341_);
  or (_15276_, _15275_, _14518_);
  and (_15277_, _15276_, _07417_);
  and (_15278_, _15277_, _15273_);
  and (_15279_, _15278_, _14156_);
  or (_15280_, _15279_, _15099_);
  and (_15281_, _15280_, _14162_);
  nand (_15282_, _11973_, _06310_);
  or (_15283_, _12152_, _06310_);
  and (_15284_, _15283_, _15282_);
  and (_15285_, _15284_, _07764_);
  and (_15286_, _15285_, _14328_);
  or (_41020_, _15286_, _15281_);
  or (_15287_, _14156_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_15288_, _15287_, _14162_);
  nor (_15289_, _09216_, _09207_);
  nor (_15290_, _15289_, _09217_);
  or (_15291_, _15290_, _07169_);
  not (_15292_, _05820_);
  nor (_15293_, _06129_, _15292_);
  nor (_15294_, _12181_, _05846_);
  and (_15295_, _10295_, _07126_);
  not (_15296_, _12580_);
  and (_15297_, _15296_, _12579_);
  or (_15298_, _15297_, _08398_);
  nor (_15299_, _08544_, _08014_);
  or (_15300_, _15299_, _08545_);
  and (_15301_, _15300_, _06162_);
  or (_15302_, _09207_, _07065_);
  nor (_15303_, _08354_, _08347_);
  nor (_15304_, _15303_, _08355_);
  nor (_15305_, _15304_, _08443_);
  nand (_15306_, _12181_, _06581_);
  or (_15307_, _06581_, \oc8051_golden_model_1.ACC [6]);
  and (_15308_, _15307_, _15306_);
  and (_15309_, _15308_, _08443_);
  or (_15310_, _15309_, _07064_);
  or (_15311_, _15310_, _15305_);
  and (_15312_, _15311_, _08429_);
  and (_15313_, _15312_, _15302_);
  or (_15314_, _15313_, _15301_);
  and (_15315_, _15314_, _08428_);
  or (_15316_, _12580_, _12579_);
  and (_15317_, _15316_, _06159_);
  or (_15318_, _15317_, _07485_);
  or (_15319_, _15318_, _15315_);
  nor (_15320_, _12180_, _05764_);
  nor (_15321_, _15320_, _07076_);
  and (_15322_, _15321_, _15319_);
  and (_15323_, _08012_, _07076_);
  or (_15324_, _15323_, _07086_);
  or (_15325_, _15324_, _15322_);
  and (_15326_, _15325_, _15298_);
  or (_15327_, _15326_, _06151_);
  nand (_15328_, _08014_, _06151_);
  and (_15329_, _15328_, _06149_);
  and (_15330_, _15329_, _15327_);
  not (_15331_, _12581_);
  and (_15332_, _15316_, _15331_);
  and (_15333_, _15332_, _06148_);
  or (_15334_, _15333_, _15330_);
  and (_15335_, _15334_, _05760_);
  or (_15336_, _12181_, _05760_);
  nand (_15337_, _15336_, _06251_);
  or (_15338_, _15337_, _15335_);
  nand (_15339_, _08014_, _06252_);
  and (_15340_, _15339_, _15338_);
  or (_15341_, _15340_, _06701_);
  and (_15342_, _09207_, _06172_);
  or (_15343_, _07959_, _07104_);
  or (_15344_, _15343_, _15342_);
  and (_15345_, _15344_, _08580_);
  and (_15346_, _15345_, _15341_);
  and (_15347_, _12580_, \oc8051_golden_model_1.PSW [7]);
  or (_15348_, _15347_, _15297_);
  and (_15349_, _15348_, _07103_);
  or (_15350_, _15349_, _05791_);
  or (_15351_, _15350_, _15346_);
  and (_15352_, _12181_, _05791_);
  nor (_15353_, _15352_, _08591_);
  and (_15354_, _15353_, _15351_);
  and (_15355_, _08012_, _08591_);
  or (_15356_, _15355_, _08595_);
  or (_15357_, _15356_, _15354_);
  or (_15358_, _09207_, _08601_);
  and (_15359_, _15358_, _08600_);
  and (_15360_, _15359_, _15357_);
  and (_15361_, _08395_, _08012_);
  and (_15362_, _08738_, \oc8051_golden_model_1.ACC [6]);
  and (_15363_, _08741_, \oc8051_golden_model_1.B [6]);
  or (_15364_, _15363_, _15362_);
  and (_15365_, _08734_, \oc8051_golden_model_1.PSW [6]);
  or (_15366_, _15365_, _15364_);
  and (_15367_, _08752_, \oc8051_golden_model_1.SBUF [6]);
  and (_15368_, _08749_, \oc8051_golden_model_1.IE [6]);
  or (_15369_, _15368_, _15367_);
  and (_15370_, _08746_, \oc8051_golden_model_1.IP [6]);
  or (_15371_, _15370_, _15369_);
  or (_15372_, _15371_, _15366_);
  and (_15373_, _08724_, \oc8051_golden_model_1.TL1 [6]);
  and (_15374_, _08706_, \oc8051_golden_model_1.TH0 [6]);
  and (_15375_, _08710_, \oc8051_golden_model_1.TH1 [6]);
  and (_15376_, _08718_, \oc8051_golden_model_1.SCON [6]);
  or (_15377_, _15376_, _15375_);
  or (_15378_, _15377_, _15374_);
  or (_15379_, _15378_, _15373_);
  or (_15380_, _15379_, _15372_);
  and (_15381_, _08765_, \oc8051_golden_model_1.DPL [6]);
  and (_15382_, _08758_, \oc8051_golden_model_1.SP [6]);
  and (_15383_, _08760_, \oc8051_golden_model_1.DPH [6]);
  or (_15384_, _15383_, _15382_);
  or (_15385_, _15384_, _15381_);
  and (_15386_, _08773_, \oc8051_golden_model_1.TL0 [6]);
  and (_15387_, _08775_, \oc8051_golden_model_1.TMOD [6]);
  or (_15388_, _15387_, _15386_);
  and (_15389_, _08770_, \oc8051_golden_model_1.PCON [6]);
  and (_15390_, _08726_, \oc8051_golden_model_1.TCON [6]);
  or (_15391_, _15390_, _15389_);
  or (_15392_, _15391_, _15388_);
  or (_15393_, _15392_, _15385_);
  or (_15394_, _15393_, _15380_);
  or (_15395_, _15394_, _15361_);
  and (_15396_, _15395_, _08599_);
  or (_15397_, _15396_, _08788_);
  or (_15398_, _15397_, _15360_);
  and (_15399_, _08788_, _06203_);
  nor (_15400_, _15399_, _06112_);
  and (_15401_, _15400_, _15398_);
  not (_15402_, _08638_);
  and (_15403_, _15402_, _06112_);
  or (_15404_, _15403_, _06076_);
  or (_15405_, _15404_, _15401_);
  or (_15406_, _12180_, _05836_);
  and (_15407_, _15406_, _15405_);
  or (_15408_, _15407_, _07128_);
  not (_15409_, _07128_);
  nand (_15410_, _08638_, _08014_);
  nor (_15411_, _08638_, _08014_);
  not (_15412_, _15411_);
  and (_15413_, _15412_, _15410_);
  or (_15414_, _15413_, _15409_);
  and (_15415_, _15414_, _08807_);
  and (_15416_, _15415_, _15408_);
  or (_15417_, _15416_, _15295_);
  and (_15418_, _15417_, _08806_);
  and (_15419_, _15411_, _07133_);
  or (_15420_, _15419_, _15418_);
  and (_15421_, _15420_, _08364_);
  and (_15422_, _10266_, _07131_);
  or (_15423_, _15422_, _07124_);
  or (_15424_, _15423_, _15421_);
  nor (_15425_, _12180_, _05848_);
  nor (_15426_, _15425_, _08820_);
  and (_15427_, _15426_, _15424_);
  and (_15428_, _15410_, _08820_);
  or (_15429_, _15428_, _08825_);
  or (_15430_, _15429_, _15427_);
  nand (_15431_, _10294_, _08825_);
  and (_15432_, _15431_, _05846_);
  and (_15433_, _15432_, _15430_);
  or (_15434_, _15433_, _15294_);
  and (_15435_, _15434_, _08361_);
  nor (_15436_, _15304_, _08361_);
  or (_15437_, _15436_, _07325_);
  nor (_15438_, _15437_, _15435_);
  and (_15439_, _15304_, _07325_);
  or (_15440_, _15439_, _14487_);
  nor (_15441_, _15440_, _15438_);
  nor (_15442_, _09165_, _08883_);
  nor (_15443_, _15442_, _09166_);
  nand (_15444_, _15443_, _06276_);
  and (_15445_, _15444_, _07153_);
  or (_15446_, _15445_, _15441_);
  nand (_15447_, _15443_, _14495_);
  and (_15448_, _15447_, _08837_);
  and (_15449_, _15448_, _15446_);
  and (_15450_, _15300_, _07152_);
  or (_15451_, _15450_, _06310_);
  or (_15452_, _15451_, _15449_);
  nand (_15453_, _12006_, _06310_);
  and (_15454_, _15453_, _12730_);
  and (_15455_, _15454_, _15452_);
  and (_15456_, _12180_, _05823_);
  or (_15457_, _15456_, _06073_);
  or (_15458_, _15457_, _15455_);
  and (_15459_, _06539_, _07369_);
  nor (_15460_, _15297_, _06074_);
  nor (_15461_, _15460_, _15459_);
  and (_15462_, _15461_, _15458_);
  nor (_15463_, _09199_, _08012_);
  nor (_15464_, _15463_, _09200_);
  and (_15465_, _15464_, _15459_);
  or (_15466_, _15465_, _15462_);
  or (_15467_, _15466_, _15293_);
  not (_15468_, _15293_);
  nor (_15469_, _15464_, _15468_);
  nor (_15470_, _15469_, _07394_);
  and (_15471_, _15470_, _15467_);
  and (_15472_, _15464_, _07394_);
  or (_15473_, _15472_, _07168_);
  or (_15474_, _15473_, _15471_);
  and (_15475_, _15474_, _15291_);
  or (_15476_, _15475_, _07167_);
  nor (_15477_, _08341_, _08015_);
  nor (_15478_, _15477_, _08342_);
  or (_15479_, _15478_, _14518_);
  and (_15480_, _15479_, _07417_);
  and (_15481_, _15480_, _15476_);
  or (_15482_, _15481_, _14164_);
  and (_15483_, _15482_, _15288_);
  nand (_15484_, _11966_, _06310_);
  or (_15485_, _12146_, _06310_);
  and (_15486_, _15485_, _15484_);
  and (_15487_, _15486_, _07764_);
  and (_15488_, _15487_, _14328_);
  or (_41021_, _15488_, _15483_);
  or (_15489_, _14156_, \oc8051_golden_model_1.IRAM[0] [7]);
  nand (_15490_, _14156_, _09225_);
  and (_15491_, _15490_, _15489_);
  or (_15492_, _15491_, _14161_);
  or (_15493_, _14162_, _09258_);
  and (_41022_, _15493_, _15492_);
  and (_15494_, _14153_, _07345_);
  and (_15495_, _15494_, _14152_);
  not (_15496_, _15495_);
  or (_15497_, _15496_, _14324_);
  or (_15498_, _15495_, \oc8051_golden_model_1.IRAM[1] [0]);
  not (_15499_, _07764_);
  nand (_15500_, _14159_, _07476_);
  or (_15501_, _15500_, _15499_);
  and (_15502_, _15501_, _15498_);
  and (_15503_, _15502_, _15497_);
  and (_15504_, _07764_, _07476_);
  and (_15505_, _15504_, _14159_);
  and (_15506_, _15505_, _14332_);
  or (_41027_, _15506_, _15503_);
  or (_15507_, _15496_, _14521_);
  or (_15508_, _15495_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_15509_, _15508_, _15501_);
  and (_15510_, _15509_, _15507_);
  and (_15511_, _15505_, _14527_);
  or (_41028_, _15511_, _15510_);
  or (_15512_, _15496_, _14713_);
  or (_15513_, _15495_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_15514_, _15513_, _15501_);
  and (_15515_, _15514_, _15512_);
  and (_15516_, _15505_, _14719_);
  or (_41029_, _15516_, _15515_);
  or (_15517_, _15496_, _14900_);
  or (_15518_, _15495_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_15519_, _15518_, _15501_);
  and (_15520_, _15519_, _15517_);
  and (_15521_, _15505_, _14906_);
  or (_41030_, _15521_, _15520_);
  or (_15522_, _15496_, _15090_);
  or (_15523_, _15495_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_15524_, _15523_, _15501_);
  and (_15525_, _15524_, _15522_);
  and (_15526_, _15505_, _15097_);
  or (_41031_, _15526_, _15525_);
  or (_15527_, _15496_, _15278_);
  or (_15528_, _15495_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_15529_, _15528_, _15501_);
  and (_15530_, _15529_, _15527_);
  and (_15531_, _15505_, _15285_);
  or (_41033_, _15531_, _15530_);
  or (_15532_, _15496_, _15481_);
  or (_15533_, _15495_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_15534_, _15533_, _15501_);
  and (_15535_, _15534_, _15532_);
  and (_15536_, _15505_, _15487_);
  or (_41034_, _15536_, _15535_);
  or (_15537_, _15496_, _09226_);
  or (_15538_, _15495_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_15539_, _15538_, _15501_);
  and (_15540_, _15539_, _15537_);
  and (_15541_, _15505_, _09259_);
  or (_41035_, _15541_, _15540_);
  and (_15542_, _07419_, _07174_);
  and (_15543_, _15542_, _14152_);
  not (_15544_, _15543_);
  or (_15545_, _15544_, _14324_);
  or (_15546_, _15543_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand (_15547_, _14159_, _08449_);
  or (_15548_, _15547_, _15499_);
  and (_15549_, _15548_, _15546_);
  and (_15550_, _15549_, _15545_);
  and (_15551_, _08449_, _07764_);
  and (_15552_, _15551_, _14159_);
  and (_15553_, _15552_, _14332_);
  or (_41038_, _15553_, _15550_);
  or (_15554_, _15544_, _14521_);
  or (_15555_, _15543_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_15556_, _15555_, _15548_);
  and (_15557_, _15556_, _15554_);
  and (_15558_, _15552_, _14527_);
  or (_41041_, _15558_, _15557_);
  or (_15559_, _15544_, _14713_);
  or (_15560_, _15543_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_15561_, _15560_, _15548_);
  and (_15562_, _15561_, _15559_);
  and (_15563_, _15552_, _14719_);
  or (_41042_, _15563_, _15562_);
  or (_15564_, _15544_, _14900_);
  or (_15565_, _15543_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_15566_, _15565_, _15548_);
  and (_15567_, _15566_, _15564_);
  and (_15568_, _15552_, _14906_);
  or (_41043_, _15568_, _15567_);
  or (_15569_, _15544_, _15090_);
  or (_15570_, _15543_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_15571_, _15570_, _15548_);
  and (_15572_, _15571_, _15569_);
  and (_15573_, _15552_, _15097_);
  or (_41044_, _15573_, _15572_);
  or (_15574_, _15544_, _15278_);
  or (_15575_, _15543_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_15576_, _15575_, _15548_);
  and (_15577_, _15576_, _15574_);
  and (_15578_, _15552_, _15285_);
  or (_41045_, _15578_, _15577_);
  or (_15579_, _15544_, _15481_);
  or (_15580_, _15543_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_15581_, _15580_, _15548_);
  and (_15582_, _15581_, _15579_);
  and (_15583_, _15552_, _15487_);
  or (_41047_, _15583_, _15582_);
  and (_15584_, _15543_, _09226_);
  or (_15585_, _15543_, _07871_);
  nand (_15586_, _15585_, _15548_);
  or (_15587_, _15586_, _15584_);
  or (_15588_, _15548_, _09258_);
  and (_41048_, _15588_, _15587_);
  and (_15589_, _14152_, _07421_);
  or (_15590_, _15589_, \oc8051_golden_model_1.IRAM[3] [0]);
  nand (_15591_, _14159_, _07177_);
  or (_15592_, _15591_, _15499_);
  and (_15593_, _15592_, _15590_);
  not (_15594_, _15589_);
  or (_15595_, _15594_, _14324_);
  and (_15596_, _15595_, _15593_);
  and (_15597_, _07764_, _07177_);
  and (_15598_, _15597_, _14159_);
  and (_15599_, _15598_, _14332_);
  or (_41052_, _15599_, _15596_);
  or (_15600_, _15589_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_15601_, _15600_, _15592_);
  or (_15602_, _15594_, _14521_);
  and (_15603_, _15602_, _15601_);
  and (_15604_, _15598_, _14527_);
  or (_41053_, _15604_, _15603_);
  or (_15605_, _15589_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_15606_, _15605_, _15592_);
  or (_15607_, _15594_, _14713_);
  and (_15608_, _15607_, _15606_);
  and (_15609_, _15598_, _14719_);
  or (_41054_, _15609_, _15608_);
  or (_15610_, _15589_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_15611_, _15610_, _15592_);
  or (_15612_, _15594_, _14900_);
  and (_15613_, _15612_, _15611_);
  and (_15614_, _15598_, _14906_);
  or (_41055_, _15614_, _15613_);
  or (_15615_, _15589_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_15616_, _15615_, _15592_);
  or (_15617_, _15594_, _15090_);
  and (_15618_, _15617_, _15616_);
  and (_15619_, _15598_, _15097_);
  or (_41056_, _15619_, _15618_);
  or (_15620_, _15589_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_15621_, _15620_, _15592_);
  or (_15622_, _15594_, _15278_);
  and (_15623_, _15622_, _15621_);
  and (_15624_, _15598_, _15285_);
  or (_41058_, _15624_, _15623_);
  or (_15625_, _15589_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_15626_, _15625_, _15592_);
  or (_15627_, _15594_, _15481_);
  and (_15628_, _15627_, _15626_);
  and (_15629_, _15598_, _15487_);
  or (_41059_, _15629_, _15628_);
  or (_15630_, _15589_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_15631_, _15630_, _15592_);
  or (_15632_, _15594_, _09226_);
  and (_15633_, _15632_, _15631_);
  and (_15634_, _15598_, _09259_);
  or (_41060_, _15634_, _15633_);
  and (_15635_, _07747_, _07593_);
  and (_15636_, _15635_, _14154_);
  not (_15637_, _15636_);
  or (_15638_, _15637_, _14324_);
  not (_15639_, _07759_);
  and (_15640_, _14158_, _15639_);
  and (_15641_, _15640_, _07178_);
  not (_15642_, _15641_);
  or (_15643_, _15636_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_15644_, _15643_, _15642_);
  and (_15645_, _15644_, _15638_);
  and (_15646_, _15641_, _14332_);
  or (_41063_, _15646_, _15645_);
  or (_15647_, _15637_, _14521_);
  or (_15648_, _15636_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_15649_, _15648_, _15642_);
  and (_15650_, _15649_, _15647_);
  and (_15651_, _15641_, _14527_);
  or (_41066_, _15651_, _15650_);
  or (_15652_, _15637_, _14713_);
  or (_15653_, _15636_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_15654_, _15653_, _15642_);
  and (_15655_, _15654_, _15652_);
  and (_15656_, _15641_, _14719_);
  or (_41067_, _15656_, _15655_);
  or (_15657_, _15637_, _14900_);
  or (_15658_, _15636_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_15659_, _15658_, _15642_);
  and (_15660_, _15659_, _15657_);
  and (_15661_, _15641_, _14906_);
  or (_41068_, _15661_, _15660_);
  or (_15662_, _15637_, _15090_);
  or (_15663_, _15636_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_15664_, _15663_, _15642_);
  and (_15665_, _15664_, _15662_);
  and (_15666_, _15641_, _15097_);
  or (_41069_, _15666_, _15665_);
  or (_15667_, _15637_, _15278_);
  or (_15668_, _15636_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_15669_, _15668_, _15642_);
  and (_15670_, _15669_, _15667_);
  and (_15671_, _15641_, _15285_);
  or (_41070_, _15671_, _15670_);
  or (_15672_, _15637_, _15481_);
  or (_15673_, _15636_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_15674_, _15673_, _15642_);
  and (_15675_, _15674_, _15672_);
  and (_15676_, _15641_, _15487_);
  or (_41071_, _15676_, _15675_);
  or (_15677_, _15637_, _09226_);
  or (_15678_, _15636_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_15679_, _15678_, _15642_);
  and (_15680_, _15679_, _15677_);
  and (_15681_, _15641_, _09259_);
  or (_41072_, _15681_, _15680_);
  and (_15682_, _15635_, _15494_);
  not (_15683_, _15682_);
  or (_15684_, _15683_, _14324_);
  and (_15685_, _15640_, _07476_);
  not (_15686_, _15685_);
  or (_15687_, _15682_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_15688_, _15687_, _15686_);
  and (_15689_, _15688_, _15684_);
  and (_15690_, _15685_, _14332_);
  or (_41075_, _15690_, _15689_);
  or (_15691_, _15683_, _14521_);
  or (_15692_, _15682_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_15693_, _15692_, _15686_);
  and (_15694_, _15693_, _15691_);
  and (_15695_, _15685_, _14527_);
  or (_41077_, _15695_, _15694_);
  or (_15696_, _15683_, _14713_);
  or (_15697_, _15682_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_15698_, _15697_, _15686_);
  and (_15699_, _15698_, _15696_);
  and (_15700_, _15685_, _14719_);
  or (_41078_, _15700_, _15699_);
  or (_15701_, _15683_, _14900_);
  or (_15702_, _15682_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_15703_, _15702_, _15686_);
  and (_15704_, _15703_, _15701_);
  and (_15705_, _15685_, _14906_);
  or (_41079_, _15705_, _15704_);
  or (_15706_, _15683_, _15090_);
  or (_15707_, _15682_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_15708_, _15707_, _15686_);
  and (_15709_, _15708_, _15706_);
  and (_15710_, _15685_, _15097_);
  or (_41080_, _15710_, _15709_);
  or (_15711_, _15683_, _15278_);
  or (_15712_, _15682_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_15713_, _15712_, _15686_);
  and (_15714_, _15713_, _15711_);
  and (_15715_, _15685_, _15285_);
  or (_41081_, _15715_, _15714_);
  or (_15716_, _15683_, _15481_);
  or (_15717_, _15682_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_15718_, _15717_, _15686_);
  and (_15719_, _15718_, _15716_);
  and (_15720_, _15685_, _15487_);
  or (_41083_, _15720_, _15719_);
  or (_15721_, _15683_, _09226_);
  or (_15722_, _15682_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_15723_, _15722_, _15686_);
  and (_15724_, _15723_, _15721_);
  and (_15725_, _15685_, _09259_);
  or (_41084_, _15725_, _15724_);
  and (_15726_, _15635_, _15542_);
  not (_15727_, _15726_);
  or (_15728_, _15727_, _14324_);
  and (_15729_, _15640_, _08449_);
  not (_15730_, _15729_);
  or (_15731_, _15726_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_15732_, _15731_, _15730_);
  and (_15733_, _15732_, _15728_);
  and (_15734_, _15729_, _14332_);
  or (_41088_, _15734_, _15733_);
  or (_15735_, _15727_, _14521_);
  or (_15736_, _15726_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_15737_, _15736_, _15730_);
  and (_15738_, _15737_, _15735_);
  and (_15739_, _15729_, _14527_);
  or (_41089_, _15739_, _15738_);
  or (_15740_, _15727_, _14713_);
  or (_15741_, _15726_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_15742_, _15741_, _15730_);
  and (_15743_, _15742_, _15740_);
  and (_15744_, _15729_, _14719_);
  or (_41090_, _15744_, _15743_);
  or (_15745_, _15727_, _14900_);
  or (_15746_, _15726_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_15747_, _15746_, _15730_);
  and (_15748_, _15747_, _15745_);
  and (_15749_, _15729_, _14906_);
  or (_41091_, _15749_, _15748_);
  or (_15750_, _15727_, _15090_);
  or (_15751_, _15726_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_15752_, _15751_, _15730_);
  and (_15753_, _15752_, _15750_);
  and (_15754_, _15729_, _15097_);
  or (_41092_, _15754_, _15753_);
  or (_15755_, _15727_, _15278_);
  or (_15756_, _15726_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_15757_, _15756_, _15730_);
  and (_15758_, _15757_, _15755_);
  and (_15759_, _15729_, _15285_);
  or (_41094_, _15759_, _15758_);
  or (_15760_, _15727_, _15481_);
  or (_15761_, _15726_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_15762_, _15761_, _15730_);
  and (_15763_, _15762_, _15760_);
  and (_15764_, _15729_, _15487_);
  or (_41095_, _15764_, _15763_);
  or (_15765_, _15727_, _09226_);
  or (_15766_, _15726_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_15767_, _15766_, _15730_);
  and (_15768_, _15767_, _15765_);
  and (_15769_, _15729_, _09259_);
  or (_41096_, _15769_, _15768_);
  and (_15770_, _15640_, _07177_);
  not (_15771_, _15770_);
  or (_15772_, _15771_, _14332_);
  and (_15773_, _15635_, _07421_);
  and (_15774_, _15773_, _14324_);
  nor (_15775_, _15773_, _07007_);
  or (_15776_, _15775_, _15770_);
  or (_15777_, _15776_, _15774_);
  and (_41100_, _15777_, _15772_);
  nor (_15778_, _15773_, _07207_);
  and (_15779_, _15773_, _14521_);
  or (_15780_, _15779_, _15778_);
  and (_15781_, _15780_, _15771_);
  and (_15782_, _15770_, _14527_);
  or (_41101_, _15782_, _15781_);
  or (_15783_, _15773_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_15784_, _15783_, _15771_);
  not (_15785_, _15773_);
  or (_15786_, _15785_, _14713_);
  and (_15787_, _15786_, _15784_);
  and (_15788_, _15770_, _14719_);
  or (_41102_, _15788_, _15787_);
  or (_15789_, _15773_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_15790_, _15789_, _15771_);
  or (_15791_, _15785_, _14900_);
  and (_15792_, _15791_, _15790_);
  and (_15793_, _15770_, _14906_);
  or (_41103_, _15793_, _15792_);
  or (_15794_, _15773_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_15795_, _15794_, _15771_);
  or (_15796_, _15785_, _15090_);
  and (_15797_, _15796_, _15795_);
  and (_15798_, _15770_, _15097_);
  or (_41104_, _15798_, _15797_);
  or (_15799_, _15773_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_15800_, _15799_, _15771_);
  or (_15801_, _15785_, _15278_);
  and (_15802_, _15801_, _15800_);
  and (_15803_, _15770_, _15285_);
  or (_41106_, _15803_, _15802_);
  or (_15804_, _15773_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_15805_, _15804_, _15771_);
  or (_15806_, _15785_, _15481_);
  and (_15807_, _15806_, _15805_);
  and (_15808_, _15770_, _15487_);
  or (_41107_, _15808_, _15807_);
  or (_15809_, _15773_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_15810_, _15809_, _15771_);
  or (_15811_, _15785_, _09226_);
  and (_15812_, _15811_, _15810_);
  and (_15813_, _15770_, _09259_);
  or (_41108_, _15813_, _15812_);
  and (_15814_, _14151_, _07746_);
  and (_15815_, _15814_, _14154_);
  not (_15816_, _15815_);
  or (_15817_, _15816_, _14324_);
  or (_15818_, _15815_, \oc8051_golden_model_1.IRAM[8] [0]);
  not (_15819_, _07755_);
  and (_15820_, _07765_, _15819_);
  and (_15821_, _15820_, _07178_);
  not (_15822_, _15821_);
  and (_15823_, _15822_, _15818_);
  and (_15824_, _15823_, _15817_);
  and (_15825_, _15821_, _14332_);
  or (_41112_, _15825_, _15824_);
  or (_15826_, _15816_, _14521_);
  or (_15827_, _15815_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_15828_, _15827_, _15822_);
  and (_15829_, _15828_, _15826_);
  and (_15830_, _15821_, _14527_);
  or (_41114_, _15830_, _15829_);
  or (_15831_, _15816_, _14713_);
  nand (_15832_, _07765_, _07753_);
  or (_15833_, _15815_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_15834_, _15833_, _15832_);
  and (_15835_, _15834_, _15831_);
  and (_15836_, _15821_, _14719_);
  or (_41115_, _15836_, _15835_);
  or (_15837_, _15816_, _14900_);
  or (_15838_, _15815_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_15839_, _15838_, _15832_);
  and (_15840_, _15839_, _15837_);
  and (_15841_, _15821_, _14906_);
  or (_41116_, _15841_, _15840_);
  or (_15842_, _15816_, _15090_);
  or (_15843_, _15815_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_15844_, _15843_, _15832_);
  and (_15845_, _15844_, _15842_);
  and (_15846_, _15821_, _15097_);
  or (_41117_, _15846_, _15845_);
  or (_15847_, _15816_, _15278_);
  or (_15848_, _15815_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_15849_, _15848_, _15832_);
  and (_15850_, _15849_, _15847_);
  and (_15851_, _15821_, _15285_);
  or (_41118_, _15851_, _15850_);
  or (_15852_, _15816_, _15481_);
  or (_15853_, _15815_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_15854_, _15853_, _15832_);
  and (_15855_, _15854_, _15852_);
  and (_15856_, _15821_, _15487_);
  or (_41120_, _15856_, _15855_);
  and (_15857_, _15815_, _09226_);
  or (_15858_, _15815_, _07899_);
  nand (_15859_, _15858_, _15832_);
  or (_15860_, _15859_, _15857_);
  or (_15861_, _15822_, _09259_);
  and (_41121_, _15861_, _15860_);
  and (_15862_, _15814_, _15494_);
  not (_15863_, _15862_);
  or (_15864_, _15863_, _14324_);
  or (_15865_, _15862_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_15866_, _15820_, _07476_);
  not (_15867_, _15866_);
  and (_15868_, _15867_, _15865_);
  and (_15869_, _15868_, _15864_);
  and (_15870_, _15866_, _14332_);
  or (_41123_, _15870_, _15869_);
  or (_15871_, _15863_, _14521_);
  or (_15872_, _15862_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_15873_, _15872_, _15867_);
  and (_15874_, _15873_, _15871_);
  and (_15875_, _15866_, _14527_);
  or (_41124_, _15875_, _15874_);
  or (_15876_, _15863_, _14713_);
  nand (_15877_, _07765_, _07477_);
  or (_15878_, _15862_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_15879_, _15878_, _15877_);
  and (_15880_, _15879_, _15876_);
  and (_15881_, _15866_, _14719_);
  or (_41125_, _15881_, _15880_);
  or (_15882_, _15863_, _14900_);
  or (_15883_, _15862_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_15884_, _15883_, _15877_);
  and (_15885_, _15884_, _15882_);
  and (_15886_, _15866_, _14906_);
  or (_41126_, _15886_, _15885_);
  or (_15887_, _15863_, _15090_);
  or (_15888_, _15862_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_15889_, _15888_, _15877_);
  and (_15890_, _15889_, _15887_);
  and (_15891_, _15866_, _15097_);
  or (_41127_, _15891_, _15890_);
  or (_15892_, _15863_, _15278_);
  or (_15893_, _15862_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_15894_, _15893_, _15877_);
  and (_15895_, _15894_, _15892_);
  and (_15896_, _15866_, _15285_);
  or (_41128_, _15896_, _15895_);
  or (_15897_, _15863_, _15481_);
  or (_15898_, _15862_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_15899_, _15898_, _15877_);
  and (_15900_, _15899_, _15897_);
  and (_15901_, _15866_, _15487_);
  or (_41131_, _15901_, _15900_);
  and (_15902_, _15862_, _09226_);
  or (_15903_, _15862_, _07901_);
  nand (_15904_, _15903_, _15877_);
  or (_15905_, _15904_, _15902_);
  or (_15906_, _15867_, _09259_);
  and (_41132_, _15906_, _15905_);
  and (_15907_, _15814_, _15542_);
  not (_15908_, _15907_);
  or (_15909_, _15908_, _14324_);
  and (_15910_, _15820_, _08449_);
  not (_15911_, _15910_);
  or (_15912_, _15907_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_15913_, _15912_, _15911_);
  and (_15914_, _15913_, _15909_);
  and (_15915_, _15910_, _14332_);
  or (_41136_, _15915_, _15914_);
  or (_15916_, _15908_, _14521_);
  or (_15917_, _15907_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_15918_, _15917_, _15911_);
  and (_15919_, _15918_, _15916_);
  and (_15920_, _15910_, _14527_);
  or (_41137_, _15920_, _15919_);
  or (_15921_, _15908_, _14713_);
  or (_15922_, _15907_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_15923_, _15922_, _15911_);
  and (_15924_, _15923_, _15921_);
  and (_15925_, _15910_, _14719_);
  or (_41138_, _15925_, _15924_);
  or (_15926_, _15908_, _14900_);
  or (_15927_, _15907_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_15928_, _15927_, _15911_);
  and (_15929_, _15928_, _15926_);
  and (_15930_, _15910_, _14906_);
  or (_41139_, _15930_, _15929_);
  or (_15931_, _15908_, _15090_);
  or (_15932_, _15907_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_15933_, _15932_, _15911_);
  and (_15934_, _15933_, _15931_);
  and (_15935_, _15910_, _15097_);
  or (_41140_, _15935_, _15934_);
  or (_15936_, _15908_, _15278_);
  or (_15937_, _15907_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_15938_, _15937_, _15911_);
  and (_15939_, _15938_, _15936_);
  and (_15940_, _15910_, _15285_);
  or (_41142_, _15940_, _15939_);
  or (_15941_, _15908_, _15481_);
  or (_15942_, _15907_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_15943_, _15942_, _15911_);
  and (_15944_, _15943_, _15941_);
  and (_15945_, _15910_, _15487_);
  or (_41143_, _15945_, _15944_);
  or (_15946_, _15908_, _09226_);
  or (_15947_, _15907_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_15948_, _15947_, _15911_);
  and (_15949_, _15948_, _15946_);
  and (_15950_, _15910_, _09259_);
  or (_41144_, _15950_, _15949_);
  not (_15951_, _07345_);
  and (_15952_, _14153_, _15951_);
  and (_15953_, _15814_, _15952_);
  not (_15954_, _15953_);
  or (_15955_, _15954_, _14324_);
  and (_15956_, _15820_, _07177_);
  not (_15957_, _15956_);
  or (_15958_, _15953_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_15959_, _15958_, _15957_);
  and (_15960_, _15959_, _15955_);
  and (_15961_, _15956_, _14332_);
  or (_41148_, _15961_, _15960_);
  or (_15962_, _15954_, _14521_);
  or (_15963_, _15953_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_15964_, _15963_, _15957_);
  and (_15965_, _15964_, _15962_);
  and (_15966_, _15956_, _14527_);
  or (_41149_, _15966_, _15965_);
  or (_15967_, _15954_, _14713_);
  or (_15968_, _15953_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_15969_, _15968_, _15957_);
  and (_15970_, _15969_, _15967_);
  and (_15971_, _15956_, _14719_);
  or (_41150_, _15971_, _15970_);
  and (_15972_, _15814_, _07421_);
  or (_15973_, _15972_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_15974_, _15973_, _15957_);
  not (_15975_, _15972_);
  or (_15976_, _15975_, _14900_);
  and (_15977_, _15976_, _15974_);
  and (_15978_, _15956_, _14906_);
  or (_41151_, _15978_, _15977_);
  or (_15979_, _15972_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_15980_, _15979_, _15957_);
  or (_15981_, _15975_, _15090_);
  and (_15982_, _15981_, _15980_);
  and (_15983_, _15956_, _15097_);
  or (_41152_, _15983_, _15982_);
  or (_15984_, _15972_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_15985_, _15984_, _15957_);
  or (_15986_, _15975_, _15278_);
  and (_15987_, _15986_, _15985_);
  and (_15988_, _15956_, _15285_);
  or (_41153_, _15988_, _15987_);
  or (_15989_, _15972_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_15990_, _15989_, _15957_);
  or (_15991_, _15975_, _15481_);
  and (_15992_, _15991_, _15990_);
  and (_15993_, _15956_, _15487_);
  or (_41154_, _15993_, _15992_);
  or (_15994_, _15972_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_15995_, _15994_, _15957_);
  or (_15996_, _15975_, _09226_);
  and (_15997_, _15996_, _15995_);
  and (_15998_, _15956_, _09259_);
  or (_41155_, _15998_, _15997_);
  not (_15999_, _07178_);
  nand (_16000_, _14158_, _07759_);
  or (_16001_, _16000_, _15999_);
  or (_16002_, _16001_, _14332_);
  and (_16003_, _14154_, _07749_);
  and (_16004_, _16003_, _14324_);
  or (_16005_, _16003_, _07039_);
  nand (_16006_, _16005_, _16001_);
  or (_16007_, _16006_, _16004_);
  and (_41158_, _16007_, _16002_);
  not (_16008_, _07746_);
  and (_16009_, _14151_, _16008_);
  and (_16010_, _14154_, _16009_);
  not (_16011_, _16010_);
  or (_16012_, _16011_, _14521_);
  and (_16013_, _07766_, _07178_);
  not (_16014_, _16013_);
  or (_16015_, _16010_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_16016_, _16015_, _16014_);
  and (_16017_, _16016_, _16012_);
  and (_16018_, _16013_, _14527_);
  or (_41159_, _16018_, _16017_);
  or (_16019_, _16003_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_16020_, _16019_, _16014_);
  or (_16021_, _16011_, _14713_);
  and (_16022_, _16021_, _16020_);
  and (_16023_, _16013_, _14719_);
  or (_41160_, _16023_, _16022_);
  or (_16024_, _16003_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_16025_, _16024_, _16014_);
  or (_16026_, _16011_, _14900_);
  and (_16027_, _16026_, _16025_);
  and (_16028_, _16013_, _14906_);
  or (_41162_, _16028_, _16027_);
  or (_16029_, _16003_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_16030_, _16029_, _16014_);
  or (_16031_, _16011_, _15090_);
  and (_16032_, _16031_, _16030_);
  and (_16033_, _16013_, _15097_);
  or (_41163_, _16033_, _16032_);
  or (_16034_, _16011_, _15278_);
  or (_16035_, _16003_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_16036_, _16035_, _16014_);
  and (_16037_, _16036_, _16034_);
  and (_16038_, _16013_, _15285_);
  or (_41164_, _16038_, _16037_);
  or (_16039_, _16003_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_16040_, _16039_, _16014_);
  or (_16041_, _16011_, _15481_);
  and (_16042_, _16041_, _16040_);
  and (_16043_, _16013_, _15487_);
  or (_41165_, _16043_, _16042_);
  and (_16044_, _16003_, _09226_);
  or (_16045_, _16003_, _07913_);
  nand (_16046_, _16045_, _16001_);
  or (_16047_, _16046_, _16044_);
  or (_16048_, _16014_, _09259_);
  and (_41166_, _16048_, _16047_);
  and (_16049_, _07766_, _07476_);
  not (_16050_, _16049_);
  or (_16051_, _16050_, _14332_);
  and (_16052_, _15494_, _07749_);
  and (_16053_, _16052_, _14324_);
  nor (_16054_, _16052_, _07041_);
  or (_16055_, _16054_, _16049_);
  or (_16056_, _16055_, _16053_);
  and (_41169_, _16056_, _16051_);
  and (_16057_, _15494_, _16009_);
  not (_16058_, _16057_);
  or (_16059_, _16058_, _14521_);
  or (_16060_, _16057_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_16061_, _16060_, _16050_);
  and (_16062_, _16061_, _16059_);
  and (_16063_, _16049_, _14527_);
  or (_41170_, _16063_, _16062_);
  or (_16064_, _16052_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_16065_, _16064_, _16050_);
  or (_16066_, _16058_, _14713_);
  and (_16067_, _16066_, _16065_);
  and (_16068_, _16049_, _14719_);
  or (_41171_, _16068_, _16067_);
  or (_16069_, _16052_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_16070_, _16069_, _16050_);
  or (_16071_, _16058_, _14900_);
  and (_16072_, _16071_, _16070_);
  and (_16073_, _16049_, _14906_);
  or (_41173_, _16073_, _16072_);
  or (_16074_, _16052_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_16075_, _16074_, _16050_);
  or (_16076_, _16058_, _15090_);
  and (_16077_, _16076_, _16075_);
  and (_16078_, _16049_, _15097_);
  or (_41174_, _16078_, _16077_);
  and (_16079_, _16049_, _15285_);
  or (_16080_, _16052_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_16081_, _16080_, _16050_);
  or (_16082_, _16058_, _15278_);
  and (_16083_, _16082_, _16081_);
  or (_41175_, _16083_, _16079_);
  or (_16084_, _16058_, _15481_);
  or (_16085_, _16052_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_16086_, _16085_, _16050_);
  and (_16087_, _16086_, _16084_);
  and (_16088_, _16049_, _15487_);
  or (_41176_, _16088_, _16087_);
  and (_16089_, _16049_, _09259_);
  or (_16090_, _16052_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_16091_, _16090_, _16050_);
  or (_16092_, _16058_, _09226_);
  and (_16093_, _16092_, _16091_);
  or (_41177_, _16093_, _16089_);
  and (_16094_, _15542_, _16009_);
  not (_16095_, _16094_);
  or (_16096_, _16095_, _14324_);
  and (_16097_, _15542_, _07749_);
  or (_16098_, _16097_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_16099_, _08449_, _07766_);
  not (_16100_, _16099_);
  and (_16101_, _16100_, _16098_);
  and (_16102_, _16101_, _16096_);
  and (_16103_, _16099_, _14332_);
  or (_41181_, _16103_, _16102_);
  or (_16104_, _16095_, _14521_);
  or (_16105_, _16094_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_16106_, _16105_, _16100_);
  and (_16107_, _16106_, _16104_);
  and (_16108_, _16099_, _14527_);
  or (_41182_, _16108_, _16107_);
  or (_16109_, _16097_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_16110_, _16109_, _16100_);
  or (_16111_, _16095_, _14713_);
  and (_16112_, _16111_, _16110_);
  and (_16113_, _16099_, _14719_);
  or (_41184_, _16113_, _16112_);
  or (_16114_, _16097_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_16115_, _16114_, _16100_);
  or (_16116_, _16095_, _14900_);
  and (_16117_, _16116_, _16115_);
  and (_16118_, _16099_, _14906_);
  or (_41185_, _16118_, _16117_);
  or (_16119_, _16095_, _15090_);
  or (_16120_, _16097_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_16121_, _16120_, _16100_);
  and (_16122_, _16121_, _16119_);
  and (_16123_, _16099_, _15097_);
  or (_41186_, _16123_, _16122_);
  or (_16124_, _16097_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_16125_, _16124_, _16100_);
  or (_16126_, _16095_, _15278_);
  and (_16127_, _16126_, _16125_);
  and (_16128_, _16099_, _15285_);
  or (_41187_, _16128_, _16127_);
  or (_16129_, _16097_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_16130_, _16129_, _16100_);
  or (_16131_, _16095_, _15481_);
  and (_16132_, _16131_, _16130_);
  and (_16133_, _16099_, _15487_);
  or (_41188_, _16133_, _16132_);
  nor (_16134_, _16094_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_16135_, _16095_, _09226_);
  or (_16136_, _16135_, _16134_);
  nand (_16137_, _16136_, _16100_);
  or (_16138_, _16100_, _09259_);
  and (_41190_, _16138_, _16137_);
  not (_16139_, _07177_);
  or (_16140_, _16000_, _16139_);
  or (_16141_, _14332_, _16140_);
  and (_16142_, _14324_, _07750_);
  or (_16143_, _07750_, _07034_);
  nand (_16144_, _16143_, _16140_);
  or (_16145_, _16144_, _16142_);
  and (_41193_, _16145_, _16141_);
  nor (_16146_, _07750_, _07237_);
  and (_16147_, _14521_, _07750_);
  or (_16148_, _16147_, _16146_);
  and (_16149_, _16148_, _16140_);
  and (_16150_, _14527_, _07767_);
  or (_41194_, _16150_, _16149_);
  or (_16151_, _07750_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_16152_, _16151_, _07768_);
  or (_16153_, _14713_, _07770_);
  and (_16154_, _16153_, _16152_);
  and (_16155_, _14719_, _07767_);
  or (_41196_, _16155_, _16154_);
  or (_16156_, _07750_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_16157_, _16156_, _07768_);
  or (_16158_, _14900_, _07770_);
  and (_16159_, _16158_, _16157_);
  and (_16160_, _14906_, _07767_);
  or (_41197_, _16160_, _16159_);
  or (_16161_, _07750_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_16162_, _16161_, _07768_);
  or (_16163_, _15090_, _07770_);
  and (_16164_, _16163_, _16162_);
  and (_16165_, _15097_, _07767_);
  or (_41198_, _16165_, _16164_);
  or (_16166_, _07750_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_16167_, _16166_, _07768_);
  or (_16168_, _15278_, _07770_);
  and (_16169_, _16168_, _16167_);
  and (_16170_, _15285_, _07767_);
  or (_41199_, _16170_, _16169_);
  or (_16171_, _07750_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_16172_, _16171_, _07768_);
  or (_16173_, _15481_, _07770_);
  and (_16174_, _16173_, _16172_);
  and (_16175_, _15487_, _07767_);
  or (_41200_, _16175_, _16174_);
  nor (_16176_, _01317_, _09899_);
  nor (_16177_, _07841_, _09899_);
  and (_16178_, _07841_, _07049_);
  or (_16179_, _16178_, _16177_);
  or (_16180_, _16179_, _07075_);
  nor (_16181_, _08211_, _10243_);
  or (_16182_, _16181_, _16177_);
  or (_16183_, _16182_, _06161_);
  and (_16184_, _07841_, \oc8051_golden_model_1.ACC [0]);
  or (_16185_, _16184_, _16177_);
  and (_16186_, _16185_, _07056_);
  nor (_16187_, _07056_, _09899_);
  or (_16188_, _16187_, _06160_);
  or (_16189_, _16188_, _16186_);
  and (_16190_, _16189_, _06157_);
  and (_16191_, _16190_, _16183_);
  nor (_16192_, _08420_, _09899_);
  and (_16193_, _14169_, _08420_);
  or (_16194_, _16193_, _16192_);
  and (_16195_, _16194_, _06156_);
  or (_16196_, _16195_, _16191_);
  or (_16197_, _16196_, _06217_);
  and (_16198_, _16197_, _16180_);
  or (_16199_, _16198_, _06220_);
  or (_16200_, _16185_, _06229_);
  and (_16201_, _16200_, _06153_);
  and (_16202_, _16201_, _16199_);
  and (_16203_, _16177_, _06152_);
  or (_16204_, _16203_, _06145_);
  or (_16205_, _16204_, _16202_);
  or (_16206_, _16182_, _06146_);
  and (_16207_, _16206_, _16205_);
  or (_16208_, _16207_, _09295_);
  nor (_16209_, _09793_, _09790_);
  nor (_16210_, _16209_, _09795_);
  or (_16211_, _16210_, _09301_);
  and (_16212_, _16211_, _06140_);
  and (_16213_, _16212_, _16208_);
  or (_16214_, _16192_, _14170_);
  and (_16215_, _16214_, _06139_);
  and (_16216_, _16215_, _16194_);
  or (_16217_, _16216_, _09842_);
  or (_16218_, _16217_, _16213_);
  or (_16219_, _16179_, _06132_);
  and (_16220_, _16219_, _06117_);
  and (_16221_, _16220_, _16218_);
  and (_16222_, _09160_, _07841_);
  or (_16223_, _16222_, _16177_);
  and (_16224_, _16223_, _06116_);
  or (_16225_, _16224_, _05787_);
  or (_16226_, _16225_, _16221_);
  and (_16227_, _14260_, _07841_);
  or (_16228_, _16177_, _06114_);
  or (_16229_, _16228_, _16227_);
  and (_16230_, _16229_, _09861_);
  and (_16231_, _16230_, _16226_);
  nand (_16232_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  or (_16233_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_16234_, _16233_, _16232_);
  or (_16235_, _10209_, _16234_);
  nand (_16236_, _10209_, _05855_);
  and (_16237_, _16236_, _09855_);
  and (_16238_, _16237_, _16235_);
  or (_16239_, _16238_, _11136_);
  or (_16240_, _16239_, _16231_);
  and (_16241_, _14275_, _07841_);
  or (_16242_, _16177_, _07127_);
  or (_16243_, _16242_, _16241_);
  and (_16244_, _07841_, _08708_);
  or (_16245_, _16244_, _16177_);
  or (_16246_, _16245_, _06111_);
  and (_16247_, _16246_, _07125_);
  and (_16248_, _16247_, _16243_);
  and (_16249_, _16248_, _16240_);
  nor (_16250_, _12321_, _10243_);
  or (_16251_, _16250_, _16177_);
  nand (_16252_, _10276_, _07841_);
  and (_16253_, _16252_, _06402_);
  and (_16254_, _16253_, _16251_);
  or (_16255_, _16254_, _16249_);
  and (_16256_, _16255_, _07132_);
  nand (_16257_, _16245_, _06306_);
  nor (_16258_, _16257_, _16181_);
  or (_16259_, _16258_, _06411_);
  or (_16260_, _16259_, _16256_);
  nor (_16261_, _16177_, _07130_);
  nand (_16262_, _16261_, _16252_);
  and (_16263_, _16262_, _16260_);
  or (_16264_, _16263_, _06303_);
  and (_16265_, _14167_, _07841_);
  or (_16266_, _16177_, _08819_);
  or (_16267_, _16266_, _16265_);
  and (_16268_, _16267_, _08824_);
  and (_16269_, _16268_, _16264_);
  and (_16270_, _16251_, _06396_);
  or (_16271_, _16270_, _06433_);
  or (_16272_, _16271_, _16269_);
  or (_16273_, _16182_, _06829_);
  and (_16274_, _16273_, _16272_);
  or (_16275_, _16274_, _05748_);
  or (_16276_, _16177_, _05749_);
  and (_16277_, _16276_, _16275_);
  or (_16278_, _16277_, _06440_);
  or (_16279_, _16182_, _06444_);
  and (_16280_, _16279_, _01317_);
  and (_16281_, _16280_, _16278_);
  or (_16282_, _16281_, _16176_);
  and (_43594_, _16282_, _43100_);
  nor (_16283_, _01317_, _09864_);
  nor (_16284_, _07841_, _09864_);
  nor (_16285_, _10277_, _10243_);
  or (_16286_, _16285_, _16284_);
  or (_16287_, _16286_, _08824_);
  nor (_16288_, _08420_, _09864_);
  and (_16289_, _14349_, _08420_);
  or (_16290_, _16289_, _16288_);
  and (_16291_, _16290_, _06152_);
  and (_16292_, _07841_, _07306_);
  or (_16293_, _16292_, _16284_);
  or (_16294_, _16293_, _07075_);
  or (_16295_, _07841_, \oc8051_golden_model_1.B [1]);
  and (_16296_, _14363_, _07841_);
  not (_16297_, _16296_);
  and (_16298_, _16297_, _16295_);
  or (_16299_, _16298_, _06161_);
  and (_16300_, _07841_, \oc8051_golden_model_1.ACC [1]);
  or (_16301_, _16300_, _16284_);
  and (_16302_, _16301_, _07056_);
  nor (_16303_, _07056_, _09864_);
  or (_16304_, _16303_, _06160_);
  or (_16305_, _16304_, _16302_);
  and (_16306_, _16305_, _06157_);
  and (_16307_, _16306_, _16299_);
  and (_16308_, _14367_, _08420_);
  or (_16309_, _16308_, _16288_);
  and (_16310_, _16309_, _06156_);
  or (_16311_, _16310_, _06217_);
  or (_16312_, _16311_, _16307_);
  and (_16313_, _16312_, _16294_);
  or (_16314_, _16313_, _06220_);
  or (_16315_, _16301_, _06229_);
  and (_16316_, _16315_, _06153_);
  and (_16317_, _16316_, _16314_);
  or (_16318_, _16317_, _16291_);
  and (_16319_, _16318_, _06146_);
  and (_16320_, _16308_, _14382_);
  or (_16321_, _16320_, _16288_);
  and (_16322_, _16321_, _06145_);
  or (_16323_, _16322_, _09295_);
  or (_16324_, _16323_, _16319_);
  nor (_16325_, _09798_, _09737_);
  nor (_16326_, _16325_, _09799_);
  or (_16327_, _16326_, _09301_);
  and (_16328_, _16327_, _06140_);
  and (_16329_, _16328_, _16324_);
  and (_16330_, _14351_, _08420_);
  or (_16331_, _16330_, _16288_);
  and (_16332_, _16331_, _06139_);
  or (_16333_, _16332_, _09842_);
  or (_16334_, _16333_, _16329_);
  or (_16335_, _16293_, _06132_);
  and (_16336_, _16335_, _16334_);
  or (_16337_, _16336_, _06116_);
  and (_16338_, _09115_, _07841_);
  or (_16339_, _16284_, _06117_);
  or (_16340_, _16339_, _16338_);
  and (_16341_, _16340_, _06114_);
  and (_16342_, _16341_, _16337_);
  or (_16343_, _14442_, _10243_);
  and (_16344_, _16295_, _05787_);
  and (_16345_, _16344_, _16343_);
  or (_16346_, _16345_, _09855_);
  or (_16347_, _16346_, _16342_);
  and (_16348_, _10209_, _10155_);
  nor (_16349_, _10204_, _10203_);
  or (_16350_, _16349_, _10205_);
  nor (_16351_, _16350_, _10209_);
  or (_16352_, _16351_, _16348_);
  or (_16353_, _16352_, _09861_);
  and (_16354_, _16353_, _06111_);
  and (_16355_, _16354_, _16347_);
  nand (_16356_, _07841_, _06945_);
  and (_16357_, _16356_, _06110_);
  and (_16358_, _16357_, _16295_);
  or (_16359_, _16358_, _16355_);
  and (_16360_, _16359_, _07127_);
  or (_16361_, _14346_, _10243_);
  and (_16362_, _16295_, _06297_);
  and (_16363_, _16362_, _16361_);
  or (_16364_, _16363_, _06402_);
  or (_16365_, _16364_, _16360_);
  and (_16366_, _10278_, _07841_);
  or (_16367_, _16366_, _16284_);
  or (_16368_, _16367_, _07125_);
  and (_16369_, _16368_, _07132_);
  and (_16370_, _16369_, _16365_);
  or (_16371_, _14344_, _10243_);
  and (_16372_, _16295_, _06306_);
  and (_16373_, _16372_, _16371_);
  or (_16374_, _16373_, _06411_);
  or (_16375_, _16374_, _16370_);
  and (_16376_, _16300_, _08176_);
  or (_16377_, _16284_, _07130_);
  or (_16378_, _16377_, _16376_);
  and (_16379_, _16378_, _08819_);
  and (_16380_, _16379_, _16375_);
  or (_16381_, _16356_, _08176_);
  and (_16382_, _16295_, _06303_);
  and (_16383_, _16382_, _16381_);
  or (_16384_, _16383_, _06396_);
  or (_16385_, _16384_, _16380_);
  and (_16386_, _16385_, _16287_);
  or (_16387_, _16386_, _06433_);
  or (_16388_, _16298_, _06829_);
  and (_16389_, _16388_, _05749_);
  and (_16390_, _16389_, _16387_);
  and (_16391_, _16290_, _05748_);
  or (_16392_, _16391_, _06440_);
  or (_16393_, _16392_, _16390_);
  or (_16394_, _16284_, _06444_);
  or (_16395_, _16394_, _16296_);
  and (_16396_, _16395_, _01317_);
  and (_16397_, _16396_, _16393_);
  or (_16398_, _16397_, _16283_);
  and (_43595_, _16398_, _43100_);
  nor (_16399_, _01317_, _09919_);
  nor (_16400_, _07841_, _09919_);
  and (_16401_, _07841_, _07708_);
  or (_16402_, _16401_, _16400_);
  or (_16403_, _16402_, _06132_);
  and (_16404_, _14538_, _08420_);
  and (_16405_, _16404_, _14569_);
  nor (_16406_, _08420_, _09919_);
  or (_16407_, _16406_, _06146_);
  or (_16408_, _16407_, _16405_);
  or (_16409_, _16402_, _07075_);
  and (_16410_, _14542_, _07841_);
  or (_16411_, _16410_, _16400_);
  or (_16412_, _16411_, _06161_);
  and (_16413_, _07841_, \oc8051_golden_model_1.ACC [2]);
  or (_16414_, _16413_, _16400_);
  and (_16415_, _16414_, _07056_);
  nor (_16416_, _07056_, _09919_);
  or (_16417_, _16416_, _06160_);
  or (_16418_, _16417_, _16415_);
  and (_16419_, _16418_, _06157_);
  and (_16420_, _16419_, _16412_);
  or (_16421_, _16406_, _16404_);
  and (_16422_, _16421_, _06156_);
  or (_16423_, _16422_, _06217_);
  or (_16424_, _16423_, _16420_);
  and (_16425_, _16424_, _16409_);
  or (_16426_, _16425_, _06220_);
  or (_16427_, _16414_, _06229_);
  and (_16428_, _16427_, _06153_);
  and (_16429_, _16428_, _16426_);
  and (_16430_, _14536_, _08420_);
  or (_16431_, _16430_, _16406_);
  and (_16432_, _16431_, _06152_);
  or (_16433_, _16432_, _06145_);
  or (_16434_, _16433_, _16429_);
  and (_16435_, _16434_, _16408_);
  or (_16436_, _16435_, _09295_);
  or (_16437_, _09801_, _09679_);
  and (_16438_, _16437_, _09802_);
  or (_16439_, _16438_, _09301_);
  and (_16440_, _16439_, _06140_);
  and (_16441_, _16440_, _16436_);
  and (_16442_, _14583_, _08420_);
  or (_16443_, _16442_, _16406_);
  and (_16444_, _16443_, _06139_);
  or (_16445_, _16444_, _09842_);
  or (_16446_, _16445_, _16441_);
  and (_16447_, _16446_, _16403_);
  or (_16448_, _16447_, _06116_);
  and (_16449_, _09211_, _07841_);
  or (_16450_, _16400_, _06117_);
  or (_16451_, _16450_, _16449_);
  and (_16452_, _16451_, _16448_);
  or (_16453_, _16452_, _05787_);
  and (_16454_, _14630_, _07841_);
  or (_16455_, _16400_, _06114_);
  or (_16456_, _16455_, _16454_);
  and (_16457_, _16456_, _09861_);
  and (_16458_, _16457_, _16453_);
  nor (_16459_, _10205_, _10156_);
  not (_16460_, _16459_);
  and (_16461_, _16460_, _10149_);
  nor (_16462_, _16460_, _10149_);
  nor (_16463_, _16462_, _16461_);
  or (_16464_, _16463_, _10209_);
  nand (_16465_, _10209_, _10146_);
  and (_16466_, _16465_, _09855_);
  and (_16467_, _16466_, _16464_);
  or (_16468_, _16467_, _11136_);
  or (_16469_, _16468_, _16458_);
  and (_16470_, _14646_, _07841_);
  or (_16471_, _16400_, _07127_);
  or (_16472_, _16471_, _16470_);
  and (_16473_, _07841_, _08768_);
  or (_16474_, _16473_, _16400_);
  or (_16475_, _16474_, _06111_);
  and (_16476_, _16475_, _07125_);
  and (_16477_, _16476_, _16472_);
  and (_16478_, _16477_, _16469_);
  and (_16479_, _10282_, _07841_);
  or (_16480_, _16479_, _16400_);
  and (_16481_, _16480_, _06402_);
  or (_16482_, _16481_, _16478_);
  and (_16483_, _16482_, _07132_);
  or (_16484_, _16400_, _08248_);
  and (_16485_, _16474_, _06306_);
  and (_16486_, _16485_, _16484_);
  or (_16487_, _16486_, _16483_);
  and (_16488_, _16487_, _07130_);
  and (_16489_, _16414_, _06411_);
  and (_16490_, _16489_, _16484_);
  or (_16491_, _16490_, _06303_);
  or (_16492_, _16491_, _16488_);
  and (_16493_, _14643_, _07841_);
  or (_16494_, _16400_, _08819_);
  or (_16495_, _16494_, _16493_);
  and (_16496_, _16495_, _08824_);
  and (_16497_, _16496_, _16492_);
  nor (_16498_, _10281_, _10243_);
  or (_16499_, _16498_, _16400_);
  and (_16500_, _16499_, _06396_);
  or (_16501_, _16500_, _06433_);
  or (_16502_, _16501_, _16497_);
  or (_16503_, _16411_, _06829_);
  and (_16504_, _16503_, _05749_);
  and (_16505_, _16504_, _16502_);
  and (_16506_, _16431_, _05748_);
  or (_16507_, _16506_, _06440_);
  or (_16508_, _16507_, _16505_);
  and (_16509_, _14710_, _07841_);
  or (_16510_, _16400_, _06444_);
  or (_16511_, _16510_, _16509_);
  and (_16512_, _16511_, _01317_);
  and (_16513_, _16512_, _16508_);
  or (_16514_, _16513_, _16399_);
  and (_43596_, _16514_, _43100_);
  nor (_16515_, _01317_, _09951_);
  nor (_16516_, _07841_, _09951_);
  and (_16517_, _14825_, _07841_);
  or (_16518_, _16517_, _16516_);
  and (_16519_, _16518_, _05787_);
  nor (_16520_, _08420_, _09951_);
  and (_16521_, _14735_, _08420_);
  or (_16522_, _16521_, _16520_);
  or (_16523_, _16520_, _14764_);
  and (_16524_, _16523_, _16522_);
  or (_16525_, _16524_, _06146_);
  and (_16526_, _14738_, _07841_);
  or (_16527_, _16526_, _16516_);
  or (_16528_, _16527_, _06161_);
  and (_16529_, _07841_, \oc8051_golden_model_1.ACC [3]);
  or (_16530_, _16529_, _16516_);
  and (_16531_, _16530_, _07056_);
  nor (_16532_, _07056_, _09951_);
  or (_16533_, _16532_, _06160_);
  or (_16534_, _16533_, _16531_);
  and (_16535_, _16534_, _06157_);
  and (_16536_, _16535_, _16528_);
  and (_16537_, _16522_, _06156_);
  or (_16538_, _16537_, _06217_);
  or (_16539_, _16538_, _16536_);
  and (_16540_, _07841_, _07544_);
  or (_16541_, _16540_, _16516_);
  or (_16542_, _16541_, _07075_);
  and (_16543_, _16542_, _16539_);
  or (_16544_, _16543_, _06220_);
  or (_16545_, _16530_, _06229_);
  and (_16546_, _16545_, _06153_);
  and (_16547_, _16546_, _16544_);
  and (_16548_, _14731_, _08420_);
  or (_16549_, _16548_, _16520_);
  and (_16550_, _16549_, _06152_);
  or (_16551_, _16550_, _06145_);
  or (_16552_, _16551_, _16547_);
  and (_16553_, _16552_, _16525_);
  or (_16554_, _16553_, _09295_);
  nor (_16555_, _09805_, _09621_);
  nor (_16556_, _16555_, _09807_);
  or (_16557_, _16556_, _09301_);
  and (_16558_, _16557_, _06140_);
  and (_16559_, _16558_, _16554_);
  and (_16560_, _14732_, _08420_);
  or (_16561_, _16560_, _16520_);
  and (_16562_, _16561_, _06139_);
  or (_16563_, _16562_, _09842_);
  or (_16564_, _16563_, _16559_);
  or (_16565_, _16541_, _06132_);
  and (_16566_, _16565_, _16564_);
  or (_16567_, _16566_, _06116_);
  and (_16568_, _09210_, _07841_);
  or (_16569_, _16516_, _06117_);
  or (_16570_, _16569_, _16568_);
  and (_16571_, _16570_, _06114_);
  and (_16572_, _16571_, _16567_);
  or (_16573_, _16572_, _16519_);
  and (_16574_, _16573_, _09861_);
  nor (_16575_, _16461_, _10148_);
  nor (_16576_, _16575_, _10140_);
  and (_16577_, _16575_, _10140_);
  or (_16578_, _16577_, _16576_);
  or (_16579_, _16578_, _10209_);
  not (_16580_, _10209_);
  or (_16581_, _16580_, _10137_);
  and (_16582_, _16581_, _09855_);
  and (_16583_, _16582_, _16579_);
  or (_16584_, _16583_, _11136_);
  or (_16585_, _16584_, _16574_);
  and (_16586_, _14727_, _07841_);
  or (_16587_, _16516_, _07127_);
  or (_16588_, _16587_, _16586_);
  and (_16589_, _07841_, _08712_);
  or (_16590_, _16589_, _16516_);
  or (_16591_, _16590_, _06111_);
  and (_16592_, _16591_, _07125_);
  and (_16593_, _16592_, _16588_);
  and (_16594_, _16593_, _16585_);
  and (_16595_, _12318_, _07841_);
  or (_16596_, _16595_, _16516_);
  and (_16597_, _16596_, _06402_);
  or (_16598_, _16597_, _16594_);
  and (_16599_, _16598_, _07132_);
  or (_16600_, _16516_, _08140_);
  and (_16601_, _16590_, _06306_);
  and (_16602_, _16601_, _16600_);
  or (_16603_, _16602_, _16599_);
  and (_16604_, _16603_, _07130_);
  and (_16605_, _16530_, _06411_);
  and (_16606_, _16605_, _16600_);
  or (_16607_, _16606_, _06303_);
  or (_16608_, _16607_, _16604_);
  and (_16609_, _14724_, _07841_);
  or (_16610_, _16516_, _08819_);
  or (_16611_, _16610_, _16609_);
  and (_16612_, _16611_, _08824_);
  and (_16613_, _16612_, _16608_);
  nor (_16614_, _10273_, _10243_);
  or (_16615_, _16614_, _16516_);
  and (_16616_, _16615_, _06396_);
  or (_16617_, _16616_, _06433_);
  or (_16618_, _16617_, _16613_);
  or (_16619_, _16527_, _06829_);
  and (_16620_, _16619_, _05749_);
  and (_16621_, _16620_, _16618_);
  and (_16622_, _16549_, _05748_);
  or (_16623_, _16622_, _06440_);
  or (_16624_, _16623_, _16621_);
  and (_16625_, _14897_, _07841_);
  or (_16626_, _16516_, _06444_);
  or (_16627_, _16626_, _16625_);
  and (_16628_, _16627_, _01317_);
  and (_16629_, _16628_, _16624_);
  or (_16630_, _16629_, _16515_);
  and (_43598_, _16630_, _43100_);
  nor (_16631_, _01317_, _09876_);
  nor (_16632_, _07841_, _09876_);
  and (_16633_, _15013_, _07841_);
  or (_16634_, _16633_, _16632_);
  and (_16635_, _16634_, _05787_);
  and (_16636_, _08336_, _07841_);
  or (_16637_, _16636_, _16632_);
  or (_16638_, _16637_, _06132_);
  nor (_16639_, _08420_, _09876_);
  and (_16640_, _14942_, _08420_);
  or (_16641_, _16640_, _16639_);
  and (_16642_, _16641_, _06152_);
  and (_16643_, _14928_, _07841_);
  or (_16644_, _16643_, _16632_);
  or (_16645_, _16644_, _06161_);
  and (_16646_, _07841_, \oc8051_golden_model_1.ACC [4]);
  or (_16647_, _16646_, _16632_);
  and (_16648_, _16647_, _07056_);
  nor (_16649_, _07056_, _09876_);
  or (_16650_, _16649_, _06160_);
  or (_16651_, _16650_, _16648_);
  and (_16652_, _16651_, _06157_);
  and (_16653_, _16652_, _16645_);
  and (_16654_, _14932_, _08420_);
  or (_16655_, _16654_, _16639_);
  and (_16656_, _16655_, _06156_);
  or (_16657_, _16656_, _06217_);
  or (_16658_, _16657_, _16653_);
  or (_16659_, _16637_, _07075_);
  and (_16660_, _16659_, _16658_);
  or (_16661_, _16660_, _06220_);
  or (_16662_, _16647_, _06229_);
  and (_16663_, _16662_, _06153_);
  and (_16664_, _16663_, _16661_);
  or (_16665_, _16664_, _16642_);
  and (_16666_, _16665_, _06146_);
  or (_16667_, _16639_, _14949_);
  and (_16668_, _16655_, _06145_);
  and (_16669_, _16668_, _16667_);
  or (_16670_, _16669_, _09295_);
  or (_16671_, _16670_, _16666_);
  or (_16672_, _09811_, _09808_);
  and (_16673_, _16672_, _09813_);
  or (_16674_, _16673_, _09301_);
  and (_16675_, _16674_, _06140_);
  and (_16676_, _16675_, _16671_);
  and (_16677_, _14966_, _08420_);
  or (_16678_, _16677_, _16639_);
  and (_16679_, _16678_, _06139_);
  or (_16680_, _16679_, _09842_);
  or (_16681_, _16680_, _16676_);
  and (_16682_, _16681_, _16638_);
  or (_16683_, _16682_, _06116_);
  and (_16684_, _09209_, _07841_);
  or (_16685_, _16632_, _06117_);
  or (_16686_, _16685_, _16684_);
  and (_16687_, _16686_, _06114_);
  and (_16688_, _16687_, _16683_);
  or (_16689_, _16688_, _16635_);
  and (_16690_, _16689_, _09861_);
  or (_16691_, _16580_, _10175_);
  nor (_16692_, _16575_, _10139_);
  or (_16693_, _16692_, _10138_);
  nand (_16694_, _16693_, _10178_);
  or (_16695_, _16693_, _10178_);
  and (_16696_, _16695_, _16694_);
  or (_16697_, _16696_, _10209_);
  and (_16698_, _16697_, _09855_);
  and (_16699_, _16698_, _16691_);
  or (_16700_, _16699_, _11136_);
  or (_16701_, _16700_, _16690_);
  and (_16702_, _15029_, _07841_);
  or (_16703_, _16632_, _07127_);
  or (_16704_, _16703_, _16702_);
  and (_16705_, _08715_, _07841_);
  or (_16706_, _16705_, _16632_);
  or (_16707_, _16706_, _06111_);
  and (_16708_, _16707_, _07125_);
  and (_16709_, _16708_, _16704_);
  and (_16710_, _16709_, _16701_);
  and (_16711_, _10289_, _07841_);
  or (_16712_, _16711_, _16632_);
  and (_16713_, _16712_, _06402_);
  or (_16714_, _16713_, _16710_);
  and (_16715_, _16714_, _07132_);
  or (_16716_, _16632_, _08339_);
  and (_16717_, _16706_, _06306_);
  and (_16718_, _16717_, _16716_);
  or (_16719_, _16718_, _16715_);
  and (_16720_, _16719_, _07130_);
  and (_16721_, _16647_, _06411_);
  and (_16722_, _16721_, _16716_);
  or (_16723_, _16722_, _06303_);
  or (_16724_, _16723_, _16720_);
  and (_16725_, _15026_, _07841_);
  or (_16726_, _16632_, _08819_);
  or (_16727_, _16726_, _16725_);
  and (_16728_, _16727_, _08824_);
  and (_16729_, _16728_, _16724_);
  nor (_16730_, _10288_, _10243_);
  or (_16731_, _16730_, _16632_);
  and (_16732_, _16731_, _06396_);
  or (_16733_, _16732_, _06433_);
  or (_16734_, _16733_, _16729_);
  or (_16735_, _16644_, _06829_);
  and (_16736_, _16735_, _05749_);
  and (_16737_, _16736_, _16734_);
  and (_16738_, _16641_, _05748_);
  or (_16739_, _16738_, _06440_);
  or (_16740_, _16739_, _16737_);
  and (_16741_, _15087_, _07841_);
  or (_16742_, _16632_, _06444_);
  or (_16743_, _16742_, _16741_);
  and (_16744_, _16743_, _01317_);
  and (_16745_, _16744_, _16740_);
  or (_16746_, _16745_, _16631_);
  and (_43599_, _16746_, _43100_);
  nor (_16747_, _01317_, _09877_);
  nor (_16748_, _07841_, _09877_);
  and (_16749_, _15203_, _07841_);
  or (_16750_, _16749_, _16748_);
  and (_16751_, _16750_, _05787_);
  and (_16752_, _08101_, _07841_);
  or (_16753_, _16752_, _16748_);
  or (_16754_, _16753_, _06132_);
  nor (_16755_, _08420_, _09877_);
  and (_16756_, _15104_, _08420_);
  or (_16757_, _16756_, _16755_);
  and (_16758_, _16757_, _06152_);
  and (_16759_, _15119_, _07841_);
  or (_16760_, _16759_, _16748_);
  or (_16761_, _16760_, _06161_);
  and (_16762_, _07841_, \oc8051_golden_model_1.ACC [5]);
  or (_16763_, _16762_, _16748_);
  and (_16764_, _16763_, _07056_);
  nor (_16765_, _07056_, _09877_);
  or (_16766_, _16765_, _06160_);
  or (_16767_, _16766_, _16764_);
  and (_16768_, _16767_, _06157_);
  and (_16769_, _16768_, _16761_);
  and (_16770_, _15123_, _08420_);
  or (_16771_, _16770_, _16755_);
  and (_16772_, _16771_, _06156_);
  or (_16773_, _16772_, _06217_);
  or (_16774_, _16773_, _16769_);
  or (_16775_, _16753_, _07075_);
  and (_16776_, _16775_, _16774_);
  or (_16777_, _16776_, _06220_);
  or (_16778_, _16763_, _06229_);
  and (_16779_, _16778_, _06153_);
  and (_16780_, _16779_, _16777_);
  or (_16781_, _16780_, _16758_);
  and (_16782_, _16781_, _06146_);
  or (_16783_, _16755_, _15138_);
  and (_16784_, _16771_, _06145_);
  and (_16785_, _16784_, _16783_);
  or (_16786_, _16785_, _09295_);
  or (_16787_, _16786_, _16782_);
  or (_16788_, _09492_, _09493_);
  and (_16789_, _16788_, _09814_);
  nor (_16790_, _16789_, _09816_);
  or (_16791_, _16790_, _09301_);
  and (_16792_, _16791_, _06140_);
  and (_16793_, _16792_, _16787_);
  and (_16794_, _15155_, _08420_);
  or (_16795_, _16794_, _16755_);
  and (_16796_, _16795_, _06139_);
  or (_16797_, _16796_, _09842_);
  or (_16798_, _16797_, _16793_);
  and (_16799_, _16798_, _16754_);
  or (_16800_, _16799_, _06116_);
  and (_16801_, _09208_, _07841_);
  or (_16802_, _16748_, _06117_);
  or (_16803_, _16802_, _16801_);
  and (_16804_, _16803_, _06114_);
  and (_16805_, _16804_, _16800_);
  or (_16806_, _16805_, _16751_);
  and (_16807_, _16806_, _09861_);
  not (_16808_, _10177_);
  and (_16809_, _16694_, _16808_);
  nor (_16810_, _16809_, _10189_);
  and (_16811_, _16809_, _10189_);
  or (_16812_, _16811_, _16810_);
  nor (_16813_, _10209_, _09861_);
  and (_16814_, _16813_, _16812_);
  and (_16815_, _10186_, _09855_);
  and (_16816_, _16815_, _10209_);
  or (_16817_, _16816_, _11136_);
  or (_16818_, _16817_, _16814_);
  or (_16819_, _16818_, _16807_);
  and (_16820_, _15219_, _07841_);
  or (_16821_, _16748_, _07127_);
  or (_16822_, _16821_, _16820_);
  and (_16823_, _08736_, _07841_);
  or (_16824_, _16823_, _16748_);
  or (_16825_, _16824_, _06111_);
  and (_16826_, _16825_, _07125_);
  and (_16827_, _16826_, _16822_);
  and (_16828_, _16827_, _16819_);
  and (_16829_, _12325_, _07841_);
  or (_16830_, _16829_, _16748_);
  and (_16831_, _16830_, _06402_);
  or (_16832_, _16831_, _16828_);
  and (_16833_, _16832_, _07132_);
  or (_16834_, _16748_, _08104_);
  and (_16835_, _16824_, _06306_);
  and (_16836_, _16835_, _16834_);
  or (_16837_, _16836_, _16833_);
  and (_16838_, _16837_, _07130_);
  and (_16839_, _16763_, _06411_);
  and (_16840_, _16839_, _16834_);
  or (_16841_, _16840_, _06303_);
  or (_16842_, _16841_, _16838_);
  and (_16843_, _15216_, _07841_);
  or (_16844_, _16748_, _08819_);
  or (_16845_, _16844_, _16843_);
  and (_16846_, _16845_, _08824_);
  and (_16847_, _16846_, _16842_);
  nor (_16848_, _10269_, _10243_);
  or (_16849_, _16848_, _16748_);
  and (_16850_, _16849_, _06396_);
  or (_16851_, _16850_, _06433_);
  or (_16852_, _16851_, _16847_);
  or (_16853_, _16760_, _06829_);
  and (_16854_, _16853_, _05749_);
  and (_16855_, _16854_, _16852_);
  and (_16856_, _16757_, _05748_);
  or (_16857_, _16856_, _06440_);
  or (_16858_, _16857_, _16855_);
  and (_16859_, _15275_, _07841_);
  or (_16860_, _16748_, _06444_);
  or (_16861_, _16860_, _16859_);
  and (_16862_, _16861_, _01317_);
  and (_16863_, _16862_, _16858_);
  or (_16864_, _16863_, _16747_);
  and (_43600_, _16864_, _43100_);
  nor (_16865_, _01317_, _10120_);
  nor (_16866_, _07841_, _10120_);
  and (_16867_, _15395_, _07841_);
  or (_16868_, _16867_, _16866_);
  and (_16869_, _16868_, _05787_);
  and (_16870_, _08012_, _07841_);
  or (_16871_, _16870_, _16866_);
  or (_16872_, _16871_, _06132_);
  nor (_16873_, _08420_, _10120_);
  and (_16874_, _15297_, _08420_);
  or (_16875_, _16874_, _16873_);
  and (_16876_, _16875_, _06152_);
  and (_16877_, _15300_, _07841_);
  or (_16878_, _16877_, _16866_);
  or (_16879_, _16878_, _06161_);
  and (_16880_, _07841_, \oc8051_golden_model_1.ACC [6]);
  or (_16881_, _16880_, _16866_);
  and (_16882_, _16881_, _07056_);
  nor (_16883_, _07056_, _10120_);
  or (_16884_, _16883_, _06160_);
  or (_16885_, _16884_, _16882_);
  and (_16886_, _16885_, _06157_);
  and (_16887_, _16886_, _16879_);
  and (_16888_, _15316_, _08420_);
  or (_16889_, _16888_, _16873_);
  and (_16890_, _16889_, _06156_);
  or (_16891_, _16890_, _06217_);
  or (_16892_, _16891_, _16887_);
  or (_16893_, _16871_, _07075_);
  and (_16894_, _16893_, _16892_);
  or (_16895_, _16894_, _06220_);
  or (_16896_, _16881_, _06229_);
  and (_16897_, _16896_, _06153_);
  and (_16898_, _16897_, _16895_);
  or (_16899_, _16898_, _16876_);
  and (_16900_, _16899_, _06146_);
  or (_16901_, _16873_, _15331_);
  and (_16902_, _16889_, _06145_);
  and (_16903_, _16902_, _16901_);
  or (_16904_, _16903_, _09295_);
  or (_16905_, _16904_, _16900_);
  nor (_16906_, _09834_, _09817_);
  nor (_16907_, _16906_, _09835_);
  or (_16908_, _16907_, _09301_);
  and (_16909_, _16908_, _06140_);
  and (_16910_, _16909_, _16905_);
  and (_16911_, _15348_, _08420_);
  or (_16912_, _16911_, _16873_);
  and (_16913_, _16912_, _06139_);
  or (_16914_, _16913_, _09842_);
  or (_16915_, _16914_, _16910_);
  and (_16916_, _16915_, _16872_);
  or (_16917_, _16916_, _06116_);
  and (_16918_, _09207_, _07841_);
  or (_16919_, _16866_, _06117_);
  or (_16920_, _16919_, _16918_);
  and (_16921_, _16920_, _06114_);
  and (_16922_, _16921_, _16917_);
  or (_16923_, _16922_, _16869_);
  and (_16924_, _16923_, _09861_);
  nor (_16925_, _16809_, _10187_);
  or (_16926_, _16925_, _10188_);
  and (_16927_, _16926_, _10169_);
  nor (_16928_, _16926_, _10169_);
  or (_16929_, _16928_, _16927_);
  or (_16930_, _16929_, _10209_);
  or (_16931_, _16580_, _10126_);
  and (_16932_, _16931_, _09855_);
  and (_16933_, _16932_, _16930_);
  or (_16934_, _16933_, _11136_);
  or (_16935_, _16934_, _16924_);
  and (_16936_, _15413_, _07841_);
  or (_16937_, _16866_, _07127_);
  or (_16938_, _16937_, _16936_);
  and (_16939_, _15402_, _07841_);
  or (_16940_, _16939_, _16866_);
  or (_16941_, _16940_, _06111_);
  and (_16942_, _16941_, _07125_);
  and (_16943_, _16942_, _16938_);
  and (_16944_, _16943_, _16935_);
  and (_16945_, _10295_, _07841_);
  or (_16946_, _16945_, _16866_);
  and (_16947_, _16946_, _06402_);
  or (_16948_, _16947_, _16944_);
  and (_16949_, _16948_, _07132_);
  or (_16950_, _16866_, _08015_);
  and (_16951_, _16940_, _06306_);
  and (_16952_, _16951_, _16950_);
  or (_16953_, _16952_, _16949_);
  and (_16954_, _16953_, _07130_);
  and (_16955_, _16881_, _06411_);
  and (_16956_, _16955_, _16950_);
  or (_16957_, _16956_, _06303_);
  or (_16958_, _16957_, _16954_);
  and (_16959_, _15410_, _07841_);
  or (_16960_, _16866_, _08819_);
  or (_16961_, _16960_, _16959_);
  and (_16962_, _16961_, _08824_);
  and (_16963_, _16962_, _16958_);
  nor (_16964_, _10294_, _10243_);
  or (_16965_, _16964_, _16866_);
  and (_16966_, _16965_, _06396_);
  or (_16967_, _16966_, _06433_);
  or (_16968_, _16967_, _16963_);
  or (_16969_, _16878_, _06829_);
  and (_16970_, _16969_, _05749_);
  and (_16971_, _16970_, _16968_);
  and (_16972_, _16875_, _05748_);
  or (_16973_, _16972_, _06440_);
  or (_16974_, _16973_, _16971_);
  and (_16975_, _15478_, _07841_);
  or (_16976_, _16866_, _06444_);
  or (_16977_, _16976_, _16975_);
  and (_16978_, _16977_, _01317_);
  and (_16979_, _16978_, _16974_);
  or (_16980_, _16979_, _16865_);
  and (_43601_, _16980_, _43100_);
  nor (_16981_, _01317_, _05855_);
  nand (_16982_, _10262_, _08430_);
  nand (_16983_, _12322_, _06169_);
  and (_16984_, _16983_, _10265_);
  nor (_16985_, _07049_, \oc8051_golden_model_1.ACC [0]);
  nor (_16986_, _10985_, _16985_);
  not (_16987_, _10962_);
  and (_16988_, _16987_, _16986_);
  and (_16989_, _14167_, _07809_);
  nor (_16990_, _07809_, _05855_);
  or (_16991_, _16990_, _08819_);
  or (_16992_, _16991_, _16989_);
  nor (_16993_, _09160_, \oc8051_golden_model_1.ACC [0]);
  nand (_16994_, _10841_, _16993_);
  and (_16995_, _14275_, _07809_);
  or (_16996_, _16990_, _07127_);
  or (_16997_, _16996_, _16995_);
  nand (_16998_, _06107_, _05801_);
  and (_16999_, _14260_, _07809_);
  or (_17000_, _16999_, _16990_);
  and (_17001_, _17000_, _05787_);
  and (_17002_, _07809_, _07049_);
  or (_17003_, _17002_, _16990_);
  or (_17004_, _17003_, _06132_);
  nor (_17005_, _10627_, _05855_);
  or (_17006_, _17005_, _10628_);
  or (_17007_, _17006_, _12380_);
  or (_17008_, _10458_, _07049_);
  nor (_17009_, _10473_, _07064_);
  or (_17010_, _17009_, _09160_);
  not (_17011_, _10471_);
  and (_17012_, _17011_, _07049_);
  or (_17013_, _06653_, \oc8051_golden_model_1.ACC [0]);
  nand (_17014_, _06653_, \oc8051_golden_model_1.ACC [0]);
  and (_17015_, _17014_, _17013_);
  and (_17016_, _17015_, _10471_);
  or (_17017_, _17016_, _10473_);
  or (_17018_, _17017_, _17012_);
  and (_17019_, _17018_, _05772_);
  or (_17020_, _17019_, _07064_);
  and (_17021_, _17020_, _06161_);
  and (_17022_, _17021_, _17010_);
  not (_17023_, _07809_);
  nor (_17024_, _08211_, _17023_);
  nor (_17025_, _17024_, _16990_);
  nor (_17026_, _17025_, _06161_);
  or (_17027_, _17026_, _06156_);
  or (_17028_, _17027_, _17022_);
  and (_17029_, _14169_, _08409_);
  nor (_17030_, _08409_, _05855_);
  or (_17031_, _17030_, _06157_);
  or (_17032_, _17031_, _17029_);
  and (_17033_, _17032_, _07075_);
  and (_17034_, _17033_, _17028_);
  and (_17035_, _17003_, _06217_);
  or (_17036_, _17035_, _10516_);
  or (_17037_, _17036_, _17034_);
  and (_17038_, _17037_, _17008_);
  or (_17039_, _17038_, _07081_);
  or (_17040_, _09160_, _07082_);
  and (_17041_, _17040_, _06229_);
  and (_17042_, _17041_, _17039_);
  and (_17043_, _08211_, _06220_);
  or (_17044_, _17043_, _10525_);
  or (_17045_, _17044_, _17042_);
  nand (_17046_, _10525_, _09902_);
  and (_17047_, _17046_, _17045_);
  or (_17048_, _17047_, _06152_);
  or (_17049_, _16990_, _06153_);
  and (_17050_, _17049_, _06146_);
  nand (_17051_, _17050_, _17048_);
  or (_17052_, _17025_, _06146_);
  and (_17053_, _17052_, _09301_);
  and (_17054_, _17053_, _17051_);
  nand (_17055_, _16232_, _09295_);
  nand (_17056_, _17055_, _10554_);
  nor (_17057_, _17056_, _17054_);
  nor (_17058_, _10354_, _05855_);
  nor (_17059_, _17058_, _10562_);
  or (_17060_, _17059_, _10554_);
  nand (_17061_, _17060_, _12380_);
  or (_17062_, _17061_, _17057_);
  and (_17063_, _17062_, _17007_);
  or (_17064_, _17063_, _06260_);
  nor (_17065_, _10434_, _05855_);
  or (_17066_, _17065_, _10435_);
  or (_17067_, _17066_, _06265_);
  and (_17068_, _17067_, _10388_);
  and (_17069_, _17068_, _17064_);
  nor (_17070_, _10701_, _05855_);
  or (_17071_, _17070_, _10702_);
  and (_17072_, _17071_, _10387_);
  or (_17073_, _17072_, _05870_);
  or (_17074_, _17073_, _17069_);
  nand (_17075_, _06107_, _05870_);
  and (_17076_, _17075_, _06140_);
  and (_17077_, _17076_, _17074_);
  and (_17078_, _14171_, _08409_);
  or (_17079_, _17078_, _17030_);
  and (_17080_, _17079_, _06139_);
  or (_17081_, _17080_, _09842_);
  or (_17082_, _17081_, _17077_);
  and (_17083_, _17082_, _17004_);
  or (_17084_, _17083_, _06116_);
  and (_17085_, _09160_, _07809_);
  or (_17086_, _16990_, _06117_);
  or (_17087_, _17086_, _17085_);
  and (_17088_, _17087_, _06114_);
  and (_17089_, _17088_, _17084_);
  or (_17090_, _17089_, _17001_);
  and (_17091_, _17090_, _09861_);
  or (_17092_, _16813_, _05801_);
  or (_17093_, _17092_, _17091_);
  and (_17094_, _17093_, _16998_);
  or (_17095_, _17094_, _06110_);
  and (_17096_, _07809_, _08708_);
  or (_17097_, _17096_, _16990_);
  or (_17098_, _17097_, _06111_);
  and (_17099_, _17098_, _10752_);
  and (_17100_, _17099_, _17095_);
  nor (_17101_, _10752_, _06107_);
  or (_17102_, _17101_, _06558_);
  or (_17103_, _17102_, _17100_);
  or (_17104_, _16986_, _10762_);
  and (_17105_, _06288_, _06399_);
  nor (_17106_, _17105_, _10768_);
  and (_17107_, _17106_, _17104_);
  and (_17108_, _17107_, _17103_);
  not (_17109_, _17106_);
  and (_17110_, _17109_, _16986_);
  or (_17111_, _17110_, _06771_);
  or (_17112_, _17111_, _17108_);
  not (_17113_, _06771_);
  or (_17114_, _16986_, _17113_);
  and (_17115_, _17114_, _17112_);
  or (_17116_, _17115_, _10775_);
  nor (_17117_, _11027_, _16993_);
  or (_17118_, _10776_, _17117_);
  and (_17119_, _17118_, _17116_);
  or (_17120_, _17119_, _06400_);
  nand (_17121_, _12322_, _06400_);
  and (_17122_, _17121_, _10788_);
  and (_17123_, _17122_, _17120_);
  and (_17124_, _10787_, _12339_);
  or (_17125_, _17124_, _06297_);
  or (_17126_, _17125_, _17123_);
  and (_17127_, _17126_, _16997_);
  or (_17128_, _17127_, _06402_);
  or (_17129_, _16990_, _07125_);
  and (_17130_, _17129_, _10808_);
  and (_17131_, _17130_, _17128_);
  and (_17132_, _10812_, _10985_);
  or (_17133_, _17132_, _10811_);
  or (_17134_, _17133_, _17131_);
  or (_17135_, _10816_, _11027_);
  and (_17136_, _17135_, _06410_);
  and (_17137_, _17136_, _17134_);
  or (_17138_, _10820_, _10276_);
  and (_17139_, _17138_, _10822_);
  or (_17140_, _17139_, _17137_);
  or (_17141_, _10826_, _11067_);
  and (_17142_, _17141_, _07132_);
  and (_17143_, _17142_, _17140_);
  nand (_17144_, _17097_, _06306_);
  nor (_17145_, _17144_, _17024_);
  or (_17146_, _17145_, _06524_);
  or (_17147_, _17146_, _17143_);
  and (_17148_, _06957_, _05840_);
  or (_17149_, _17148_, _06555_);
  not (_17150_, _17149_);
  nand (_17151_, _16985_, _06524_);
  and (_17152_, _17151_, _17150_);
  and (_17153_, _17152_, _17147_);
  and (_17154_, _06684_, _05840_);
  and (_17155_, _06288_, _05840_);
  or (_17156_, _17155_, _17154_);
  nor (_17157_, _17150_, _16985_);
  or (_17158_, _17157_, _17156_);
  or (_17159_, _17158_, _17153_);
  and (_17160_, _06273_, _05840_);
  not (_17161_, _17160_);
  nand (_17162_, _17156_, _16985_);
  and (_17163_, _17162_, _17161_);
  and (_17164_, _17163_, _17159_);
  nor (_17165_, _16985_, _17161_);
  or (_17166_, _17165_, _10841_);
  or (_17167_, _17166_, _17164_);
  and (_17168_, _17167_, _16994_);
  or (_17169_, _17168_, _06394_);
  nand (_17170_, _12321_, _06394_);
  and (_17171_, _17170_, _10851_);
  and (_17172_, _17171_, _17169_);
  nor (_17173_, _10851_, _12338_);
  or (_17174_, _17173_, _06303_);
  or (_17175_, _17174_, _17172_);
  and (_17176_, _17175_, _16992_);
  or (_17177_, _17176_, _10858_);
  nand (_17178_, _17059_, _10858_);
  and (_17179_, _17178_, _10867_);
  and (_17180_, _17179_, _17177_);
  and (_17181_, _10865_, _17006_);
  or (_17182_, _17181_, _06406_);
  or (_17183_, _17182_, _17180_);
  or (_17184_, _17066_, _06407_);
  and (_17185_, _17184_, _10927_);
  and (_17186_, _17185_, _17183_);
  and (_17187_, _10895_, _17071_);
  or (_17188_, _17187_, _10925_);
  or (_17189_, _17188_, _17186_);
  nand (_17190_, _10925_, _10693_);
  and (_17191_, _17190_, _10962_);
  and (_17192_, _17191_, _17189_);
  or (_17193_, _17192_, _16988_);
  and (_17194_, _17193_, _10957_);
  and (_17195_, _06284_, _05825_);
  and (_17196_, _16986_, _10956_);
  or (_17197_, _17196_, _17195_);
  or (_17198_, _17197_, _17194_);
  and (_17199_, _06281_, _05825_);
  not (_17200_, _17199_);
  not (_17201_, _17195_);
  or (_17202_, _17201_, _17117_);
  and (_17203_, _17202_, _17200_);
  and (_17204_, _17203_, _17198_);
  and (_17205_, _17117_, _17199_);
  or (_17206_, _17205_, _06169_);
  or (_17207_, _17206_, _17204_);
  and (_17208_, _17207_, _16984_);
  and (_17209_, _12339_, _10264_);
  or (_17210_, _17209_, _10262_);
  or (_17211_, _17210_, _17208_);
  and (_17212_, _17211_, _16982_);
  or (_17213_, _17212_, _06433_);
  nand (_17214_, _17025_, _06433_);
  and (_17215_, _17214_, _11090_);
  and (_17216_, _17215_, _17213_);
  nor (_17217_, _11094_, _05855_);
  nor (_17218_, _17217_, _12719_);
  or (_17219_, _17218_, _17216_);
  nand (_17220_, _11094_, _05887_);
  and (_17221_, _17220_, _05749_);
  and (_17222_, _17221_, _17219_);
  and (_17223_, _16990_, _05748_);
  or (_17224_, _17223_, _06440_);
  or (_17225_, _17224_, _17222_);
  nand (_17226_, _17025_, _06440_);
  and (_17227_, _17226_, _11113_);
  and (_17228_, _17227_, _17225_);
  nor (_17229_, _11119_, _05855_);
  nor (_17230_, _17229_, _12744_);
  or (_17231_, _17230_, _17228_);
  nand (_17232_, _11119_, _05887_);
  and (_17233_, _17232_, _01317_);
  and (_17234_, _17233_, _17231_);
  or (_17235_, _17234_, _16981_);
  and (_43603_, _17235_, _43100_);
  nor (_17236_, _01317_, _05887_);
  or (_17237_, _10906_, _10905_);
  nor (_17238_, _10907_, _06407_);
  and (_17239_, _17238_, _17237_);
  and (_17240_, _06284_, _06300_);
  not (_17241_, _17240_);
  not (_17242_, _10841_);
  or (_17243_, _17242_, _11024_);
  nor (_17244_, _10835_, _17154_);
  nor (_17245_, _10983_, _17160_);
  or (_17246_, _17245_, _17244_);
  or (_17247_, _10816_, _11023_);
  not (_17248_, _10984_);
  and (_17249_, _17106_, _10762_);
  nor (_17250_, _17249_, _17248_);
  nor (_17251_, _07809_, _05887_);
  and (_17252_, _07809_, _07306_);
  or (_17253_, _17252_, _17251_);
  or (_17254_, _17253_, _06132_);
  or (_17255_, _10458_, _07306_);
  or (_17256_, _17009_, _09115_);
  and (_17257_, _17011_, _07306_);
  or (_17258_, _06653_, \oc8051_golden_model_1.ACC [1]);
  nand (_17259_, _06653_, \oc8051_golden_model_1.ACC [1]);
  and (_17260_, _17259_, _17258_);
  and (_17261_, _17260_, _10471_);
  or (_17262_, _17261_, _10473_);
  or (_17263_, _17262_, _17257_);
  and (_17264_, _17263_, _05772_);
  or (_17265_, _17264_, _07064_);
  and (_17266_, _17265_, _17256_);
  or (_17267_, _17266_, _06160_);
  or (_17268_, _07809_, \oc8051_golden_model_1.ACC [1]);
  and (_17269_, _14363_, _07809_);
  not (_17270_, _17269_);
  and (_17271_, _17270_, _17268_);
  or (_17272_, _17271_, _06161_);
  and (_17273_, _17272_, _17267_);
  or (_17274_, _17273_, _10490_);
  nor (_17275_, _10494_, \oc8051_golden_model_1.PSW [6]);
  nor (_17276_, _17275_, \oc8051_golden_model_1.ACC [1]);
  and (_17277_, _17275_, \oc8051_golden_model_1.ACC [1]);
  nor (_17278_, _17277_, _17276_);
  nand (_17279_, _17278_, _10490_);
  and (_17280_, _17279_, _06221_);
  and (_17281_, _17280_, _17274_);
  nor (_17282_, _08409_, _05887_);
  and (_17283_, _14367_, _08409_);
  or (_17284_, _17283_, _17282_);
  and (_17285_, _17284_, _06156_);
  and (_17286_, _17253_, _06217_);
  or (_17287_, _17286_, _10516_);
  or (_17288_, _17287_, _17285_);
  or (_17289_, _17288_, _17281_);
  and (_17290_, _17289_, _17255_);
  or (_17291_, _17290_, _07081_);
  or (_17292_, _09115_, _07082_);
  and (_17293_, _17292_, _06229_);
  and (_17294_, _17293_, _17291_);
  nor (_17295_, _08175_, _06229_);
  or (_17296_, _17295_, _10525_);
  or (_17297_, _17296_, _17294_);
  nand (_17298_, _10525_, _09930_);
  and (_17299_, _17298_, _17297_);
  or (_17300_, _17299_, _06152_);
  and (_17301_, _14349_, _08409_);
  or (_17302_, _17301_, _17282_);
  or (_17303_, _17302_, _06153_);
  and (_17304_, _17303_, _06146_);
  and (_17305_, _17304_, _17300_);
  or (_17306_, _17282_, _14382_);
  and (_17307_, _17284_, _06145_);
  and (_17308_, _17307_, _17306_);
  or (_17309_, _17308_, _09295_);
  or (_17310_, _17309_, _17305_);
  nor (_17311_, _09771_, _09770_);
  or (_17312_, _17311_, _09772_);
  nand (_17313_, _17312_, _09295_);
  and (_17314_, _17313_, _10554_);
  and (_17315_, _17314_, _17310_);
  nor (_17316_, _10345_, _05855_);
  or (_17317_, _17316_, _10353_);
  or (_17318_, _17317_, _17248_);
  nand (_17319_, _17317_, _17248_);
  and (_17320_, _17319_, _17318_);
  and (_17321_, _17320_, _10557_);
  or (_17322_, _17321_, _17315_);
  and (_17323_, _17322_, _12380_);
  nor (_17324_, _10621_, _05855_);
  or (_17325_, _17324_, _10626_);
  nor (_17326_, _17325_, _11026_);
  and (_17327_, _17325_, _11026_);
  or (_17328_, _17327_, _17326_);
  and (_17329_, _17328_, _12379_);
  or (_17330_, _17329_, _17323_);
  and (_17331_, _17330_, _06265_);
  nor (_17332_, _10389_, _05855_);
  or (_17333_, _17332_, _10433_);
  nor (_17334_, _17333_, _10278_);
  and (_17335_, _17333_, _10278_);
  or (_17336_, _17335_, _10387_);
  or (_17337_, _17336_, _17334_);
  and (_17338_, _17337_, _12386_);
  or (_17339_, _17338_, _17331_);
  nor (_17340_, _06107_, \oc8051_golden_model_1.ACC [0]);
  nor (_17341_, _17340_, _11066_);
  and (_17342_, _17340_, _11066_);
  nor (_17343_, _17342_, _17341_);
  or (_17344_, _12339_, _10693_);
  and (_17345_, _17344_, _17343_);
  and (_17346_, _12340_, \oc8051_golden_model_1.PSW [7]);
  or (_17347_, _17346_, _17345_);
  or (_17348_, _17347_, _10388_);
  and (_17349_, _17348_, _17339_);
  or (_17350_, _17349_, _05870_);
  nand (_17351_, _06912_, _05870_);
  and (_17352_, _17351_, _06140_);
  and (_17353_, _17352_, _17350_);
  and (_17354_, _14351_, _08409_);
  or (_17355_, _17354_, _17282_);
  and (_17356_, _17355_, _06139_);
  or (_17357_, _17356_, _09842_);
  or (_17358_, _17357_, _17353_);
  and (_17359_, _17358_, _17254_);
  or (_17360_, _17359_, _06116_);
  and (_17361_, _09115_, _07809_);
  or (_17362_, _17251_, _06117_);
  or (_17363_, _17362_, _17361_);
  and (_17364_, _17363_, _06114_);
  and (_17365_, _17364_, _17360_);
  or (_17366_, _14442_, _17023_);
  and (_17367_, _17268_, _05787_);
  and (_17368_, _17367_, _17366_);
  or (_17369_, _17368_, _09855_);
  or (_17370_, _17369_, _17365_);
  or (_17371_, _10115_, _09861_);
  and (_17372_, _17371_, _17370_);
  or (_17373_, _17372_, _05801_);
  nand (_17374_, _06912_, _05801_);
  and (_17375_, _17374_, _06111_);
  and (_17377_, _17375_, _17373_);
  nand (_17378_, _07809_, _06945_);
  and (_17379_, _17378_, _06110_);
  and (_17380_, _17379_, _17268_);
  or (_17381_, _17380_, _10751_);
  or (_17382_, _17381_, _17377_);
  nand (_17383_, _10751_, _06912_);
  and (_17384_, _17383_, _17249_);
  and (_17385_, _17384_, _17382_);
  or (_17386_, _17385_, _17250_);
  and (_17388_, _17386_, _17113_);
  and (_17389_, _10984_, _06771_);
  or (_17390_, _17389_, _10775_);
  or (_17391_, _17390_, _17388_);
  or (_17392_, _10776_, _11026_);
  and (_17393_, _17392_, _17391_);
  or (_17394_, _17393_, _06400_);
  or (_17395_, _10278_, _06401_);
  and (_17396_, _17395_, _10788_);
  and (_17397_, _17396_, _17394_);
  and (_17399_, _10787_, _11066_);
  or (_17400_, _17399_, _17397_);
  and (_17401_, _17400_, _07127_);
  or (_17402_, _14346_, _17023_);
  and (_17403_, _17268_, _06297_);
  and (_17404_, _17403_, _17402_);
  or (_17405_, _17404_, _06402_);
  or (_17406_, _17405_, _17401_);
  and (_17407_, _06122_, _06408_);
  not (_17408_, _17407_);
  or (_17410_, _17251_, _07125_);
  and (_17411_, _17410_, _17408_);
  and (_17412_, _17411_, _17406_);
  and (_17413_, _17407_, _10982_);
  or (_17414_, _17413_, _06965_);
  or (_17415_, _17414_, _17412_);
  not (_17416_, _10807_);
  not (_17417_, _06965_);
  or (_17418_, _10982_, _17417_);
  and (_17419_, _17418_, _17416_);
  and (_17421_, _17419_, _17415_);
  and (_17422_, _10807_, _10982_);
  or (_17423_, _17422_, _10811_);
  or (_17424_, _17423_, _17421_);
  and (_17425_, _17424_, _17247_);
  or (_17426_, _17425_, _06409_);
  or (_17427_, _10275_, _06410_);
  and (_17428_, _17427_, _10826_);
  and (_17429_, _17428_, _17426_);
  and (_17430_, _10820_, _11064_);
  or (_17432_, _17430_, _17429_);
  and (_17433_, _17432_, _07132_);
  or (_17434_, _14344_, _17023_);
  and (_17435_, _17268_, _06306_);
  and (_17436_, _17435_, _17434_);
  or (_17437_, _17436_, _06524_);
  or (_17438_, _17437_, _17433_);
  nand (_17439_, _10983_, _06524_);
  and (_17440_, _17439_, _17150_);
  and (_17441_, _17440_, _17438_);
  nor (_17442_, _17150_, _10983_);
  or (_17443_, _17442_, _17156_);
  or (_17444_, _17443_, _17441_);
  and (_17445_, _17444_, _17246_);
  nor (_17446_, _10983_, _17161_);
  or (_17447_, _17446_, _10841_);
  or (_17448_, _17447_, _17445_);
  and (_17449_, _17448_, _17243_);
  or (_17450_, _17449_, _06394_);
  nand (_17451_, _10277_, _06394_);
  and (_17452_, _17451_, _10851_);
  and (_17453_, _17452_, _17450_);
  nor (_17454_, _10851_, _11065_);
  or (_17455_, _17454_, _17453_);
  and (_17456_, _17455_, _08819_);
  or (_17457_, _17378_, _08176_);
  and (_17458_, _17268_, _06303_);
  and (_17459_, _17458_, _17457_);
  or (_17460_, _17459_, _10858_);
  or (_17461_, _17460_, _17456_);
  nor (_17462_, _10355_, _10352_);
  nor (_17463_, _17462_, _10356_);
  or (_17464_, _17463_, _10380_);
  and (_17465_, _17464_, _17461_);
  and (_17466_, _17465_, _17241_);
  nor (_17467_, _10876_, _10875_);
  nor (_17468_, _17467_, _10877_);
  and (_17469_, _17468_, _17240_);
  or (_17470_, _17469_, _17466_);
  or (_17471_, _17470_, _06792_);
  or (_17472_, _17468_, _06793_);
  and (_17473_, _17472_, _06407_);
  and (_17474_, _17473_, _17471_);
  or (_17475_, _17474_, _17239_);
  and (_17476_, _17475_, _10927_);
  nor (_17477_, _10936_, _10935_);
  nor (_17478_, _17477_, _10937_);
  and (_17479_, _17478_, _10895_);
  or (_17480_, _17479_, _10925_);
  or (_17481_, _17480_, _17476_);
  nand (_17482_, _10925_, _05855_);
  and (_17483_, _17482_, _10963_);
  and (_17484_, _17483_, _17481_);
  or (_17485_, _10985_, _10984_);
  nor (_17486_, _10986_, _10963_);
  and (_17487_, _17486_, _17485_);
  or (_17488_, _17487_, _11003_);
  or (_17489_, _17488_, _17484_);
  nor (_17490_, _11027_, _11026_);
  nor (_17491_, _17490_, _11028_);
  or (_17492_, _17491_, _11041_);
  and (_17493_, _17492_, _06171_);
  and (_17494_, _17493_, _17489_);
  nor (_17495_, _10278_, _10276_);
  nor (_17496_, _17495_, _10279_);
  or (_17497_, _17496_, _10264_);
  and (_17498_, _17497_, _12691_);
  or (_17499_, _17498_, _17494_);
  nor (_17500_, _11067_, _11066_);
  nor (_17501_, _17500_, _11068_);
  or (_17502_, _17501_, _10265_);
  and (_17503_, _17502_, _12693_);
  and (_17504_, _17503_, _17499_);
  and (_17505_, _10262_, \oc8051_golden_model_1.ACC [0]);
  or (_17506_, _17505_, _06433_);
  or (_17507_, _17506_, _17504_);
  or (_17508_, _17271_, _06829_);
  and (_17509_, _17508_, _11090_);
  and (_17510_, _17509_, _17507_);
  nor (_17511_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  nor (_17512_, _11120_, _17511_);
  nor (_17513_, _17512_, _11090_);
  or (_17514_, _17513_, _11094_);
  or (_17515_, _17514_, _17510_);
  nand (_17516_, _11094_, _09981_);
  and (_17517_, _17516_, _05749_);
  and (_17518_, _17517_, _17515_);
  and (_17519_, _17302_, _05748_);
  or (_17520_, _17519_, _06440_);
  or (_17521_, _17520_, _17518_);
  or (_17522_, _17269_, _17251_);
  or (_17523_, _17522_, _06444_);
  and (_17524_, _17523_, _11113_);
  and (_17525_, _17524_, _17521_);
  and (_17526_, _17512_, _11112_);
  or (_17527_, _17526_, _11119_);
  or (_17528_, _17527_, _17525_);
  nand (_17529_, _11119_, _09981_);
  and (_17530_, _17529_, _01317_);
  and (_17531_, _17530_, _17528_);
  or (_17532_, _17531_, _17236_);
  and (_43604_, _17532_, _43100_);
  nor (_17533_, _01317_, _09981_);
  nand (_17534_, _10262_, _05887_);
  and (_17535_, _10283_, _10280_);
  nor (_17536_, _17535_, _10284_);
  or (_17537_, _17536_, _06171_);
  and (_17538_, _17537_, _10265_);
  nand (_17539_, _10908_, _10427_);
  nor (_17540_, _10909_, _06407_);
  and (_17541_, _17540_, _17539_);
  nand (_17542_, _10357_, _10344_);
  nor (_17543_, _10380_, _10358_);
  and (_17544_, _17543_, _17542_);
  nand (_17545_, _10848_, _11062_);
  and (_17546_, _06122_, _05840_);
  nand (_17547_, _17546_, _10979_);
  and (_17548_, _14646_, _07809_);
  nor (_17549_, _07809_, _09981_);
  or (_17550_, _17549_, _07127_);
  or (_17551_, _17550_, _17548_);
  or (_17552_, _10776_, _11021_);
  nor (_17553_, _10752_, _06625_);
  and (_17554_, _07809_, _07708_);
  or (_17555_, _17554_, _17549_);
  or (_17556_, _17555_, _06132_);
  and (_17557_, _08175_, \oc8051_golden_model_1.ACC [1]);
  and (_17558_, _08211_, _05855_);
  nor (_17559_, _17558_, _13920_);
  nor (_17560_, _17559_, _17557_);
  nor (_17561_, _17560_, _10282_);
  and (_17562_, _17560_, _10282_);
  nor (_17563_, _17562_, _17561_);
  and (_17564_, _12323_, \oc8051_golden_model_1.PSW [7]);
  or (_17565_, _17564_, _17563_);
  nand (_17566_, _17564_, _17563_);
  and (_17567_, _17566_, _17565_);
  or (_17568_, _17567_, _06265_);
  and (_17569_, _17568_, _10388_);
  or (_17570_, _10458_, _07708_);
  nor (_17571_, _08409_, _09981_);
  and (_17572_, _14538_, _08409_);
  or (_17573_, _17572_, _17571_);
  or (_17574_, _17573_, _06157_);
  and (_17575_, _17574_, _07075_);
  and (_17576_, _14542_, _07809_);
  or (_17577_, _17576_, _17549_);
  and (_17578_, _17577_, _06160_);
  or (_17579_, _17009_, _09211_);
  and (_17580_, _17011_, _07708_);
  or (_17581_, _06653_, \oc8051_golden_model_1.ACC [2]);
  nand (_17582_, _06653_, \oc8051_golden_model_1.ACC [2]);
  and (_17583_, _17582_, _17581_);
  and (_17584_, _17583_, _10471_);
  or (_17585_, _17584_, _10473_);
  or (_17586_, _17585_, _17580_);
  and (_17587_, _17586_, _05772_);
  or (_17588_, _17587_, _07064_);
  and (_17589_, _17588_, _06161_);
  and (_17590_, _17589_, _17579_);
  or (_17591_, _17590_, _17578_);
  and (_17592_, _17591_, _10491_);
  or (_17593_, _17276_, \oc8051_golden_model_1.ACC [2]);
  nand (_17594_, _17276_, \oc8051_golden_model_1.ACC [2]);
  and (_17595_, _17594_, _17593_);
  and (_17596_, _17595_, _10490_);
  or (_17597_, _17596_, _06156_);
  or (_17598_, _17597_, _17592_);
  and (_17599_, _17598_, _17575_);
  and (_17600_, _17555_, _06217_);
  or (_17601_, _17600_, _10516_);
  or (_17602_, _17601_, _17599_);
  and (_17603_, _17602_, _17570_);
  or (_17604_, _17603_, _07081_);
  or (_17605_, _09211_, _07082_);
  and (_17606_, _17605_, _06229_);
  and (_17607_, _17606_, _17604_);
  nor (_17608_, _08247_, _06229_);
  or (_17609_, _17608_, _10525_);
  or (_17610_, _17609_, _17607_);
  nand (_17611_, _10525_, _09883_);
  and (_17612_, _17611_, _17610_);
  or (_17613_, _17612_, _06152_);
  and (_17614_, _14536_, _08409_);
  or (_17615_, _17614_, _17571_);
  or (_17616_, _17615_, _06153_);
  and (_17617_, _17616_, _06146_);
  and (_17618_, _17617_, _17613_);
  or (_17619_, _17571_, _14569_);
  and (_17620_, _17573_, _06145_);
  and (_17621_, _17620_, _17619_);
  or (_17622_, _17621_, _09295_);
  or (_17623_, _17622_, _17618_);
  nor (_17624_, _09774_, _09772_);
  or (_17625_, _17624_, _09775_);
  nand (_17626_, _17625_, _09295_);
  and (_17627_, _17626_, _10554_);
  and (_17628_, _17627_, _17623_);
  and (_17629_, _07252_, \oc8051_golden_model_1.ACC [1]);
  and (_17630_, _07049_, _05855_);
  nor (_17631_, _17630_, _10984_);
  nor (_17632_, _17631_, _17629_);
  nor (_17633_, _10980_, _17632_);
  and (_17634_, _10980_, _17632_);
  nor (_17635_, _17634_, _17633_);
  nor (_17636_, _16986_, _10984_);
  and (_17637_, _17636_, \oc8051_golden_model_1.PSW [7]);
  nand (_17638_, _17637_, _17635_);
  or (_17639_, _17637_, _17635_);
  and (_17640_, _17639_, _10557_);
  and (_17641_, _17640_, _17638_);
  or (_17642_, _17641_, _10580_);
  or (_17643_, _17642_, _17628_);
  or (_17644_, _09115_, _05887_);
  and (_17645_, _09160_, _05855_);
  or (_17646_, _17645_, _11026_);
  and (_17647_, _17646_, _17644_);
  nor (_17648_, _11021_, _17647_);
  and (_17649_, _11021_, _17647_);
  nor (_17650_, _17649_, _17648_);
  nor (_17651_, _17117_, _11026_);
  not (_17652_, _17651_);
  or (_17653_, _17652_, _17650_);
  and (_17654_, _17653_, \oc8051_golden_model_1.PSW [7]);
  nor (_17655_, _17650_, \oc8051_golden_model_1.PSW [7]);
  nor (_17656_, _17655_, _17654_);
  and (_17657_, _17652_, _17650_);
  or (_17658_, _17657_, _17656_);
  and (_17659_, _17658_, _06276_);
  or (_17660_, _17659_, _12380_);
  and (_17661_, _17660_, _17643_);
  and (_17662_, _17658_, _06709_);
  or (_17663_, _17662_, _06260_);
  or (_17664_, _17663_, _17661_);
  and (_17665_, _17664_, _17569_);
  nor (_17666_, _17341_, _13944_);
  nor (_17667_, _11063_, _17666_);
  and (_17668_, _11063_, _17666_);
  nor (_17669_, _17668_, _17667_);
  nand (_17670_, _17346_, _17669_);
  or (_17671_, _17346_, _17669_);
  and (_17672_, _17671_, _17670_);
  and (_17673_, _17672_, _10387_);
  or (_17674_, _17673_, _05870_);
  or (_17675_, _17674_, _17665_);
  nand (_17676_, _06625_, _05870_);
  and (_17677_, _17676_, _06140_);
  and (_17678_, _17677_, _17675_);
  and (_17679_, _14583_, _08409_);
  or (_17680_, _17679_, _17571_);
  and (_17681_, _17680_, _06139_);
  or (_17682_, _17681_, _09842_);
  or (_17683_, _17682_, _17678_);
  and (_17684_, _17683_, _17556_);
  or (_17685_, _17684_, _06116_);
  and (_17686_, _09211_, _07809_);
  or (_17687_, _17549_, _06117_);
  or (_17688_, _17687_, _17686_);
  and (_17689_, _17688_, _06114_);
  and (_17690_, _17689_, _17685_);
  and (_17691_, _14630_, _07809_);
  or (_17692_, _17691_, _17549_);
  and (_17693_, _17692_, _05787_);
  or (_17694_, _17693_, _09855_);
  or (_17695_, _17694_, _17690_);
  or (_17696_, _10052_, _09861_);
  and (_17697_, _17696_, _05802_);
  and (_17698_, _17697_, _17695_);
  nor (_17699_, _06625_, _05802_);
  or (_17700_, _17699_, _06110_);
  or (_17701_, _17700_, _17698_);
  and (_17702_, _07809_, _08768_);
  or (_17703_, _17702_, _17549_);
  or (_17704_, _17703_, _06111_);
  and (_17705_, _17704_, _10752_);
  and (_17706_, _17705_, _17701_);
  or (_17707_, _17706_, _17553_);
  and (_17708_, _17707_, _10762_);
  and (_17709_, _06957_, _06399_);
  or (_17710_, _17709_, _06574_);
  and (_17711_, _10980_, _06558_);
  or (_17712_, _17711_, _17710_);
  or (_17713_, _17712_, _17708_);
  and (_17714_, _06684_, _06399_);
  nor (_17715_, _10772_, _17714_);
  nand (_17716_, _17710_, _10981_);
  and (_17717_, _17716_, _17715_);
  and (_17718_, _17717_, _17713_);
  nor (_17719_, _17715_, _10981_);
  or (_17720_, _17719_, _10775_);
  or (_17721_, _17720_, _17718_);
  and (_17722_, _17721_, _17552_);
  or (_17723_, _17722_, _06400_);
  or (_17724_, _10282_, _06401_);
  and (_17725_, _17724_, _10788_);
  and (_17726_, _17725_, _17723_);
  and (_17727_, _10787_, _11063_);
  or (_17728_, _17727_, _06297_);
  or (_17729_, _17728_, _17726_);
  and (_17730_, _17729_, _17551_);
  or (_17731_, _17730_, _06402_);
  or (_17732_, _17549_, _07125_);
  and (_17733_, _17732_, _10808_);
  and (_17734_, _17733_, _17731_);
  and (_17735_, _10812_, _10978_);
  or (_17736_, _17735_, _10811_);
  or (_17737_, _17736_, _17734_);
  or (_17738_, _10816_, _11018_);
  and (_17739_, _17738_, _06410_);
  and (_17740_, _17739_, _17737_);
  or (_17741_, _10820_, _10274_);
  and (_17742_, _17741_, _10822_);
  or (_17743_, _17742_, _17740_);
  or (_17744_, _10826_, _11061_);
  and (_17745_, _17744_, _07132_);
  and (_17746_, _17745_, _17743_);
  nand (_17747_, _17703_, _06306_);
  nor (_17748_, _17747_, _10281_);
  or (_17749_, _17748_, _17546_);
  or (_17750_, _17749_, _17746_);
  nand (_17751_, _17750_, _17547_);
  nor (_17752_, _17156_, _17148_);
  nand (_17753_, _17752_, _17751_);
  not (_17754_, _17752_);
  nand (_17755_, _17754_, _10979_);
  and (_17756_, _17755_, _17161_);
  and (_17757_, _17756_, _17753_);
  nor (_17758_, _10979_, _17161_);
  or (_17759_, _17758_, _10841_);
  or (_17760_, _17759_, _17757_);
  or (_17761_, _17242_, _11019_);
  and (_17762_, _17761_, _06395_);
  and (_17763_, _17762_, _17760_);
  nand (_17764_, _10851_, _10281_);
  and (_17765_, _17764_, _10850_);
  or (_17766_, _17765_, _17763_);
  and (_17767_, _17766_, _17545_);
  or (_17768_, _17767_, _06303_);
  and (_17769_, _14643_, _07809_);
  or (_17770_, _17549_, _08819_);
  or (_17771_, _17770_, _17769_);
  and (_17772_, _17771_, _10380_);
  and (_17773_, _17772_, _17768_);
  or (_17774_, _17773_, _17544_);
  and (_17775_, _17774_, _17241_);
  and (_17776_, _10878_, _10619_);
  nor (_17777_, _17776_, _10879_);
  and (_17778_, _17777_, _17240_);
  or (_17779_, _17778_, _17775_);
  or (_17780_, _17779_, _06792_);
  or (_17781_, _17777_, _06793_);
  and (_17782_, _17781_, _06407_);
  and (_17783_, _17782_, _17780_);
  or (_17784_, _17783_, _17541_);
  nand (_17785_, _17784_, _10927_);
  and (_17786_, _10938_, _10691_);
  or (_17787_, _10939_, _10927_);
  or (_17788_, _17787_, _17786_);
  and (_17789_, _17788_, _10926_);
  and (_17790_, _17789_, _17785_);
  nand (_17791_, _10925_, _05887_);
  nand (_17792_, _17791_, _10963_);
  or (_17793_, _17792_, _17790_);
  and (_17794_, _10987_, _10981_);
  or (_17795_, _17794_, _10988_);
  or (_17796_, _17795_, _10963_);
  and (_17797_, _17796_, _17201_);
  and (_17798_, _17797_, _17793_);
  and (_17799_, _11029_, _11022_);
  or (_17800_, _17799_, _11030_);
  or (_17801_, _17800_, _05707_);
  and (_17802_, _17801_, _11003_);
  nor (_17803_, _17802_, _17798_);
  or (_17804_, _17800_, _17200_);
  nand (_17805_, _17804_, _06171_);
  or (_17806_, _17805_, _17803_);
  and (_17807_, _17806_, _17538_);
  or (_17808_, _11070_, _11063_);
  nor (_17809_, _11071_, _10265_);
  and (_17810_, _17809_, _17808_);
  or (_17811_, _17810_, _10262_);
  or (_17812_, _17811_, _17807_);
  and (_17813_, _17812_, _17534_);
  or (_17814_, _17813_, _06433_);
  or (_17815_, _17577_, _06829_);
  and (_17816_, _17815_, _11090_);
  and (_17817_, _17816_, _17814_);
  nor (_17818_, _17511_, _09981_);
  or (_17819_, _17818_, _11095_);
  nor (_17820_, _17819_, _11094_);
  nor (_17821_, _17820_, _12719_);
  or (_17822_, _17821_, _17817_);
  nand (_17823_, _11094_, _10028_);
  and (_17824_, _17823_, _05749_);
  and (_17825_, _17824_, _17822_);
  and (_17826_, _17615_, _05748_);
  or (_17827_, _17826_, _06440_);
  or (_17828_, _17827_, _17825_);
  and (_17829_, _14710_, _07809_);
  or (_17830_, _17829_, _17549_);
  or (_17831_, _17830_, _06444_);
  and (_17832_, _17831_, _11113_);
  and (_17833_, _17832_, _17828_);
  nor (_17834_, _11120_, \oc8051_golden_model_1.ACC [2]);
  nor (_17835_, _17834_, _11121_);
  and (_17836_, _17835_, _11112_);
  or (_17837_, _17836_, _11119_);
  or (_17838_, _17837_, _17833_);
  nand (_17839_, _11119_, _10028_);
  and (_17840_, _17839_, _01317_);
  and (_17841_, _17840_, _17838_);
  or (_17842_, _17841_, _17533_);
  and (_43605_, _17842_, _43100_);
  nor (_17843_, _01317_, _10028_);
  and (_17844_, _10359_, _10337_);
  nor (_17845_, _17844_, _10360_);
  or (_17846_, _17845_, _10380_);
  not (_17847_, _10835_);
  nor (_17848_, _17847_, _10977_);
  or (_17849_, _17848_, _10841_);
  nand (_17850_, _10977_, _06524_);
  and (_17851_, _10976_, _06965_);
  and (_17852_, _17407_, _10976_);
  and (_17853_, _14727_, _07809_);
  nor (_17854_, _07809_, _10028_);
  or (_17855_, _17854_, _07127_);
  or (_17856_, _17855_, _17853_);
  nor (_17857_, _10752_, _06070_);
  and (_17858_, _07809_, _07544_);
  or (_17859_, _17858_, _17854_);
  or (_17860_, _17859_, _06132_);
  or (_17861_, _10458_, _07544_);
  nor (_17862_, _08409_, _10028_);
  and (_17863_, _14735_, _08409_);
  or (_17864_, _17863_, _17862_);
  or (_17865_, _17864_, _06157_);
  and (_17866_, _17865_, _07075_);
  and (_17867_, _14738_, _07809_);
  or (_17868_, _17867_, _17854_);
  and (_17869_, _17868_, _06160_);
  or (_17870_, _17009_, _09210_);
  and (_17871_, _17011_, _07544_);
  or (_17872_, _06653_, \oc8051_golden_model_1.ACC [3]);
  nand (_17873_, _06653_, \oc8051_golden_model_1.ACC [3]);
  and (_17874_, _17873_, _17872_);
  and (_17875_, _17874_, _10471_);
  or (_17876_, _17875_, _10473_);
  or (_17877_, _17876_, _17871_);
  and (_17878_, _17877_, _05772_);
  or (_17879_, _17878_, _07064_);
  and (_17880_, _17879_, _06161_);
  and (_17881_, _17880_, _17870_);
  or (_17882_, _17881_, _17869_);
  and (_17883_, _17882_, _10491_);
  not (_17884_, \oc8051_golden_model_1.PSW [6]);
  nor (_17885_, _10493_, _17884_);
  nor (_17886_, _17885_, \oc8051_golden_model_1.ACC [3]);
  nor (_17887_, _17886_, _10494_);
  and (_17888_, _17887_, _10490_);
  or (_17889_, _17888_, _06156_);
  or (_17890_, _17889_, _17883_);
  and (_17891_, _17890_, _17866_);
  and (_17892_, _17859_, _06217_);
  or (_17893_, _17892_, _10516_);
  or (_17894_, _17893_, _17891_);
  and (_17895_, _17894_, _17861_);
  or (_17896_, _17895_, _07081_);
  or (_17897_, _09210_, _07082_);
  and (_17898_, _17897_, _06229_);
  and (_17899_, _17898_, _17896_);
  nor (_17900_, _08139_, _06229_);
  or (_17901_, _17900_, _10525_);
  or (_17902_, _17901_, _17899_);
  nand (_17903_, _10525_, _08430_);
  and (_17904_, _17903_, _17902_);
  or (_17905_, _17904_, _06152_);
  and (_17906_, _14731_, _08409_);
  or (_17907_, _17906_, _17862_);
  or (_17908_, _17907_, _06153_);
  and (_17909_, _17908_, _06146_);
  and (_17910_, _17909_, _17905_);
  or (_17911_, _17862_, _14764_);
  and (_17912_, _17864_, _06145_);
  and (_17913_, _17912_, _17911_);
  or (_17914_, _17913_, _09295_);
  or (_17915_, _17914_, _17910_);
  nor (_17916_, _09777_, _09775_);
  or (_17917_, _17916_, _09778_);
  nand (_17918_, _17917_, _09295_);
  and (_17919_, _17918_, _10554_);
  and (_17920_, _17919_, _17915_);
  and (_17921_, _07657_, \oc8051_golden_model_1.ACC [2]);
  nor (_17922_, _17633_, _17921_);
  nor (_17923_, _10976_, _10977_);
  nor (_17924_, _17923_, _17922_);
  and (_17925_, _17923_, _17922_);
  nor (_17926_, _17925_, _17924_);
  not (_17927_, _17636_);
  nor (_17928_, _17927_, _17635_);
  nand (_17929_, _17928_, \oc8051_golden_model_1.PSW [7]);
  and (_17930_, _17929_, _17926_);
  not (_17931_, _17928_);
  nor (_17932_, _17931_, _17926_);
  and (_17933_, _17932_, \oc8051_golden_model_1.PSW [7]);
  or (_17934_, _17933_, _17930_);
  and (_17935_, _17934_, _10557_);
  or (_17936_, _17935_, _12379_);
  or (_17937_, _17936_, _17920_);
  and (_17938_, _09070_, \oc8051_golden_model_1.ACC [2]);
  nor (_17939_, _17648_, _17938_);
  nor (_17940_, _11016_, _11017_);
  not (_17941_, _17940_);
  nand (_17942_, _17941_, _17939_);
  or (_17943_, _17941_, _17939_);
  and (_17944_, _17943_, _17942_);
  or (_17945_, _17944_, _10693_);
  nand (_17946_, _17944_, _10693_);
  and (_17947_, _17946_, _17945_);
  nand (_17948_, _17947_, _17654_);
  or (_17949_, _17947_, _17654_);
  and (_17950_, _17949_, _17948_);
  or (_17951_, _17950_, _12380_);
  and (_17952_, _17951_, _06265_);
  and (_17953_, _17952_, _17937_);
  and (_17954_, _12324_, \oc8051_golden_model_1.PSW [7]);
  and (_17955_, _08247_, \oc8051_golden_model_1.ACC [2]);
  nor (_17956_, _17561_, _17955_);
  nor (_17957_, _17956_, _12318_);
  and (_17958_, _17956_, _12318_);
  nor (_17959_, _17958_, _17957_);
  not (_17960_, _12323_);
  or (_17961_, _17960_, _17563_);
  or (_17962_, _17961_, _10693_);
  and (_17963_, _17962_, _17959_);
  or (_17964_, _17963_, _10387_);
  or (_17965_, _17964_, _17954_);
  and (_17966_, _17965_, _12386_);
  or (_17967_, _17966_, _17953_);
  and (_17968_, _12341_, \oc8051_golden_model_1.PSW [7]);
  and (_17969_, _06625_, \oc8051_golden_model_1.ACC [2]);
  nor (_17970_, _17667_, _17969_);
  nor (_17971_, _12336_, _17970_);
  and (_17972_, _12336_, _17970_);
  nor (_17973_, _17972_, _17971_);
  not (_17974_, _12340_);
  or (_17975_, _17974_, _17669_);
  or (_17976_, _17975_, _10693_);
  and (_17977_, _17976_, _17973_);
  or (_17978_, _17977_, _10388_);
  or (_17979_, _17978_, _17968_);
  and (_17980_, _17979_, _17967_);
  or (_17981_, _17980_, _05870_);
  nand (_17982_, _06070_, _05870_);
  and (_17983_, _17982_, _06140_);
  and (_17984_, _17983_, _17981_);
  and (_17985_, _14732_, _08409_);
  or (_17986_, _17985_, _17862_);
  and (_17987_, _17986_, _06139_);
  or (_17988_, _17987_, _09842_);
  or (_17989_, _17988_, _17984_);
  and (_17990_, _17989_, _17860_);
  or (_17991_, _17990_, _06116_);
  and (_17992_, _09210_, _07809_);
  or (_17993_, _17854_, _06117_);
  or (_17994_, _17993_, _17992_);
  and (_17995_, _17994_, _06114_);
  and (_17996_, _17995_, _17991_);
  and (_17997_, _14825_, _07809_);
  or (_17998_, _17997_, _17854_);
  and (_17999_, _17998_, _05787_);
  or (_18001_, _17999_, _09855_);
  or (_18002_, _18001_, _17996_);
  or (_18003_, _09998_, _09861_);
  and (_18004_, _18003_, _05802_);
  and (_18005_, _18004_, _18002_);
  nor (_18006_, _06070_, _05802_);
  or (_18007_, _18006_, _06110_);
  or (_18008_, _18007_, _18005_);
  and (_18009_, _07809_, _08712_);
  or (_18010_, _18009_, _17854_);
  or (_18011_, _18010_, _06111_);
  and (_18012_, _18011_, _10752_);
  and (_18013_, _18012_, _18008_);
  or (_18014_, _18013_, _17857_);
  and (_18015_, _18014_, _10762_);
  and (_18016_, _17923_, _06558_);
  or (_18017_, _18016_, _17109_);
  or (_18018_, _18017_, _18015_);
  or (_18019_, _17106_, _17923_);
  and (_18020_, _18019_, _17113_);
  and (_18021_, _18020_, _18018_);
  and (_18022_, _17923_, _06771_);
  or (_18023_, _18022_, _18021_);
  and (_18024_, _18023_, _10776_);
  and (_18025_, _10775_, _17940_);
  or (_18026_, _18025_, _06400_);
  or (_18027_, _18026_, _18024_);
  or (_18028_, _12318_, _06401_);
  and (_18029_, _18028_, _10788_);
  and (_18030_, _18029_, _18027_);
  and (_18031_, _10787_, _12336_);
  or (_18032_, _18031_, _06297_);
  or (_18033_, _18032_, _18030_);
  and (_18034_, _18033_, _17856_);
  or (_18035_, _18034_, _06402_);
  or (_18036_, _17854_, _07125_);
  and (_18037_, _18036_, _17408_);
  and (_18038_, _18037_, _18035_);
  or (_18039_, _18038_, _17852_);
  and (_18040_, _18039_, _17417_);
  or (_18041_, _18040_, _17851_);
  and (_18042_, _18041_, _17416_);
  and (_18043_, _10807_, _10976_);
  or (_18044_, _18043_, _10811_);
  or (_18045_, _18044_, _18042_);
  or (_18046_, _10816_, _11016_);
  and (_18047_, _18046_, _06410_);
  and (_18048_, _18047_, _18045_);
  and (_18049_, _10272_, _06409_);
  or (_18050_, _18049_, _10820_);
  or (_18051_, _18050_, _18048_);
  or (_18052_, _10826_, _11059_);
  and (_18053_, _18052_, _07132_);
  and (_18054_, _18053_, _18051_);
  nand (_18055_, _18010_, _06306_);
  nor (_18056_, _18055_, _10273_);
  or (_18057_, _18056_, _06524_);
  or (_18058_, _18057_, _18054_);
  and (_18059_, _18058_, _17850_);
  or (_18060_, _18059_, _06555_);
  nand (_18061_, _10977_, _06555_);
  and (_18062_, _18061_, _18060_);
  or (_18063_, _18062_, _06975_);
  nand (_18064_, _10977_, _06975_);
  and (_18065_, _18064_, _17847_);
  and (_18066_, _18065_, _18063_);
  or (_18067_, _18066_, _17849_);
  nand (_18068_, _10841_, _11017_);
  and (_18069_, _18068_, _06395_);
  and (_18070_, _18069_, _18067_);
  nand (_18071_, _10851_, _10273_);
  and (_18072_, _18071_, _10850_);
  or (_18073_, _18072_, _18070_);
  nand (_18074_, _10848_, _11060_);
  and (_18075_, _18074_, _08819_);
  and (_18076_, _18075_, _18073_);
  and (_18077_, _14724_, _07809_);
  or (_18078_, _18077_, _17854_);
  and (_18079_, _18078_, _06303_);
  or (_18080_, _18079_, _10858_);
  or (_18081_, _18080_, _18076_);
  and (_18082_, _18081_, _17846_);
  or (_18083_, _18082_, _10865_);
  and (_18084_, _10880_, _10613_);
  nor (_18085_, _18084_, _10881_);
  or (_18086_, _18085_, _10867_);
  and (_18087_, _18086_, _06407_);
  and (_18088_, _18087_, _18083_);
  nand (_18089_, _10910_, _10422_);
  nor (_18090_, _10911_, _06407_);
  and (_18091_, _18090_, _18089_);
  or (_18092_, _18091_, _10895_);
  or (_18093_, _18092_, _18088_);
  and (_18094_, _10940_, _10685_);
  nor (_18095_, _18094_, _10941_);
  or (_18096_, _18095_, _10927_);
  and (_18097_, _18096_, _10926_);
  and (_18098_, _18097_, _18093_);
  nand (_18099_, _10925_, \oc8051_golden_model_1.ACC [2]);
  nand (_18100_, _18099_, _10963_);
  or (_18101_, _18100_, _18098_);
  and (_18102_, _10989_, _17923_);
  nor (_18103_, _10989_, _17923_);
  or (_18104_, _18103_, _18102_);
  or (_18105_, _18104_, _10963_);
  and (_18106_, _18105_, _18101_);
  or (_18107_, _18106_, _11003_);
  and (_18108_, _11031_, _17940_);
  nor (_18109_, _11031_, _17940_);
  or (_18110_, _18109_, _11041_);
  or (_18111_, _18110_, _18108_);
  and (_18112_, _18111_, _06171_);
  and (_18113_, _18112_, _18107_);
  and (_18114_, _12318_, _10285_);
  nor (_18115_, _12318_, _10285_);
  or (_18116_, _18115_, _10264_);
  or (_18117_, _18116_, _18114_);
  and (_18118_, _18117_, _12691_);
  or (_18119_, _18118_, _18113_);
  and (_18120_, _11072_, _12336_);
  nor (_18121_, _11072_, _12336_);
  or (_18122_, _18121_, _18120_);
  or (_18123_, _18122_, _10265_);
  and (_18124_, _18123_, _12693_);
  and (_18125_, _18124_, _18119_);
  and (_18126_, _10262_, \oc8051_golden_model_1.ACC [2]);
  or (_18127_, _18126_, _06433_);
  or (_18128_, _18127_, _18125_);
  or (_18129_, _17868_, _06829_);
  and (_18130_, _18129_, _11090_);
  and (_18131_, _18130_, _18128_);
  nor (_18132_, _11095_, _10028_);
  or (_18133_, _18132_, _11096_);
  and (_18134_, _18133_, _11089_);
  or (_18135_, _18134_, _11094_);
  or (_18136_, _18135_, _18131_);
  nand (_18137_, _11094_, _09902_);
  and (_18138_, _18137_, _05749_);
  and (_18139_, _18138_, _18136_);
  and (_18140_, _17907_, _05748_);
  or (_18141_, _18140_, _06440_);
  or (_18142_, _18141_, _18139_);
  and (_18143_, _14897_, _07809_);
  or (_18144_, _17854_, _06444_);
  or (_18145_, _18144_, _18143_);
  and (_18146_, _18145_, _11113_);
  and (_18147_, _18146_, _18142_);
  nor (_18148_, _11121_, \oc8051_golden_model_1.ACC [3]);
  nor (_18149_, _18148_, _11122_);
  and (_18150_, _18149_, _11112_);
  or (_18151_, _18150_, _11119_);
  or (_18152_, _18151_, _18147_);
  nand (_18153_, _11119_, _09902_);
  and (_18154_, _18153_, _01317_);
  and (_18155_, _18154_, _18152_);
  or (_18156_, _18155_, _17843_);
  and (_43606_, _18156_, _43100_);
  nor (_18157_, _01317_, _09902_);
  nand (_18158_, _10262_, _10028_);
  or (_18159_, _10289_, _10287_);
  and (_18160_, _10290_, _06169_);
  and (_18161_, _18160_, _18159_);
  or (_18162_, _11033_, _11015_);
  and (_18163_, _18162_, _11034_);
  or (_18164_, _18163_, _17201_);
  or (_18165_, _10912_, _10416_);
  and (_18166_, _18165_, _10913_);
  or (_18167_, _18166_, _06407_);
  and (_18168_, _18167_, _10927_);
  nand (_18169_, _10848_, _11057_);
  or (_18170_, _06965_, _06554_);
  and (_18171_, _18170_, _10972_);
  not (_18172_, _17105_);
  and (_18173_, _18172_, _06772_);
  nor (_18174_, _06722_, _05833_);
  and (_18175_, _06123_, _06399_);
  nor (_18176_, _18175_, _18174_);
  not (_18177_, _18176_);
  and (_18178_, _06128_, _06399_);
  nor (_18179_, _18178_, _18177_);
  and (_18180_, _18179_, _18173_);
  and (_18181_, _06277_, _06399_);
  not (_18182_, _18181_);
  nor (_18183_, _10752_, _06876_);
  nor (_18184_, _07809_, _09902_);
  and (_18185_, _08336_, _07809_);
  or (_18186_, _18185_, _18184_);
  or (_18187_, _18186_, _06132_);
  nand (_18188_, _17948_, _17945_);
  and (_18189_, _09210_, _10028_);
  or (_18191_, _09210_, _10028_);
  and (_18192_, _18191_, _17939_);
  or (_18193_, _18192_, _18189_);
  nor (_18194_, _11015_, _18193_);
  not (_18195_, _18194_);
  nand (_18196_, _11015_, _18193_);
  and (_18197_, _18196_, _18195_);
  nand (_18198_, _18197_, \oc8051_golden_model_1.PSW [7]);
  or (_18199_, _18197_, \oc8051_golden_model_1.PSW [7]);
  and (_18200_, _18199_, _18198_);
  or (_18202_, _18200_, _18188_);
  nand (_18203_, _18200_, _18188_);
  and (_18204_, _12379_, _18203_);
  and (_18205_, _18204_, _18202_);
  nor (_18206_, _17932_, _10693_);
  and (_18207_, _07544_, _10028_);
  or (_18208_, _07544_, _10028_);
  and (_18209_, _18208_, _17922_);
  or (_18210_, _18209_, _18207_);
  nor (_18211_, _10975_, _18210_);
  and (_18213_, _10975_, _18210_);
  nor (_18214_, _18213_, _18211_);
  and (_18215_, _18214_, \oc8051_golden_model_1.PSW [7]);
  nor (_18216_, _18214_, \oc8051_golden_model_1.PSW [7]);
  nor (_18217_, _18216_, _18215_);
  and (_18218_, _18217_, _18206_);
  nor (_18219_, _18217_, _18206_);
  nor (_18220_, _18219_, _18218_);
  and (_18221_, _18220_, _10557_);
  or (_18222_, _10458_, _08336_);
  nor (_18224_, _08409_, _09902_);
  and (_18225_, _14932_, _08409_);
  or (_18226_, _18225_, _18224_);
  or (_18227_, _18226_, _06157_);
  and (_18228_, _18227_, _07075_);
  and (_18229_, _14928_, _07809_);
  or (_18230_, _18229_, _18184_);
  and (_18231_, _18230_, _06160_);
  or (_18232_, _10474_, _09209_);
  and (_18233_, _17011_, _08336_);
  or (_18235_, _06653_, \oc8051_golden_model_1.ACC [4]);
  nand (_18236_, _06653_, \oc8051_golden_model_1.ACC [4]);
  and (_18237_, _18236_, _18235_);
  and (_18238_, _18237_, _10471_);
  or (_18239_, _18238_, _10473_);
  or (_18240_, _18239_, _18233_);
  and (_18241_, _18240_, _10484_);
  and (_18242_, _18241_, _18232_);
  or (_18243_, _18242_, _18231_);
  and (_18244_, _18243_, _10491_);
  nor (_18246_, _10494_, \oc8051_golden_model_1.ACC [4]);
  nor (_18247_, _18246_, _10495_);
  and (_18248_, _18247_, _10490_);
  or (_18249_, _18248_, _06156_);
  or (_18250_, _18249_, _18244_);
  and (_18251_, _18250_, _18228_);
  and (_18252_, _18186_, _06217_);
  or (_18253_, _18252_, _10516_);
  or (_18254_, _18253_, _18251_);
  and (_18255_, _18254_, _18222_);
  or (_18257_, _18255_, _07081_);
  or (_18258_, _09209_, _07082_);
  and (_18259_, _18258_, _06229_);
  and (_18260_, _18259_, _18257_);
  nor (_18261_, _08338_, _06229_);
  or (_18262_, _18261_, _10525_);
  or (_18263_, _18262_, _18260_);
  nand (_18264_, _10525_, _05855_);
  and (_18265_, _18264_, _18263_);
  or (_18266_, _18265_, _06152_);
  and (_18268_, _14942_, _08409_);
  or (_18269_, _18268_, _18224_);
  or (_18270_, _18269_, _06153_);
  and (_18271_, _18270_, _06146_);
  and (_18272_, _18271_, _18266_);
  or (_18273_, _18224_, _14949_);
  and (_18274_, _18226_, _06145_);
  and (_18275_, _18274_, _18273_);
  or (_18276_, _18275_, _09295_);
  or (_18277_, _18276_, _18272_);
  nor (_18279_, _09780_, _09778_);
  nor (_18280_, _18279_, _09781_);
  or (_18281_, _18280_, _09301_);
  and (_18282_, _18281_, _10554_);
  and (_18283_, _18282_, _18277_);
  or (_18284_, _18283_, _18221_);
  and (_18285_, _18284_, _12380_);
  or (_18286_, _18285_, _18205_);
  and (_18287_, _18286_, _06265_);
  nor (_18288_, _12324_, _10693_);
  or (_18290_, _17956_, _13917_);
  and (_18291_, _18290_, _13915_);
  nor (_18292_, _18291_, _10289_);
  and (_18293_, _18291_, _10289_);
  nor (_18294_, _18293_, _18292_);
  and (_18295_, _18294_, \oc8051_golden_model_1.PSW [7]);
  nor (_18296_, _18294_, \oc8051_golden_model_1.PSW [7]);
  nor (_18297_, _18296_, _18295_);
  or (_18298_, _18297_, _18288_);
  and (_18299_, _18297_, _18288_);
  nor (_18301_, _18299_, _06265_);
  and (_18302_, _18301_, _18298_);
  or (_18303_, _18302_, _18287_);
  and (_18304_, _18303_, _10388_);
  nor (_18305_, _12341_, _10693_);
  or (_18306_, _17970_, _13950_);
  and (_18307_, _18306_, _13949_);
  nor (_18308_, _11058_, _18307_);
  and (_18309_, _11058_, _18307_);
  nor (_18310_, _18309_, _18308_);
  and (_18312_, _18310_, \oc8051_golden_model_1.PSW [7]);
  nor (_18313_, _18310_, \oc8051_golden_model_1.PSW [7]);
  nor (_18314_, _18313_, _18312_);
  or (_18315_, _18314_, _18305_);
  and (_18316_, _18314_, _18305_);
  nor (_18317_, _18316_, _10388_);
  and (_18318_, _18317_, _18315_);
  or (_18319_, _18318_, _05870_);
  or (_18320_, _18319_, _18304_);
  nand (_18321_, _06876_, _05870_);
  and (_18323_, _18321_, _06140_);
  and (_18324_, _18323_, _18320_);
  and (_18325_, _14966_, _08409_);
  or (_18326_, _18325_, _18224_);
  and (_18327_, _18326_, _06139_);
  or (_18328_, _18327_, _09842_);
  or (_18329_, _18328_, _18324_);
  and (_18330_, _18329_, _18187_);
  or (_18331_, _18330_, _06116_);
  and (_18332_, _09209_, _07809_);
  or (_18334_, _18184_, _06117_);
  or (_18335_, _18334_, _18332_);
  and (_18336_, _18335_, _06114_);
  and (_18337_, _18336_, _18331_);
  and (_18338_, _15013_, _07809_);
  or (_18339_, _18338_, _18184_);
  and (_18340_, _18339_, _05787_);
  or (_18341_, _18340_, _09855_);
  or (_18342_, _18341_, _18337_);
  or (_18343_, _09947_, _09861_);
  and (_18345_, _18343_, _05802_);
  and (_18346_, _18345_, _18342_);
  nor (_18347_, _06876_, _05802_);
  or (_18348_, _18347_, _06110_);
  or (_18349_, _18348_, _18346_);
  and (_18350_, _08715_, _07809_);
  or (_18351_, _18350_, _18184_);
  or (_18352_, _18351_, _06111_);
  and (_18353_, _18352_, _10752_);
  and (_18354_, _18353_, _18349_);
  or (_18356_, _18354_, _18183_);
  and (_18357_, _18356_, _18182_);
  and (_18358_, _10975_, _18181_);
  nor (_18359_, _18358_, _18357_);
  nand (_18360_, _18359_, _18180_);
  or (_18361_, _18180_, _10975_);
  and (_18362_, _18361_, _10776_);
  and (_18363_, _18362_, _18360_);
  and (_18364_, _10775_, _11015_);
  or (_18365_, _18364_, _06400_);
  or (_18366_, _18365_, _18363_);
  or (_18367_, _10289_, _06401_);
  and (_18368_, _18367_, _18366_);
  and (_18369_, _18368_, _10788_);
  and (_18370_, _10787_, _11058_);
  or (_18371_, _18370_, _06297_);
  or (_18372_, _18371_, _18369_);
  and (_18373_, _15029_, _07809_);
  or (_18374_, _18184_, _07127_);
  or (_18375_, _18374_, _18373_);
  and (_18377_, _18375_, _07125_);
  and (_18378_, _18377_, _18372_);
  and (_18379_, _18184_, _06402_);
  or (_18380_, _18379_, _06557_);
  or (_18381_, _18380_, _18378_);
  and (_18382_, _10972_, _05742_);
  or (_18383_, _18382_, _17408_);
  and (_18384_, _18383_, _17417_);
  and (_18385_, _18384_, _18381_);
  or (_18386_, _18385_, _18171_);
  and (_18388_, _18386_, _17416_);
  and (_18389_, _10807_, _10972_);
  or (_18390_, _18389_, _10811_);
  or (_18391_, _18390_, _18388_);
  or (_18392_, _10816_, _11012_);
  and (_18393_, _18392_, _06410_);
  and (_18394_, _18393_, _18391_);
  or (_18395_, _10820_, _10270_);
  and (_18396_, _18395_, _10822_);
  or (_18397_, _18396_, _18394_);
  or (_18399_, _10826_, _11055_);
  and (_18400_, _18399_, _07132_);
  and (_18401_, _18400_, _18397_);
  nand (_18402_, _18351_, _06306_);
  nor (_18403_, _18402_, _10288_);
  or (_18404_, _18403_, _06524_);
  or (_18405_, _18404_, _18401_);
  not (_18406_, _06524_);
  or (_18407_, _10973_, _18406_);
  and (_18408_, _18407_, _10837_);
  and (_18410_, _18408_, _18405_);
  not (_18411_, _10837_);
  and (_18412_, _18411_, _10973_);
  or (_18413_, _18412_, _10841_);
  or (_18414_, _18413_, _18410_);
  or (_18415_, _17242_, _11014_);
  and (_18416_, _18415_, _06395_);
  and (_18417_, _18416_, _18414_);
  nand (_18418_, _10851_, _10288_);
  and (_18419_, _18418_, _10850_);
  or (_18421_, _18419_, _18417_);
  and (_18422_, _18421_, _18169_);
  or (_18423_, _18422_, _06303_);
  and (_18424_, _15026_, _07809_);
  or (_18425_, _18184_, _08819_);
  or (_18426_, _18425_, _18424_);
  and (_18427_, _18426_, _10380_);
  and (_18428_, _18427_, _18423_);
  or (_18429_, _10361_, _10330_);
  and (_18430_, _18429_, _10362_);
  and (_18432_, _18430_, _10858_);
  or (_18433_, _18432_, _17240_);
  or (_18434_, _18433_, _18428_);
  or (_18435_, _10882_, _10606_);
  and (_18436_, _18435_, _10883_);
  and (_18437_, _18436_, _06276_);
  or (_18438_, _18437_, _10867_);
  and (_18439_, _18438_, _18434_);
  and (_18440_, _18436_, _06792_);
  or (_18441_, _18440_, _06406_);
  or (_18443_, _18441_, _18439_);
  and (_18444_, _18443_, _18168_);
  or (_18445_, _10942_, _10679_);
  and (_18446_, _10943_, _10895_);
  and (_18447_, _18446_, _18445_);
  or (_18448_, _18447_, _10925_);
  or (_18449_, _18448_, _18444_);
  nand (_18450_, _10925_, _10028_);
  and (_18451_, _18450_, _10963_);
  and (_18452_, _18451_, _18449_);
  not (_18454_, _10963_);
  nor (_18455_, _10991_, _10975_);
  nor (_18456_, _18455_, _10992_);
  and (_18457_, _18456_, _18454_);
  or (_18458_, _18457_, _17195_);
  or (_18459_, _18458_, _18452_);
  and (_18460_, _18459_, _18164_);
  or (_18461_, _18460_, _17199_);
  or (_18462_, _18163_, _17200_);
  and (_18463_, _18462_, _06171_);
  and (_18465_, _18463_, _18461_);
  or (_18466_, _18465_, _18161_);
  and (_18467_, _18466_, _10265_);
  or (_18468_, _11074_, _11058_);
  and (_18469_, _11075_, _10264_);
  and (_18470_, _18469_, _18468_);
  or (_18471_, _18470_, _10262_);
  or (_18472_, _18471_, _18467_);
  and (_18473_, _18472_, _18158_);
  or (_18474_, _18473_, _06433_);
  or (_18476_, _18230_, _06829_);
  and (_18477_, _18476_, _11090_);
  and (_18478_, _18477_, _18474_);
  nor (_18479_, _11096_, _09902_);
  or (_18480_, _18479_, _11097_);
  and (_18481_, _18480_, _11089_);
  or (_18482_, _18481_, _11094_);
  or (_18483_, _18482_, _18478_);
  nand (_18484_, _11094_, _09930_);
  and (_18485_, _18484_, _05749_);
  and (_18487_, _18485_, _18483_);
  and (_18488_, _18269_, _05748_);
  or (_18489_, _18488_, _06440_);
  or (_18490_, _18489_, _18487_);
  and (_18491_, _15087_, _07809_);
  or (_18492_, _18184_, _06444_);
  or (_18493_, _18492_, _18491_);
  and (_18494_, _18493_, _11113_);
  and (_18495_, _18494_, _18490_);
  nor (_18496_, _11122_, \oc8051_golden_model_1.ACC [4]);
  nor (_18498_, _18496_, _11123_);
  and (_18499_, _18498_, _11112_);
  or (_18500_, _18499_, _11119_);
  or (_18501_, _18500_, _18495_);
  nand (_18502_, _11119_, _09930_);
  and (_18503_, _18502_, _01317_);
  and (_18504_, _18503_, _18501_);
  or (_18505_, _18504_, _18157_);
  and (_43607_, _18505_, _43100_);
  nor (_18506_, _01317_, _09930_);
  and (_18508_, _10363_, _10323_);
  nor (_18509_, _18508_, _10364_);
  or (_18510_, _18509_, _10380_);
  and (_18511_, _15219_, _07809_);
  nor (_18512_, _07809_, _09930_);
  or (_18513_, _18512_, _07127_);
  or (_18514_, _18513_, _18511_);
  nor (_18515_, _10971_, _10970_);
  nor (_18516_, _18178_, _10772_);
  not (_18517_, _18516_);
  and (_18519_, _18517_, _18515_);
  nor (_18520_, _10752_, _06477_);
  and (_18521_, _08101_, _07809_);
  or (_18522_, _18521_, _18512_);
  or (_18523_, _18522_, _06132_);
  and (_18524_, _06876_, \oc8051_golden_model_1.ACC [4]);
  nor (_18525_, _18308_, _18524_);
  nor (_18526_, _12342_, _18525_);
  and (_18527_, _12342_, _18525_);
  nor (_18528_, _18527_, _18526_);
  and (_18530_, _18528_, \oc8051_golden_model_1.PSW [7]);
  nor (_18531_, _18528_, \oc8051_golden_model_1.PSW [7]);
  nor (_18532_, _18531_, _18530_);
  nor (_18533_, _18316_, _18312_);
  not (_18534_, _18533_);
  and (_18535_, _18534_, _18532_);
  nor (_18536_, _18534_, _18532_);
  nor (_18537_, _18536_, _18535_);
  or (_18538_, _18537_, _10388_);
  and (_18539_, _08980_, \oc8051_golden_model_1.ACC [4]);
  nor (_18541_, _18194_, _18539_);
  or (_18542_, _11011_, _18541_);
  nand (_18543_, _11011_, _18541_);
  and (_18544_, _18543_, _18542_);
  or (_18545_, _18544_, _10693_);
  nand (_18546_, _18544_, _10693_);
  and (_18547_, _18546_, _18545_);
  nand (_18548_, _18203_, _18198_);
  nand (_18549_, _18548_, _18547_);
  or (_18550_, _18548_, _18547_);
  and (_18552_, _18550_, _18549_);
  or (_18553_, _18552_, _12380_);
  or (_18554_, _10458_, _08101_);
  or (_18555_, _10474_, _09208_);
  and (_18556_, _17011_, _08101_);
  or (_18557_, _06653_, \oc8051_golden_model_1.ACC [5]);
  nand (_18558_, _06653_, \oc8051_golden_model_1.ACC [5]);
  and (_18559_, _18558_, _18557_);
  and (_18560_, _18559_, _10471_);
  or (_18561_, _18560_, _10473_);
  or (_18563_, _18561_, _18556_);
  and (_18564_, _18563_, _10484_);
  and (_18565_, _18564_, _18555_);
  and (_18566_, _15119_, _07809_);
  or (_18567_, _18566_, _18512_);
  and (_18568_, _18567_, _06160_);
  or (_18569_, _18568_, _10490_);
  or (_18570_, _18569_, _18565_);
  nor (_18571_, _13858_, _10502_);
  nand (_18572_, _13858_, _10502_);
  nand (_18574_, _18572_, _10490_);
  or (_18575_, _18574_, _18571_);
  and (_18576_, _18575_, _06221_);
  and (_18577_, _18576_, _18570_);
  nor (_18578_, _08409_, _09930_);
  and (_18579_, _15123_, _08409_);
  or (_18580_, _18579_, _18578_);
  and (_18581_, _18580_, _06156_);
  and (_18582_, _18522_, _06217_);
  or (_18583_, _18582_, _10516_);
  or (_18585_, _18583_, _18581_);
  or (_18586_, _18585_, _18577_);
  and (_18587_, _18586_, _18554_);
  or (_18588_, _18587_, _07081_);
  or (_18589_, _09208_, _07082_);
  and (_18590_, _18589_, _06229_);
  and (_18591_, _18590_, _18588_);
  nor (_18592_, _08103_, _06229_);
  or (_18593_, _18592_, _10525_);
  or (_18594_, _18593_, _18591_);
  nand (_18596_, _10525_, _05887_);
  and (_18597_, _18596_, _18594_);
  or (_18598_, _18597_, _06152_);
  and (_18599_, _15104_, _08409_);
  or (_18600_, _18599_, _18578_);
  or (_18601_, _18600_, _06153_);
  and (_18602_, _18601_, _06146_);
  and (_18603_, _18602_, _18598_);
  or (_18604_, _18578_, _15138_);
  and (_18605_, _18580_, _06145_);
  and (_18607_, _18605_, _18604_);
  or (_18608_, _18607_, _18603_);
  and (_18609_, _18608_, _09301_);
  or (_18610_, _09783_, _09781_);
  nor (_18611_, _09784_, _09301_);
  and (_18612_, _18611_, _18610_);
  nor (_18613_, _06129_, _05803_);
  or (_18614_, _18613_, _10547_);
  or (_18615_, _18614_, _18612_);
  or (_18616_, _18615_, _18609_);
  and (_18618_, _06119_, _05790_);
  not (_18619_, _18618_);
  and (_18620_, _08349_, \oc8051_golden_model_1.ACC [4]);
  nor (_18621_, _18211_, _18620_);
  nor (_18622_, _18515_, _18621_);
  and (_18623_, _18515_, _18621_);
  nor (_18624_, _18623_, _18622_);
  and (_18625_, _18624_, \oc8051_golden_model_1.PSW [7]);
  nor (_18626_, _18624_, \oc8051_golden_model_1.PSW [7]);
  nor (_18627_, _18626_, _18625_);
  nor (_18629_, _18218_, _18215_);
  not (_18630_, _18629_);
  and (_18631_, _18630_, _18627_);
  nor (_18632_, _18630_, _18627_);
  nor (_18633_, _18632_, _18631_);
  and (_18634_, _18633_, _18619_);
  or (_18635_, _18634_, _10554_);
  and (_18636_, _18635_, _18616_);
  and (_18637_, _18633_, _18618_);
  or (_18638_, _18637_, _12379_);
  or (_18640_, _18638_, _18636_);
  and (_18641_, _18640_, _06265_);
  and (_18642_, _18641_, _18553_);
  and (_18643_, _08338_, \oc8051_golden_model_1.ACC [4]);
  nor (_18644_, _18292_, _18643_);
  nor (_18645_, _18644_, _12325_);
  and (_18646_, _18644_, _12325_);
  nor (_18647_, _18646_, _18645_);
  and (_18648_, _18647_, \oc8051_golden_model_1.PSW [7]);
  nor (_18649_, _18647_, \oc8051_golden_model_1.PSW [7]);
  nor (_18651_, _18649_, _18648_);
  nor (_18652_, _18299_, _18295_);
  not (_18653_, _18652_);
  or (_18654_, _18653_, _18651_);
  and (_18655_, _18653_, _18651_);
  nor (_18656_, _18655_, _06265_);
  and (_18657_, _18656_, _18654_);
  or (_18658_, _18657_, _10387_);
  or (_18659_, _18658_, _18642_);
  and (_18660_, _18659_, _18538_);
  or (_18661_, _18660_, _05870_);
  nand (_18662_, _06477_, _05870_);
  and (_18663_, _18662_, _06140_);
  and (_18664_, _18663_, _18661_);
  and (_18665_, _15155_, _08409_);
  or (_18666_, _18665_, _18578_);
  and (_18667_, _18666_, _06139_);
  or (_18668_, _18667_, _09842_);
  or (_18669_, _18668_, _18664_);
  and (_18670_, _18669_, _18523_);
  or (_18673_, _18670_, _06116_);
  and (_18674_, _09208_, _07809_);
  or (_18675_, _18512_, _06117_);
  or (_18676_, _18675_, _18674_);
  and (_18677_, _18676_, _06114_);
  and (_18678_, _18677_, _18673_);
  and (_18679_, _15203_, _07809_);
  or (_18680_, _18679_, _18512_);
  and (_18681_, _18680_, _05787_);
  or (_18682_, _18681_, _09855_);
  or (_18684_, _18682_, _18678_);
  or (_18685_, _09916_, _09861_);
  and (_18686_, _18685_, _05802_);
  and (_18687_, _18686_, _18684_);
  nor (_18688_, _06477_, _05802_);
  or (_18689_, _18688_, _06110_);
  or (_18690_, _18689_, _18687_);
  and (_18691_, _08736_, _07809_);
  or (_18692_, _18691_, _18512_);
  or (_18693_, _18692_, _06111_);
  and (_18694_, _18693_, _10752_);
  and (_18695_, _18694_, _18690_);
  or (_18696_, _18695_, _18520_);
  and (_18697_, _18696_, _10762_);
  and (_18698_, _18515_, _06558_);
  or (_18699_, _18698_, _06574_);
  or (_18700_, _18699_, _18697_);
  not (_18701_, _06574_);
  or (_18702_, _18515_, _18701_);
  and (_18703_, _18702_, _18516_);
  and (_18706_, _18703_, _18700_);
  or (_18707_, _18706_, _18519_);
  and (_18708_, _18707_, _10776_);
  nor (_18709_, _10776_, _11011_);
  or (_18710_, _18709_, _06400_);
  or (_18711_, _18710_, _18708_);
  or (_18712_, _12325_, _06401_);
  and (_18713_, _18712_, _10788_);
  and (_18714_, _18713_, _18711_);
  and (_18715_, _10787_, _12342_);
  or (_18717_, _18715_, _06297_);
  or (_18718_, _18717_, _18714_);
  and (_18719_, _18718_, _18514_);
  or (_18720_, _18719_, _06402_);
  and (_18721_, _06957_, _06408_);
  not (_18722_, _18721_);
  and (_18723_, _06684_, _06408_);
  and (_18724_, _06288_, _06408_);
  nor (_18725_, _18724_, _18723_);
  and (_18726_, _18725_, _18722_);
  and (_18727_, _18726_, _17408_);
  or (_18728_, _18512_, _07125_);
  and (_18729_, _18728_, _18727_);
  and (_18730_, _18729_, _18720_);
  and (_18731_, _06273_, _06408_);
  or (_18732_, _10970_, _18731_);
  and (_18733_, _18732_, _10812_);
  or (_18734_, _18733_, _18730_);
  not (_18735_, _18731_);
  or (_18736_, _10970_, _18735_);
  and (_18739_, _18736_, _18734_);
  or (_18740_, _18739_, _10811_);
  or (_18741_, _10816_, _11009_);
  and (_18742_, _18741_, _06410_);
  and (_18743_, _18742_, _18740_);
  or (_18744_, _10820_, _10268_);
  and (_18745_, _18744_, _10822_);
  or (_18746_, _18745_, _18743_);
  or (_18747_, _10826_, _11053_);
  and (_18748_, _18747_, _07132_);
  and (_18750_, _18748_, _18746_);
  nand (_18751_, _18692_, _06306_);
  nor (_18752_, _18751_, _10269_);
  or (_18753_, _18752_, _06524_);
  or (_18754_, _18753_, _18750_);
  nand (_18755_, _10971_, _06524_);
  and (_18756_, _18755_, _17150_);
  and (_18757_, _18756_, _18754_);
  nor (_18758_, _17150_, _10971_);
  or (_18759_, _18758_, _17156_);
  or (_18760_, _18759_, _18757_);
  nand (_18761_, _17156_, _10971_);
  and (_18762_, _18761_, _17161_);
  and (_18763_, _18762_, _18760_);
  nor (_18764_, _10971_, _17161_);
  or (_18765_, _18764_, _10841_);
  or (_18766_, _18765_, _18763_);
  nand (_18767_, _10841_, _09930_);
  or (_18768_, _18767_, _09208_);
  and (_18769_, _18768_, _06395_);
  and (_18772_, _18769_, _18766_);
  nand (_18773_, _10851_, _10269_);
  and (_18774_, _18773_, _10850_);
  or (_18775_, _18774_, _18772_);
  nand (_18776_, _10848_, _11054_);
  and (_18777_, _18776_, _08819_);
  and (_18778_, _18777_, _18775_);
  and (_18779_, _15216_, _07809_);
  or (_18780_, _18779_, _18512_);
  and (_18781_, _18780_, _06303_);
  or (_18783_, _18781_, _10858_);
  or (_18784_, _18783_, _18778_);
  and (_18785_, _18784_, _18510_);
  or (_18786_, _18785_, _10865_);
  and (_18787_, _10884_, _10599_);
  nor (_18788_, _18787_, _10885_);
  or (_18789_, _18788_, _10867_);
  and (_18790_, _18789_, _06407_);
  and (_18791_, _18790_, _18786_);
  and (_18792_, _10914_, _10410_);
  nor (_18793_, _18792_, _10915_);
  or (_18794_, _18793_, _10895_);
  and (_18795_, _18794_, _10897_);
  or (_18796_, _18795_, _18791_);
  and (_18797_, _10944_, _10676_);
  nor (_18798_, _18797_, _10945_);
  or (_18799_, _18798_, _10927_);
  and (_18800_, _18799_, _10926_);
  and (_18801_, _18800_, _18796_);
  nand (_18802_, _10925_, \oc8051_golden_model_1.ACC [4]);
  nand (_18805_, _18802_, _10963_);
  or (_18806_, _18805_, _18801_);
  and (_18807_, _10993_, _18515_);
  nor (_18808_, _10993_, _18515_);
  or (_18809_, _18808_, _18807_);
  or (_18810_, _18809_, _10963_);
  and (_18811_, _18810_, _18806_);
  or (_18812_, _18811_, _11003_);
  and (_18813_, _11035_, _11011_);
  nor (_18814_, _18813_, _11036_);
  or (_18816_, _18814_, _11041_);
  and (_18817_, _18816_, _06171_);
  and (_18818_, _18817_, _18812_);
  and (_18819_, _12325_, _10291_);
  nor (_18820_, _12325_, _10291_);
  or (_18821_, _18820_, _10264_);
  or (_18822_, _18821_, _18819_);
  and (_18823_, _18822_, _12691_);
  or (_18824_, _18823_, _18818_);
  and (_18825_, _11076_, _12342_);
  nor (_18826_, _11076_, _12342_);
  or (_18827_, _18826_, _10265_);
  or (_18828_, _18827_, _18825_);
  and (_18829_, _18828_, _12693_);
  and (_18830_, _18829_, _18824_);
  and (_18831_, _10262_, \oc8051_golden_model_1.ACC [4]);
  or (_18832_, _18831_, _06433_);
  or (_18833_, _18832_, _18830_);
  or (_18834_, _18567_, _06829_);
  and (_18835_, _18834_, _11090_);
  and (_18838_, _18835_, _18833_);
  nor (_18839_, _11097_, _09930_);
  or (_18840_, _18839_, _11098_);
  and (_18841_, _18840_, _11089_);
  or (_18842_, _18841_, _11094_);
  or (_18843_, _18842_, _18838_);
  nand (_18844_, _11094_, _09883_);
  and (_18845_, _18844_, _05749_);
  and (_18846_, _18845_, _18843_);
  and (_18847_, _18600_, _05748_);
  or (_18849_, _18847_, _06440_);
  or (_18850_, _18849_, _18846_);
  and (_18851_, _15275_, _07809_);
  or (_18852_, _18512_, _06444_);
  or (_18853_, _18852_, _18851_);
  and (_18854_, _18853_, _11113_);
  and (_18855_, _18854_, _18850_);
  nor (_18856_, _11123_, \oc8051_golden_model_1.ACC [5]);
  nor (_18857_, _18856_, _11124_);
  and (_18858_, _18857_, _11112_);
  or (_18859_, _18858_, _11119_);
  or (_18860_, _18859_, _18855_);
  nand (_18861_, _11119_, _09883_);
  and (_18862_, _18861_, _01317_);
  and (_18863_, _18862_, _18860_);
  or (_18864_, _18863_, _18506_);
  and (_43608_, _18864_, _43100_);
  nor (_18865_, _01317_, _09883_);
  nor (_18866_, _11037_, _11008_);
  nor (_18867_, _18866_, _11038_);
  or (_18870_, _18867_, _17201_);
  nor (_18871_, _10916_, _10448_);
  nor (_18872_, _18871_, _10917_);
  or (_18873_, _18872_, _06407_);
  and (_18874_, _18873_, _10927_);
  nand (_18875_, _10848_, _11051_);
  or (_18876_, _10967_, _18406_);
  and (_18877_, _15413_, _07809_);
  nor (_18878_, _07809_, _09883_);
  or (_18879_, _18878_, _07127_);
  or (_18881_, _18879_, _18877_);
  and (_18882_, _18178_, _10969_);
  and (_18883_, _15395_, _07809_);
  or (_18884_, _18883_, _18878_);
  and (_18885_, _18884_, _05787_);
  and (_18886_, _08012_, _07809_);
  or (_18887_, _18886_, _18878_);
  or (_18888_, _18887_, _06132_);
  or (_18889_, _09208_, _09930_);
  and (_18890_, _09208_, _09930_);
  or (_18892_, _18541_, _18890_);
  and (_18893_, _18892_, _18889_);
  nor (_18894_, _18893_, _11008_);
  and (_18895_, _18893_, _11008_);
  nor (_18896_, _18895_, _18894_);
  and (_18897_, _18549_, _18545_);
  nand (_18898_, _18897_, \oc8051_golden_model_1.PSW [7]);
  nor (_18899_, _18898_, _18896_);
  and (_18900_, _18898_, _18896_);
  or (_18901_, _18900_, _18899_);
  or (_18903_, _18901_, _12380_);
  or (_18904_, _10458_, _08012_);
  or (_18905_, _10474_, _09207_);
  and (_18906_, _17011_, _08012_);
  or (_18907_, _06653_, \oc8051_golden_model_1.ACC [6]);
  nand (_18908_, _06653_, \oc8051_golden_model_1.ACC [6]);
  and (_18909_, _18908_, _18907_);
  and (_18910_, _18909_, _10471_);
  or (_18911_, _18910_, _10473_);
  or (_18912_, _18911_, _18906_);
  and (_18914_, _18912_, _10484_);
  and (_18915_, _18914_, _18905_);
  and (_18916_, _15300_, _07809_);
  or (_18917_, _18916_, _18878_);
  and (_18918_, _18917_, _06160_);
  or (_18919_, _18918_, _10490_);
  or (_18920_, _18919_, _18915_);
  not (_18921_, _10504_);
  nor (_18922_, _18571_, _18921_);
  nand (_18923_, _10508_, _10505_);
  nand (_18925_, _18923_, _10490_);
  or (_18926_, _18925_, _18922_);
  and (_18927_, _18926_, _06221_);
  and (_18928_, _18927_, _18920_);
  nor (_18929_, _08409_, _09883_);
  and (_18930_, _15316_, _08409_);
  or (_18931_, _18930_, _18929_);
  and (_18932_, _18931_, _06156_);
  and (_18933_, _18887_, _06217_);
  or (_18934_, _18933_, _10516_);
  or (_18936_, _18934_, _18932_);
  or (_18937_, _18936_, _18928_);
  and (_18938_, _18937_, _18904_);
  or (_18939_, _18938_, _07081_);
  or (_18940_, _09207_, _07082_);
  and (_18941_, _18940_, _06229_);
  and (_18942_, _18941_, _18939_);
  nor (_18943_, _08014_, _06229_);
  or (_18944_, _18943_, _10525_);
  or (_18945_, _18944_, _18942_);
  nand (_18947_, _10525_, _09981_);
  and (_18948_, _18947_, _18945_);
  or (_18949_, _18948_, _06152_);
  and (_18950_, _15297_, _08409_);
  or (_18951_, _18950_, _18929_);
  or (_18952_, _18951_, _06153_);
  and (_18953_, _18952_, _06146_);
  and (_18954_, _18953_, _18949_);
  or (_18955_, _18929_, _15331_);
  and (_18956_, _18931_, _06145_);
  and (_18958_, _18956_, _18955_);
  or (_18959_, _18958_, _09295_);
  or (_18960_, _18959_, _18954_);
  nor (_18961_, _09786_, _09784_);
  nor (_18962_, _18961_, _09787_);
  or (_18963_, _18962_, _09301_);
  and (_18964_, _18963_, _10554_);
  and (_18965_, _18964_, _18960_);
  or (_18966_, _08101_, _09930_);
  and (_18967_, _08101_, _09930_);
  or (_18969_, _18621_, _18967_);
  and (_18970_, _18969_, _18966_);
  nor (_18971_, _18970_, _10969_);
  and (_18972_, _18970_, _10969_);
  nor (_18973_, _18972_, _18971_);
  nor (_18974_, _18631_, _18625_);
  and (_18975_, _18974_, \oc8051_golden_model_1.PSW [7]);
  or (_18976_, _18975_, _18973_);
  nand (_18977_, _18975_, _18973_);
  and (_18978_, _18977_, _18976_);
  nand (_18980_, _18978_, _10557_);
  nand (_18981_, _18980_, _12380_);
  or (_18982_, _18981_, _18965_);
  and (_18983_, _18982_, _06265_);
  and (_18984_, _18983_, _18903_);
  nor (_18985_, _18655_, _18648_);
  or (_18986_, _18644_, _13929_);
  and (_18987_, _18986_, _13927_);
  nor (_18988_, _18987_, _10295_);
  and (_18989_, _18987_, _10295_);
  nor (_18991_, _18989_, _18988_);
  nor (_18992_, _18991_, _10693_);
  and (_18993_, _18991_, _10693_);
  nor (_18994_, _18993_, _18992_);
  nand (_18995_, _18994_, _18985_);
  or (_18996_, _18994_, _18985_);
  and (_18997_, _18996_, _06260_);
  and (_18998_, _18997_, _18995_);
  or (_18999_, _18998_, _18984_);
  and (_19000_, _18999_, _10388_);
  or (_19002_, _18525_, _13957_);
  and (_19003_, _19002_, _13956_);
  nor (_19004_, _19003_, _11052_);
  and (_19005_, _19003_, _11052_);
  nor (_19006_, _19005_, _19004_);
  nor (_19007_, _18535_, _18530_);
  and (_19008_, _19007_, \oc8051_golden_model_1.PSW [7]);
  or (_19009_, _19008_, _19006_);
  nand (_19010_, _19008_, _19006_);
  and (_19011_, _19010_, _10387_);
  and (_19013_, _19011_, _19009_);
  or (_19014_, _19013_, _05870_);
  or (_19015_, _19014_, _19000_);
  nand (_19016_, _06203_, _05870_);
  and (_19017_, _19016_, _06140_);
  and (_19018_, _19017_, _19015_);
  and (_19019_, _15348_, _08409_);
  or (_19020_, _19019_, _18929_);
  and (_19021_, _19020_, _06139_);
  or (_19022_, _19021_, _09842_);
  or (_19024_, _19022_, _19018_);
  and (_19025_, _19024_, _18888_);
  or (_19026_, _19025_, _06116_);
  and (_19027_, _09207_, _07809_);
  or (_19028_, _18878_, _06117_);
  or (_19029_, _19028_, _19027_);
  and (_19030_, _19029_, _06114_);
  and (_19031_, _19030_, _19026_);
  or (_19032_, _19031_, _18885_);
  and (_19033_, _19032_, _11922_);
  nor (_19035_, _06203_, _05802_);
  not (_19036_, _09888_);
  nor (_19037_, _19036_, _09884_);
  and (_19038_, _19037_, _05799_);
  and (_19039_, _19038_, _09855_);
  or (_19040_, _19039_, _19035_);
  or (_19041_, _19040_, _19033_);
  and (_19042_, _19041_, _06111_);
  and (_19043_, _15402_, _07809_);
  or (_19044_, _19043_, _18878_);
  and (_19046_, _19044_, _06110_);
  or (_19047_, _19046_, _10751_);
  or (_19048_, _19047_, _19042_);
  nand (_19049_, _10751_, _06203_);
  and (_19050_, _19049_, _18182_);
  and (_19051_, _19050_, _19048_);
  and (_19052_, _10969_, _18181_);
  nor (_19053_, _19052_, _19051_);
  or (_19054_, _19053_, _18174_);
  nand (_19055_, _10969_, _18174_);
  and (_19057_, _19055_, _19054_);
  nor (_19058_, _19057_, _18175_);
  and (_19059_, _10969_, _18175_);
  or (_19060_, _19059_, _06574_);
  or (_19061_, _19060_, _19058_);
  nor (_19062_, _10969_, _18701_);
  or (_19063_, _19062_, _17709_);
  nor (_19064_, _19063_, _17714_);
  and (_19065_, _19064_, _19061_);
  or (_19066_, _19065_, _18882_);
  and (_19068_, _19066_, _18172_);
  and (_19069_, _17105_, _10969_);
  or (_19070_, _19069_, _06771_);
  or (_19071_, _19070_, _19068_);
  or (_19072_, _10969_, _17113_);
  and (_19073_, _19072_, _10776_);
  and (_19074_, _19073_, _19071_);
  and (_19075_, _10775_, _11008_);
  or (_19076_, _19075_, _06400_);
  or (_19077_, _19076_, _19074_);
  or (_19079_, _10295_, _06401_);
  and (_19080_, _19079_, _10788_);
  and (_19081_, _19080_, _19077_);
  and (_19082_, _10787_, _11052_);
  or (_19083_, _19082_, _06297_);
  or (_19084_, _19083_, _19081_);
  and (_19085_, _19084_, _18881_);
  or (_19086_, _19085_, _06402_);
  or (_19087_, _18878_, _07125_);
  and (_19088_, _19087_, _10808_);
  and (_19090_, _19088_, _19086_);
  and (_19091_, _10812_, _10966_);
  or (_19092_, _19091_, _10811_);
  or (_19093_, _19092_, _19090_);
  or (_19094_, _10816_, _11005_);
  and (_19095_, _19094_, _06410_);
  and (_19096_, _19095_, _19093_);
  and (_19097_, _10266_, _06409_);
  or (_19098_, _19097_, _10820_);
  or (_19099_, _19098_, _19096_);
  or (_19101_, _10826_, _11049_);
  and (_19102_, _19101_, _07132_);
  and (_19103_, _19102_, _19099_);
  nand (_19104_, _19044_, _06306_);
  nor (_19105_, _19104_, _10294_);
  or (_19106_, _19105_, _06524_);
  or (_19107_, _19106_, _19103_);
  and (_19108_, _19107_, _18876_);
  or (_19109_, _19108_, _06555_);
  nor (_19110_, _10967_, _10834_);
  nor (_19112_, _19110_, _06975_);
  and (_19113_, _19112_, _19109_);
  and (_19114_, _10967_, _06975_);
  or (_19115_, _19114_, _19113_);
  and (_19116_, _19115_, _17847_);
  and (_19117_, _10835_, _10967_);
  or (_19118_, _19117_, _10841_);
  or (_19119_, _19118_, _19116_);
  or (_19120_, _17242_, _11006_);
  and (_19121_, _19120_, _06395_);
  and (_19123_, _19121_, _19119_);
  nand (_19124_, _10851_, _10294_);
  and (_19125_, _19124_, _10850_);
  or (_19126_, _19125_, _19123_);
  and (_19127_, _19126_, _18875_);
  or (_19128_, _19127_, _06303_);
  and (_19129_, _15410_, _07809_);
  or (_19130_, _18878_, _08819_);
  or (_19131_, _19130_, _19129_);
  and (_19132_, _19131_, _10380_);
  and (_19134_, _19132_, _19128_);
  or (_19135_, _10365_, _10316_);
  and (_19136_, _10858_, _10366_);
  and (_19137_, _19136_, _19135_);
  or (_19138_, _19137_, _19134_);
  or (_19139_, _19138_, _17240_);
  or (_19140_, _10886_, _10641_);
  and (_19141_, _19140_, _10887_);
  and (_19142_, _19141_, _06276_);
  or (_19143_, _19142_, _10867_);
  and (_19145_, _19143_, _19139_);
  and (_19146_, _19141_, _06792_);
  or (_19147_, _19146_, _06406_);
  or (_19148_, _19147_, _19145_);
  and (_19149_, _19148_, _18874_);
  or (_19150_, _10946_, _10714_);
  nor (_19151_, _10947_, _10927_);
  and (_19152_, _19151_, _19150_);
  or (_19153_, _19152_, _10925_);
  or (_19154_, _19153_, _19149_);
  nand (_19156_, _10925_, _09930_);
  and (_19157_, _19156_, _10963_);
  and (_19158_, _19157_, _19154_);
  nor (_19159_, _10995_, _10969_);
  nor (_19160_, _19159_, _10996_);
  and (_19161_, _19160_, _18454_);
  or (_19162_, _19161_, _17195_);
  or (_19163_, _19162_, _19158_);
  and (_19164_, _19163_, _18870_);
  or (_19165_, _19164_, _17199_);
  or (_19167_, _18867_, _17200_);
  and (_19168_, _19167_, _06171_);
  and (_19169_, _19168_, _19165_);
  or (_19170_, _10295_, _10293_);
  and (_19171_, _19170_, _10296_);
  or (_19172_, _19171_, _10264_);
  and (_19173_, _19172_, _12691_);
  or (_19174_, _19173_, _19169_);
  or (_19175_, _11078_, _11052_);
  and (_19176_, _19175_, _11079_);
  or (_19178_, _19176_, _10265_);
  and (_19179_, _19178_, _12693_);
  and (_19180_, _19179_, _19174_);
  and (_19181_, _10262_, \oc8051_golden_model_1.ACC [5]);
  or (_19182_, _19181_, _06433_);
  or (_19183_, _19182_, _19180_);
  or (_19184_, _18917_, _06829_);
  and (_19185_, _19184_, _11090_);
  and (_19186_, _19185_, _19183_);
  nor (_19187_, _11098_, _09883_);
  or (_19189_, _19187_, _11099_);
  and (_19190_, _19189_, _11089_);
  or (_19191_, _19190_, _11094_);
  or (_19192_, _19191_, _19186_);
  nand (_19193_, _11094_, _08430_);
  and (_19194_, _19193_, _05749_);
  and (_19195_, _19194_, _19192_);
  and (_19196_, _18951_, _05748_);
  or (_19197_, _19196_, _06440_);
  or (_19198_, _19197_, _19195_);
  and (_19200_, _15478_, _07809_);
  or (_19201_, _18878_, _06444_);
  or (_19202_, _19201_, _19200_);
  and (_19203_, _19202_, _11113_);
  and (_19204_, _19203_, _19198_);
  nor (_19205_, _11124_, \oc8051_golden_model_1.ACC [6]);
  nor (_19206_, _19205_, _11125_);
  and (_19207_, _19206_, _11112_);
  or (_19208_, _19207_, _11119_);
  or (_19209_, _19208_, _19204_);
  nand (_19211_, _11119_, _08430_);
  and (_19212_, _19211_, _01317_);
  and (_19213_, _19212_, _19209_);
  or (_19214_, _19213_, _18865_);
  and (_43609_, _19214_, _43100_);
  not (_19215_, \oc8051_golden_model_1.PCON [0]);
  nor (_19216_, _01317_, _19215_);
  and (_19217_, _07856_, \oc8051_golden_model_1.ACC [0]);
  and (_19218_, _19217_, _08211_);
  nor (_19219_, _07856_, _19215_);
  or (_19221_, _19219_, _07130_);
  or (_19222_, _19221_, _19218_);
  nor (_19223_, _08211_, _11137_);
  or (_19224_, _19223_, _19219_);
  or (_19225_, _19224_, _06161_);
  or (_19226_, _19219_, _19217_);
  and (_19227_, _19226_, _07056_);
  nor (_19228_, _07056_, _19215_);
  or (_19229_, _19228_, _06160_);
  or (_19230_, _19229_, _19227_);
  and (_19232_, _19230_, _07075_);
  and (_19233_, _19232_, _19225_);
  and (_19234_, _07856_, _07049_);
  or (_19235_, _19234_, _19219_);
  and (_19236_, _19235_, _06217_);
  or (_19237_, _19236_, _19233_);
  and (_19238_, _19237_, _06229_);
  and (_19239_, _19226_, _06220_);
  or (_19240_, _19239_, _09842_);
  or (_19241_, _19240_, _19238_);
  or (_19243_, _19235_, _06132_);
  and (_19244_, _19243_, _19241_);
  or (_19245_, _19244_, _06116_);
  and (_19246_, _09160_, _07856_);
  or (_19247_, _19219_, _06117_);
  or (_19248_, _19247_, _19246_);
  and (_19249_, _19248_, _19245_);
  or (_19250_, _19249_, _05787_);
  and (_19251_, _14260_, _07856_);
  or (_19252_, _19219_, _06114_);
  or (_19254_, _19252_, _19251_);
  and (_19255_, _19254_, _06111_);
  and (_19256_, _19255_, _19250_);
  and (_19257_, _07856_, _08708_);
  or (_19258_, _19257_, _19219_);
  and (_19259_, _19258_, _06110_);
  or (_19260_, _19259_, _06297_);
  or (_19261_, _19260_, _19256_);
  and (_19262_, _14275_, _07856_);
  or (_19263_, _19262_, _19219_);
  or (_19265_, _19263_, _07127_);
  and (_19266_, _19265_, _07125_);
  and (_19267_, _19266_, _19261_);
  nor (_19268_, _12321_, _11137_);
  or (_19269_, _19268_, _19219_);
  nor (_19270_, _19218_, _07125_);
  and (_19271_, _19270_, _19269_);
  or (_19272_, _19271_, _19267_);
  and (_19273_, _19272_, _07132_);
  nand (_19274_, _19258_, _06306_);
  nor (_19276_, _19274_, _19223_);
  or (_19277_, _19276_, _06411_);
  or (_19278_, _19277_, _19273_);
  and (_19279_, _19278_, _19222_);
  or (_19280_, _19279_, _06303_);
  and (_19281_, _14167_, _07856_);
  or (_19282_, _19219_, _08819_);
  or (_19283_, _19282_, _19281_);
  and (_19284_, _19283_, _08824_);
  and (_19285_, _19284_, _19280_);
  not (_19287_, _06630_);
  and (_19288_, _19269_, _06396_);
  or (_19289_, _19288_, _19287_);
  or (_19290_, _19289_, _19285_);
  or (_19291_, _19224_, _06630_);
  and (_19292_, _19291_, _01317_);
  and (_19293_, _19292_, _19290_);
  or (_19294_, _19293_, _19216_);
  and (_43611_, _19294_, _43100_);
  not (_19295_, \oc8051_golden_model_1.PCON [1]);
  nor (_19297_, _01317_, _19295_);
  or (_19298_, _14442_, _11137_);
  or (_19299_, _07856_, \oc8051_golden_model_1.PCON [1]);
  and (_19300_, _19299_, _05787_);
  and (_19301_, _19300_, _19298_);
  and (_19302_, _09115_, _07856_);
  nor (_19303_, _07856_, _19295_);
  or (_19304_, _19303_, _06117_);
  or (_19305_, _19304_, _19302_);
  and (_19306_, _07856_, _07306_);
  or (_19308_, _19306_, _19303_);
  or (_19309_, _19308_, _06132_);
  and (_19310_, _14363_, _07856_);
  not (_19311_, _19310_);
  and (_19312_, _19311_, _19299_);
  or (_19313_, _19312_, _06161_);
  and (_19314_, _07856_, \oc8051_golden_model_1.ACC [1]);
  or (_19315_, _19314_, _19303_);
  and (_19316_, _19315_, _07056_);
  nor (_19317_, _07056_, _19295_);
  or (_19319_, _19317_, _06160_);
  or (_19320_, _19319_, _19316_);
  and (_19321_, _19320_, _07075_);
  and (_19322_, _19321_, _19313_);
  and (_19323_, _19308_, _06217_);
  or (_19324_, _19323_, _19322_);
  and (_19325_, _19324_, _06229_);
  and (_19326_, _19315_, _06220_);
  or (_19327_, _19326_, _09842_);
  or (_19328_, _19327_, _19325_);
  and (_19330_, _19328_, _19309_);
  or (_19331_, _19330_, _06116_);
  and (_19332_, _19331_, _06114_);
  and (_19333_, _19332_, _19305_);
  or (_19334_, _19333_, _19301_);
  and (_19335_, _19334_, _06298_);
  or (_19336_, _14346_, _11137_);
  and (_19337_, _19299_, _06297_);
  and (_19338_, _19337_, _19336_);
  nand (_19339_, _07856_, _06945_);
  and (_19341_, _19299_, _06110_);
  and (_19342_, _19341_, _19339_);
  or (_19343_, _19342_, _06402_);
  or (_19344_, _19343_, _19338_);
  or (_19345_, _19344_, _19335_);
  and (_19346_, _10278_, _07856_);
  or (_19347_, _19346_, _19303_);
  or (_19348_, _19347_, _07125_);
  and (_19349_, _19348_, _07132_);
  and (_19350_, _19349_, _19345_);
  or (_19352_, _14344_, _11137_);
  and (_19353_, _19299_, _06306_);
  and (_19354_, _19353_, _19352_);
  or (_19355_, _19354_, _06411_);
  or (_19356_, _19355_, _19350_);
  and (_19357_, _19314_, _08176_);
  or (_19358_, _19303_, _07130_);
  or (_19359_, _19358_, _19357_);
  and (_19360_, _19359_, _08819_);
  and (_19361_, _19360_, _19356_);
  or (_19363_, _19339_, _08176_);
  and (_19364_, _19299_, _06303_);
  and (_19365_, _19364_, _19363_);
  or (_19366_, _19365_, _06396_);
  or (_19367_, _19366_, _19361_);
  nor (_19368_, _10277_, _11137_);
  or (_19369_, _19368_, _19303_);
  or (_19370_, _19369_, _08824_);
  and (_19371_, _19370_, _19367_);
  and (_19372_, _19371_, _06829_);
  and (_19374_, _19312_, _06433_);
  or (_19375_, _19374_, _06440_);
  or (_19376_, _19375_, _19372_);
  or (_19377_, _19303_, _06444_);
  or (_19378_, _19377_, _19310_);
  and (_19379_, _19378_, _01317_);
  and (_19380_, _19379_, _19376_);
  or (_19381_, _19380_, _19297_);
  and (_43612_, _19381_, _43100_);
  not (_19382_, \oc8051_golden_model_1.PCON [2]);
  nor (_19384_, _01317_, _19382_);
  nor (_19385_, _07856_, _19382_);
  and (_19386_, _07856_, _07708_);
  or (_19387_, _19386_, _19385_);
  or (_19388_, _19387_, _06132_);
  and (_19389_, _14542_, _07856_);
  or (_19390_, _19389_, _19385_);
  and (_19391_, _19390_, _06160_);
  nor (_19392_, _07056_, _19382_);
  and (_19393_, _07856_, \oc8051_golden_model_1.ACC [2]);
  or (_19395_, _19393_, _19385_);
  and (_19396_, _19395_, _07056_);
  or (_19397_, _19396_, _19392_);
  and (_19398_, _19397_, _06161_);
  or (_19399_, _19398_, _06217_);
  or (_19400_, _19399_, _19391_);
  or (_19401_, _19387_, _07075_);
  and (_19402_, _19401_, _06229_);
  and (_19403_, _19402_, _19400_);
  and (_19404_, _19395_, _06220_);
  or (_19406_, _19404_, _09842_);
  or (_19407_, _19406_, _19403_);
  and (_19408_, _19407_, _19388_);
  or (_19409_, _19408_, _06116_);
  and (_19410_, _09211_, _07856_);
  or (_19411_, _19385_, _06117_);
  or (_19412_, _19411_, _19410_);
  and (_19413_, _19412_, _19409_);
  or (_19414_, _19413_, _05787_);
  and (_19415_, _14630_, _07856_);
  or (_19417_, _19415_, _19385_);
  or (_19418_, _19417_, _06114_);
  and (_19419_, _19418_, _06111_);
  and (_19420_, _19419_, _19414_);
  and (_19421_, _07856_, _08768_);
  or (_19422_, _19421_, _19385_);
  and (_19423_, _19422_, _06110_);
  or (_19424_, _19423_, _06297_);
  or (_19425_, _19424_, _19420_);
  and (_19426_, _14646_, _07856_);
  or (_19428_, _19385_, _07127_);
  or (_19429_, _19428_, _19426_);
  and (_19430_, _19429_, _07125_);
  and (_19431_, _19430_, _19425_);
  and (_19432_, _10282_, _07856_);
  or (_19433_, _19432_, _19385_);
  and (_19434_, _19433_, _06402_);
  or (_19435_, _19434_, _19431_);
  and (_19436_, _19435_, _07132_);
  or (_19437_, _19385_, _08248_);
  and (_19439_, _19422_, _06306_);
  and (_19440_, _19439_, _19437_);
  or (_19441_, _19440_, _19436_);
  and (_19442_, _19441_, _07130_);
  and (_19443_, _19395_, _06411_);
  and (_19444_, _19443_, _19437_);
  or (_19445_, _19444_, _06303_);
  or (_19446_, _19445_, _19442_);
  and (_19447_, _14643_, _07856_);
  or (_19448_, _19385_, _08819_);
  or (_19450_, _19448_, _19447_);
  and (_19451_, _19450_, _08824_);
  and (_19452_, _19451_, _19446_);
  nor (_19453_, _10281_, _11137_);
  or (_19454_, _19453_, _19385_);
  and (_19455_, _19454_, _06396_);
  or (_19456_, _19455_, _19452_);
  and (_19457_, _19456_, _06829_);
  and (_19458_, _19390_, _06433_);
  or (_19459_, _19458_, _06440_);
  or (_19461_, _19459_, _19457_);
  and (_19462_, _14710_, _07856_);
  or (_19463_, _19385_, _06444_);
  or (_19464_, _19463_, _19462_);
  and (_19465_, _19464_, _01317_);
  and (_19466_, _19465_, _19461_);
  or (_19467_, _19466_, _19384_);
  and (_43613_, _19467_, _43100_);
  and (_19468_, _11137_, \oc8051_golden_model_1.PCON [3]);
  and (_19469_, _14738_, _07856_);
  or (_19471_, _19469_, _19468_);
  or (_19472_, _19471_, _06161_);
  and (_19473_, _07856_, \oc8051_golden_model_1.ACC [3]);
  or (_19474_, _19473_, _19468_);
  and (_19475_, _19474_, _07056_);
  and (_19476_, _07057_, \oc8051_golden_model_1.PCON [3]);
  or (_19477_, _19476_, _06160_);
  or (_19478_, _19477_, _19475_);
  and (_19479_, _19478_, _07075_);
  and (_19480_, _19479_, _19472_);
  and (_19482_, _07856_, _07544_);
  or (_19483_, _19482_, _19468_);
  and (_19484_, _19483_, _06217_);
  or (_19485_, _19484_, _19480_);
  and (_19486_, _19485_, _06229_);
  and (_19487_, _19474_, _06220_);
  or (_19488_, _19487_, _09842_);
  or (_19489_, _19488_, _19486_);
  or (_19490_, _19483_, _06132_);
  and (_19491_, _19490_, _06117_);
  and (_19493_, _19491_, _19489_);
  and (_19494_, _09210_, _07856_);
  or (_19495_, _19494_, _19468_);
  and (_19496_, _19495_, _06116_);
  or (_19497_, _19496_, _05787_);
  or (_19498_, _19497_, _19493_);
  and (_19499_, _14825_, _07856_);
  or (_19500_, _19499_, _19468_);
  or (_19501_, _19500_, _06114_);
  and (_19502_, _19501_, _06111_);
  and (_19504_, _19502_, _19498_);
  and (_19505_, _07856_, _08712_);
  or (_19506_, _19505_, _19468_);
  and (_19507_, _19506_, _06110_);
  or (_19508_, _19507_, _06297_);
  or (_19509_, _19508_, _19504_);
  and (_19510_, _14727_, _07856_);
  or (_19511_, _19510_, _19468_);
  or (_19512_, _19511_, _07127_);
  and (_19513_, _19512_, _07125_);
  and (_19515_, _19513_, _19509_);
  and (_19516_, _12318_, _07856_);
  or (_19517_, _19516_, _19468_);
  and (_19518_, _19517_, _06402_);
  or (_19519_, _19518_, _19515_);
  and (_19520_, _19519_, _07132_);
  or (_19521_, _19468_, _08140_);
  and (_19522_, _19506_, _06306_);
  and (_19523_, _19522_, _19521_);
  or (_19524_, _19523_, _19520_);
  and (_19526_, _19524_, _07130_);
  and (_19527_, _19474_, _06411_);
  and (_19528_, _19527_, _19521_);
  or (_19529_, _19528_, _06303_);
  or (_19530_, _19529_, _19526_);
  and (_19531_, _14724_, _07856_);
  or (_19532_, _19468_, _08819_);
  or (_19533_, _19532_, _19531_);
  and (_19534_, _19533_, _08824_);
  and (_19535_, _19534_, _19530_);
  nor (_19537_, _10273_, _11137_);
  or (_19538_, _19537_, _19468_);
  and (_19539_, _19538_, _06396_);
  or (_19540_, _19539_, _06433_);
  or (_19541_, _19540_, _19535_);
  or (_19542_, _19471_, _06829_);
  and (_19543_, _19542_, _06444_);
  and (_19544_, _19543_, _19541_);
  and (_19545_, _14897_, _07856_);
  or (_19546_, _19545_, _19468_);
  and (_19548_, _19546_, _06440_);
  or (_19549_, _19548_, _01321_);
  or (_19550_, _19549_, _19544_);
  or (_19551_, _01317_, \oc8051_golden_model_1.PCON [3]);
  and (_19552_, _19551_, _43100_);
  and (_43614_, _19552_, _19550_);
  and (_19553_, _11137_, \oc8051_golden_model_1.PCON [4]);
  and (_19554_, _08336_, _07856_);
  or (_19555_, _19554_, _19553_);
  or (_19556_, _19555_, _06132_);
  and (_19558_, _14928_, _07856_);
  or (_19559_, _19558_, _19553_);
  or (_19560_, _19559_, _06161_);
  and (_19561_, _07856_, \oc8051_golden_model_1.ACC [4]);
  or (_19562_, _19561_, _19553_);
  and (_19563_, _19562_, _07056_);
  and (_19564_, _07057_, \oc8051_golden_model_1.PCON [4]);
  or (_19565_, _19564_, _06160_);
  or (_19566_, _19565_, _19563_);
  and (_19567_, _19566_, _07075_);
  and (_19569_, _19567_, _19560_);
  and (_19570_, _19555_, _06217_);
  or (_19571_, _19570_, _19569_);
  and (_19572_, _19571_, _06229_);
  and (_19573_, _19562_, _06220_);
  or (_19574_, _19573_, _09842_);
  or (_19575_, _19574_, _19572_);
  and (_19576_, _19575_, _19556_);
  or (_19577_, _19576_, _06116_);
  and (_19578_, _09209_, _07856_);
  or (_19580_, _19553_, _06117_);
  or (_19581_, _19580_, _19578_);
  and (_19582_, _19581_, _06114_);
  and (_19583_, _19582_, _19577_);
  and (_19584_, _15013_, _07856_);
  or (_19585_, _19584_, _19553_);
  and (_19586_, _19585_, _05787_);
  or (_19587_, _19586_, _19583_);
  or (_19588_, _19587_, _11136_);
  and (_19589_, _15029_, _07856_);
  or (_19591_, _19553_, _07127_);
  or (_19592_, _19591_, _19589_);
  and (_19593_, _08715_, _07856_);
  or (_19594_, _19593_, _19553_);
  or (_19595_, _19594_, _06111_);
  and (_19596_, _19595_, _07125_);
  and (_19597_, _19596_, _19592_);
  and (_19598_, _19597_, _19588_);
  and (_19599_, _10289_, _07856_);
  or (_19600_, _19599_, _19553_);
  and (_19602_, _19600_, _06402_);
  or (_19603_, _19602_, _19598_);
  and (_19604_, _19603_, _07132_);
  or (_19605_, _19553_, _08339_);
  and (_19606_, _19594_, _06306_);
  and (_19607_, _19606_, _19605_);
  or (_19608_, _19607_, _19604_);
  and (_19609_, _19608_, _07130_);
  and (_19610_, _19562_, _06411_);
  and (_19611_, _19610_, _19605_);
  or (_19613_, _19611_, _06303_);
  or (_19614_, _19613_, _19609_);
  and (_19615_, _15026_, _07856_);
  or (_19616_, _19553_, _08819_);
  or (_19617_, _19616_, _19615_);
  and (_19618_, _19617_, _08824_);
  and (_19619_, _19618_, _19614_);
  nor (_19620_, _10288_, _11137_);
  or (_19621_, _19620_, _19553_);
  and (_19622_, _19621_, _06396_);
  or (_19624_, _19622_, _06433_);
  or (_19625_, _19624_, _19619_);
  or (_19626_, _19559_, _06829_);
  and (_19627_, _19626_, _06444_);
  and (_19628_, _19627_, _19625_);
  and (_19629_, _15087_, _07856_);
  or (_19630_, _19629_, _19553_);
  and (_19631_, _19630_, _06440_);
  or (_19632_, _19631_, _01321_);
  or (_19633_, _19632_, _19628_);
  or (_19635_, _01317_, \oc8051_golden_model_1.PCON [4]);
  and (_19636_, _19635_, _43100_);
  and (_43615_, _19636_, _19633_);
  and (_19637_, _11137_, \oc8051_golden_model_1.PCON [5]);
  or (_19638_, _19637_, _08104_);
  and (_19639_, _08736_, _07856_);
  or (_19640_, _19639_, _19637_);
  and (_19641_, _19640_, _06306_);
  and (_19642_, _19641_, _19638_);
  and (_19643_, _15119_, _07856_);
  or (_19645_, _19643_, _19637_);
  or (_19646_, _19645_, _06161_);
  and (_19647_, _07856_, \oc8051_golden_model_1.ACC [5]);
  or (_19648_, _19647_, _19637_);
  and (_19649_, _19648_, _07056_);
  and (_19650_, _07057_, \oc8051_golden_model_1.PCON [5]);
  or (_19651_, _19650_, _06160_);
  or (_19652_, _19651_, _19649_);
  and (_19653_, _19652_, _07075_);
  and (_19654_, _19653_, _19646_);
  and (_19656_, _08101_, _07856_);
  or (_19657_, _19656_, _19637_);
  and (_19658_, _19657_, _06217_);
  or (_19659_, _19658_, _19654_);
  and (_19660_, _19659_, _06229_);
  and (_19661_, _19648_, _06220_);
  or (_19662_, _19661_, _09842_);
  or (_19663_, _19662_, _19660_);
  or (_19664_, _19657_, _06132_);
  and (_19665_, _19664_, _19663_);
  or (_19667_, _19665_, _06116_);
  and (_19668_, _09208_, _07856_);
  or (_19669_, _19637_, _06117_);
  or (_19670_, _19669_, _19668_);
  and (_19671_, _19670_, _06114_);
  and (_19672_, _19671_, _19667_);
  and (_19673_, _15203_, _07856_);
  or (_19674_, _19673_, _19637_);
  and (_19675_, _19674_, _05787_);
  or (_19676_, _19675_, _11136_);
  or (_19678_, _19676_, _19672_);
  and (_19679_, _15219_, _07856_);
  or (_19680_, _19637_, _07127_);
  or (_19681_, _19680_, _19679_);
  or (_19682_, _19640_, _06111_);
  and (_19683_, _19682_, _07125_);
  and (_19684_, _19683_, _19681_);
  and (_19685_, _19684_, _19678_);
  and (_19686_, _12325_, _07856_);
  or (_19687_, _19686_, _19637_);
  and (_19689_, _19687_, _06402_);
  or (_19690_, _19689_, _19685_);
  and (_19691_, _19690_, _07132_);
  or (_19692_, _19691_, _19642_);
  and (_19693_, _19692_, _07130_);
  and (_19694_, _19648_, _06411_);
  and (_19695_, _19694_, _19638_);
  or (_19696_, _19695_, _06303_);
  or (_19697_, _19696_, _19693_);
  and (_19698_, _15216_, _07856_);
  or (_19700_, _19637_, _08819_);
  or (_19701_, _19700_, _19698_);
  and (_19702_, _19701_, _08824_);
  and (_19703_, _19702_, _19697_);
  nor (_19704_, _10269_, _11137_);
  or (_19705_, _19704_, _19637_);
  and (_19706_, _19705_, _06396_);
  or (_19707_, _19706_, _06433_);
  or (_19708_, _19707_, _19703_);
  or (_19709_, _19645_, _06829_);
  and (_19711_, _19709_, _06444_);
  and (_19712_, _19711_, _19708_);
  and (_19713_, _15275_, _07856_);
  or (_19714_, _19713_, _19637_);
  and (_19715_, _19714_, _06440_);
  or (_19716_, _19715_, _01321_);
  or (_19717_, _19716_, _19712_);
  or (_19718_, _01317_, \oc8051_golden_model_1.PCON [5]);
  and (_19719_, _19718_, _43100_);
  and (_43617_, _19719_, _19717_);
  and (_19721_, _11137_, \oc8051_golden_model_1.PCON [6]);
  or (_19722_, _19721_, _08015_);
  and (_19723_, _15402_, _07856_);
  or (_19724_, _19723_, _19721_);
  and (_19725_, _19724_, _06306_);
  and (_19726_, _19725_, _19722_);
  and (_19727_, _15300_, _07856_);
  or (_19728_, _19727_, _19721_);
  or (_19729_, _19728_, _06161_);
  and (_19730_, _07856_, \oc8051_golden_model_1.ACC [6]);
  or (_19732_, _19730_, _19721_);
  and (_19733_, _19732_, _07056_);
  and (_19734_, _07057_, \oc8051_golden_model_1.PCON [6]);
  or (_19735_, _19734_, _06160_);
  or (_19736_, _19735_, _19733_);
  and (_19737_, _19736_, _07075_);
  and (_19738_, _19737_, _19729_);
  and (_19739_, _08012_, _07856_);
  or (_19740_, _19739_, _19721_);
  and (_19741_, _19740_, _06217_);
  or (_19743_, _19741_, _19738_);
  and (_19744_, _19743_, _06229_);
  and (_19745_, _19732_, _06220_);
  or (_19746_, _19745_, _09842_);
  or (_19747_, _19746_, _19744_);
  or (_19748_, _19740_, _06132_);
  and (_19749_, _19748_, _19747_);
  or (_19750_, _19749_, _06116_);
  and (_19751_, _09207_, _07856_);
  or (_19752_, _19721_, _06117_);
  or (_19754_, _19752_, _19751_);
  and (_19755_, _19754_, _06114_);
  and (_19756_, _19755_, _19750_);
  and (_19757_, _15395_, _07856_);
  or (_19758_, _19757_, _19721_);
  and (_19759_, _19758_, _05787_);
  or (_19760_, _19759_, _11136_);
  or (_19761_, _19760_, _19756_);
  and (_19762_, _15413_, _07856_);
  or (_19763_, _19721_, _07127_);
  or (_19765_, _19763_, _19762_);
  or (_19766_, _19724_, _06111_);
  and (_19767_, _19766_, _07125_);
  and (_19768_, _19767_, _19765_);
  and (_19769_, _19768_, _19761_);
  and (_19770_, _10295_, _07856_);
  or (_19771_, _19770_, _19721_);
  and (_19772_, _19771_, _06402_);
  or (_19773_, _19772_, _19769_);
  and (_19774_, _19773_, _07132_);
  or (_19776_, _19774_, _19726_);
  and (_19777_, _19776_, _07130_);
  and (_19778_, _19732_, _06411_);
  and (_19779_, _19778_, _19722_);
  or (_19780_, _19779_, _06303_);
  or (_19781_, _19780_, _19777_);
  and (_19782_, _15410_, _07856_);
  or (_19783_, _19721_, _08819_);
  or (_19784_, _19783_, _19782_);
  and (_19785_, _19784_, _08824_);
  and (_19787_, _19785_, _19781_);
  nor (_19788_, _10294_, _11137_);
  or (_19789_, _19788_, _19721_);
  and (_19790_, _19789_, _06396_);
  or (_19791_, _19790_, _06433_);
  or (_19792_, _19791_, _19787_);
  or (_19793_, _19728_, _06829_);
  and (_19794_, _19793_, _06444_);
  and (_19795_, _19794_, _19792_);
  and (_19796_, _15478_, _07856_);
  or (_19798_, _19796_, _19721_);
  and (_19799_, _19798_, _06440_);
  or (_19800_, _19799_, _01321_);
  or (_19801_, _19800_, _19795_);
  or (_19802_, _01317_, \oc8051_golden_model_1.PCON [6]);
  and (_19803_, _19802_, _43100_);
  and (_43618_, _19803_, _19801_);
  not (_19804_, \oc8051_golden_model_1.TMOD [0]);
  nor (_19805_, _01317_, _19804_);
  nand (_19806_, _10276_, _07812_);
  nor (_19808_, _07812_, _19804_);
  nor (_19809_, _19808_, _07130_);
  nand (_19810_, _19809_, _19806_);
  and (_19811_, _07812_, _07049_);
  or (_19812_, _19811_, _19808_);
  or (_19813_, _19812_, _06132_);
  nor (_19814_, _08211_, _11214_);
  or (_19815_, _19814_, _19808_);
  or (_19816_, _19815_, _06161_);
  and (_19817_, _07812_, \oc8051_golden_model_1.ACC [0]);
  or (_19819_, _19817_, _19808_);
  and (_19820_, _19819_, _07056_);
  nor (_19821_, _07056_, _19804_);
  or (_19822_, _19821_, _06160_);
  or (_19823_, _19822_, _19820_);
  and (_19824_, _19823_, _07075_);
  and (_19825_, _19824_, _19816_);
  and (_19826_, _19812_, _06217_);
  or (_19827_, _19826_, _19825_);
  and (_19828_, _19827_, _06229_);
  and (_19830_, _19819_, _06220_);
  or (_19831_, _19830_, _09842_);
  or (_19832_, _19831_, _19828_);
  and (_19833_, _19832_, _19813_);
  or (_19834_, _19833_, _06116_);
  and (_19835_, _09160_, _07812_);
  or (_19836_, _19808_, _06117_);
  or (_19837_, _19836_, _19835_);
  and (_19838_, _19837_, _19834_);
  or (_19839_, _19838_, _05787_);
  and (_19841_, _14260_, _07812_);
  or (_19842_, _19808_, _06114_);
  or (_19843_, _19842_, _19841_);
  and (_19844_, _19843_, _06111_);
  and (_19845_, _19844_, _19839_);
  and (_19846_, _07812_, _08708_);
  or (_19847_, _19846_, _19808_);
  and (_19848_, _19847_, _06110_);
  or (_19849_, _19848_, _06297_);
  or (_19850_, _19849_, _19845_);
  and (_19852_, _14275_, _07812_);
  or (_19853_, _19808_, _07127_);
  or (_19854_, _19853_, _19852_);
  and (_19855_, _19854_, _07125_);
  and (_19856_, _19855_, _19850_);
  nor (_19857_, _12321_, _11214_);
  or (_19858_, _19857_, _19808_);
  and (_19859_, _19806_, _06402_);
  and (_19860_, _19859_, _19858_);
  or (_19861_, _19860_, _19856_);
  and (_19864_, _19861_, _07132_);
  nand (_19865_, _19847_, _06306_);
  nor (_19866_, _19865_, _19814_);
  or (_19867_, _19866_, _06411_);
  or (_19868_, _19867_, _19864_);
  and (_19869_, _19868_, _19810_);
  or (_19870_, _19869_, _06303_);
  and (_19871_, _14167_, _07812_);
  or (_19872_, _19808_, _08819_);
  or (_19873_, _19872_, _19871_);
  and (_19876_, _19873_, _08824_);
  and (_19877_, _19876_, _19870_);
  and (_19878_, _19858_, _06396_);
  or (_19879_, _19878_, _19287_);
  or (_19880_, _19879_, _19877_);
  or (_19881_, _19815_, _06630_);
  and (_19882_, _19881_, _01317_);
  and (_19883_, _19882_, _19880_);
  or (_19884_, _19883_, _19805_);
  and (_43619_, _19884_, _43100_);
  and (_19887_, _11214_, \oc8051_golden_model_1.TMOD [1]);
  nor (_19888_, _10277_, _11214_);
  or (_19889_, _19888_, _19887_);
  or (_19890_, _19889_, _08824_);
  or (_19891_, _14442_, _11214_);
  or (_19892_, _07812_, \oc8051_golden_model_1.TMOD [1]);
  and (_19893_, _19892_, _05787_);
  and (_19894_, _19893_, _19891_);
  and (_19895_, _09115_, _07812_);
  or (_19896_, _19887_, _06117_);
  or (_19899_, _19896_, _19895_);
  and (_19900_, _14363_, _07812_);
  not (_19901_, _19900_);
  and (_19902_, _19901_, _19892_);
  or (_19903_, _19902_, _06161_);
  and (_19904_, _07812_, \oc8051_golden_model_1.ACC [1]);
  or (_19905_, _19904_, _19887_);
  and (_19906_, _19905_, _07056_);
  and (_19907_, _07057_, \oc8051_golden_model_1.TMOD [1]);
  or (_19908_, _19907_, _06160_);
  or (_19911_, _19908_, _19906_);
  and (_19912_, _19911_, _07075_);
  and (_19913_, _19912_, _19903_);
  and (_19914_, _07812_, _07306_);
  or (_19915_, _19914_, _19887_);
  and (_19916_, _19915_, _06217_);
  or (_19917_, _19916_, _19913_);
  and (_19918_, _19917_, _06229_);
  and (_19919_, _19905_, _06220_);
  or (_19920_, _19919_, _09842_);
  or (_19923_, _19920_, _19918_);
  or (_19924_, _19915_, _06132_);
  and (_19925_, _19924_, _19923_);
  or (_19926_, _19925_, _06116_);
  and (_19927_, _19926_, _06114_);
  and (_19928_, _19927_, _19899_);
  or (_19929_, _19928_, _19894_);
  and (_19930_, _19929_, _06298_);
  or (_19931_, _14346_, _11214_);
  and (_19932_, _19931_, _06297_);
  nand (_19935_, _07812_, _06945_);
  and (_19936_, _19935_, _06110_);
  or (_19937_, _19936_, _19932_);
  and (_19938_, _19937_, _19892_);
  or (_19939_, _19938_, _06402_);
  or (_19940_, _19939_, _19930_);
  nand (_19941_, _10275_, _07812_);
  and (_19942_, _19941_, _19889_);
  or (_19943_, _19942_, _07125_);
  and (_19944_, _19943_, _07132_);
  and (_19946_, _19944_, _19940_);
  or (_19947_, _14344_, _11214_);
  and (_19948_, _19892_, _06306_);
  and (_19949_, _19948_, _19947_);
  or (_19950_, _19949_, _06411_);
  or (_19951_, _19950_, _19946_);
  nor (_19952_, _19887_, _07130_);
  nand (_19953_, _19952_, _19941_);
  and (_19954_, _19953_, _08819_);
  and (_19955_, _19954_, _19951_);
  or (_19957_, _19935_, _08176_);
  and (_19958_, _19892_, _06303_);
  and (_19959_, _19958_, _19957_);
  or (_19960_, _19959_, _06396_);
  or (_19961_, _19960_, _19955_);
  and (_19962_, _19961_, _19890_);
  or (_19963_, _19962_, _06433_);
  or (_19964_, _19902_, _06829_);
  and (_19965_, _19964_, _06444_);
  and (_19966_, _19965_, _19963_);
  or (_19968_, _19900_, _19887_);
  and (_19969_, _19968_, _06440_);
  or (_19970_, _19969_, _01321_);
  or (_19971_, _19970_, _19966_);
  or (_19972_, _01317_, \oc8051_golden_model_1.TMOD [1]);
  and (_19973_, _19972_, _43100_);
  and (_43621_, _19973_, _19971_);
  and (_19974_, _01321_, \oc8051_golden_model_1.TMOD [2]);
  and (_19975_, _11214_, \oc8051_golden_model_1.TMOD [2]);
  and (_19976_, _09211_, _07812_);
  or (_19978_, _19976_, _19975_);
  and (_19979_, _19978_, _06116_);
  and (_19980_, _14542_, _07812_);
  or (_19981_, _19980_, _19975_);
  or (_19982_, _19981_, _06161_);
  and (_19983_, _07812_, \oc8051_golden_model_1.ACC [2]);
  or (_19984_, _19983_, _19975_);
  and (_19985_, _19984_, _07056_);
  and (_19986_, _07057_, \oc8051_golden_model_1.TMOD [2]);
  or (_19987_, _19986_, _06160_);
  or (_19989_, _19987_, _19985_);
  and (_19990_, _19989_, _07075_);
  and (_19991_, _19990_, _19982_);
  and (_19992_, _07812_, _07708_);
  or (_19993_, _19992_, _19975_);
  and (_19994_, _19993_, _06217_);
  or (_19995_, _19994_, _19991_);
  and (_19996_, _19995_, _06229_);
  and (_19997_, _19984_, _06220_);
  or (_19998_, _19997_, _09842_);
  or (_20000_, _19998_, _19996_);
  or (_20001_, _19993_, _06132_);
  and (_20002_, _20001_, _06117_);
  and (_20003_, _20002_, _20000_);
  or (_20004_, _20003_, _05787_);
  or (_20005_, _20004_, _19979_);
  and (_20006_, _14630_, _07812_);
  or (_20007_, _20006_, _19975_);
  or (_20008_, _20007_, _06114_);
  and (_20009_, _20008_, _06111_);
  and (_20011_, _20009_, _20005_);
  and (_20012_, _07812_, _08768_);
  or (_20013_, _20012_, _19975_);
  and (_20014_, _20013_, _06110_);
  or (_20015_, _20014_, _06297_);
  or (_20016_, _20015_, _20011_);
  and (_20017_, _14646_, _07812_);
  or (_20018_, _19975_, _07127_);
  or (_20019_, _20018_, _20017_);
  and (_20020_, _20019_, _07125_);
  and (_20022_, _20020_, _20016_);
  and (_20023_, _10282_, _07812_);
  or (_20024_, _20023_, _19975_);
  and (_20025_, _20024_, _06402_);
  or (_20026_, _20025_, _20022_);
  and (_20027_, _20026_, _07132_);
  or (_20028_, _19975_, _08248_);
  and (_20029_, _20013_, _06306_);
  and (_20030_, _20029_, _20028_);
  or (_20031_, _20030_, _20027_);
  and (_20033_, _20031_, _07130_);
  and (_20034_, _19984_, _06411_);
  and (_20035_, _20034_, _20028_);
  or (_20036_, _20035_, _06303_);
  or (_20037_, _20036_, _20033_);
  and (_20038_, _14643_, _07812_);
  or (_20039_, _19975_, _08819_);
  or (_20040_, _20039_, _20038_);
  and (_20041_, _20040_, _08824_);
  and (_20042_, _20041_, _20037_);
  nor (_20044_, _10281_, _11214_);
  or (_20045_, _20044_, _19975_);
  and (_20046_, _20045_, _06396_);
  or (_20047_, _20046_, _20042_);
  and (_20048_, _20047_, _06829_);
  and (_20049_, _19981_, _06433_);
  or (_20050_, _20049_, _06440_);
  or (_20051_, _20050_, _20048_);
  and (_20052_, _14710_, _07812_);
  or (_20053_, _19975_, _06444_);
  or (_20055_, _20053_, _20052_);
  and (_20056_, _20055_, _01317_);
  and (_20057_, _20056_, _20051_);
  or (_20058_, _20057_, _19974_);
  and (_43622_, _20058_, _43100_);
  and (_20059_, _11214_, \oc8051_golden_model_1.TMOD [3]);
  and (_20060_, _14738_, _07812_);
  or (_20061_, _20060_, _20059_);
  or (_20062_, _20061_, _06161_);
  and (_20063_, _07812_, \oc8051_golden_model_1.ACC [3]);
  or (_20065_, _20063_, _20059_);
  and (_20066_, _20065_, _07056_);
  and (_20067_, _07057_, \oc8051_golden_model_1.TMOD [3]);
  or (_20068_, _20067_, _06160_);
  or (_20069_, _20068_, _20066_);
  and (_20070_, _20069_, _07075_);
  and (_20071_, _20070_, _20062_);
  and (_20072_, _07812_, _07544_);
  or (_20073_, _20072_, _20059_);
  and (_20074_, _20073_, _06217_);
  or (_20076_, _20074_, _20071_);
  and (_20077_, _20076_, _06229_);
  and (_20078_, _20065_, _06220_);
  or (_20079_, _20078_, _09842_);
  or (_20080_, _20079_, _20077_);
  or (_20081_, _20073_, _06132_);
  and (_20082_, _20081_, _20080_);
  or (_20083_, _20082_, _06116_);
  and (_20084_, _09210_, _07812_);
  or (_20085_, _20059_, _06117_);
  or (_20087_, _20085_, _20084_);
  and (_20088_, _20087_, _06114_);
  and (_20089_, _20088_, _20083_);
  and (_20090_, _14825_, _07812_);
  or (_20091_, _20090_, _20059_);
  and (_20092_, _20091_, _05787_);
  or (_20093_, _20092_, _11136_);
  or (_20094_, _20093_, _20089_);
  and (_20095_, _14727_, _07812_);
  or (_20096_, _20059_, _07127_);
  or (_20098_, _20096_, _20095_);
  and (_20099_, _07812_, _08712_);
  or (_20100_, _20099_, _20059_);
  or (_20101_, _20100_, _06111_);
  and (_20102_, _20101_, _07125_);
  and (_20103_, _20102_, _20098_);
  and (_20104_, _20103_, _20094_);
  and (_20105_, _12318_, _07812_);
  or (_20106_, _20105_, _20059_);
  and (_20107_, _20106_, _06402_);
  or (_20109_, _20107_, _20104_);
  and (_20110_, _20109_, _07132_);
  or (_20111_, _20059_, _08140_);
  and (_20112_, _20100_, _06306_);
  and (_20113_, _20112_, _20111_);
  or (_20114_, _20113_, _20110_);
  and (_20115_, _20114_, _07130_);
  and (_20116_, _20065_, _06411_);
  and (_20117_, _20116_, _20111_);
  or (_20118_, _20117_, _06303_);
  or (_20120_, _20118_, _20115_);
  and (_20121_, _14724_, _07812_);
  or (_20122_, _20059_, _08819_);
  or (_20123_, _20122_, _20121_);
  and (_20124_, _20123_, _08824_);
  and (_20125_, _20124_, _20120_);
  nor (_20126_, _10273_, _11214_);
  or (_20127_, _20126_, _20059_);
  and (_20128_, _20127_, _06396_);
  or (_20129_, _20128_, _06433_);
  or (_20131_, _20129_, _20125_);
  or (_20132_, _20061_, _06829_);
  and (_20133_, _20132_, _06444_);
  and (_20134_, _20133_, _20131_);
  and (_20135_, _14897_, _07812_);
  or (_20136_, _20135_, _20059_);
  and (_20137_, _20136_, _06440_);
  or (_20138_, _20137_, _01321_);
  or (_20139_, _20138_, _20134_);
  or (_20140_, _01317_, \oc8051_golden_model_1.TMOD [3]);
  and (_20142_, _20140_, _43100_);
  and (_43623_, _20142_, _20139_);
  and (_20143_, _11214_, \oc8051_golden_model_1.TMOD [4]);
  and (_20144_, _08336_, _07812_);
  or (_20145_, _20144_, _20143_);
  or (_20146_, _20145_, _06132_);
  and (_20147_, _14928_, _07812_);
  or (_20148_, _20147_, _20143_);
  or (_20149_, _20148_, _06161_);
  and (_20150_, _07812_, \oc8051_golden_model_1.ACC [4]);
  or (_20152_, _20150_, _20143_);
  and (_20153_, _20152_, _07056_);
  and (_20154_, _07057_, \oc8051_golden_model_1.TMOD [4]);
  or (_20155_, _20154_, _06160_);
  or (_20156_, _20155_, _20153_);
  and (_20157_, _20156_, _07075_);
  and (_20158_, _20157_, _20149_);
  and (_20159_, _20145_, _06217_);
  or (_20160_, _20159_, _20158_);
  and (_20161_, _20160_, _06229_);
  and (_20163_, _20152_, _06220_);
  or (_20164_, _20163_, _09842_);
  or (_20165_, _20164_, _20161_);
  and (_20166_, _20165_, _20146_);
  or (_20167_, _20166_, _06116_);
  and (_20168_, _09209_, _07812_);
  or (_20169_, _20143_, _06117_);
  or (_20170_, _20169_, _20168_);
  and (_20171_, _20170_, _06114_);
  and (_20172_, _20171_, _20167_);
  and (_20174_, _15013_, _07812_);
  or (_20175_, _20174_, _20143_);
  and (_20176_, _20175_, _05787_);
  or (_20177_, _20176_, _20172_);
  or (_20178_, _20177_, _11136_);
  and (_20179_, _15029_, _07812_);
  or (_20180_, _20143_, _07127_);
  or (_20181_, _20180_, _20179_);
  and (_20182_, _08715_, _07812_);
  or (_20183_, _20182_, _20143_);
  or (_20185_, _20183_, _06111_);
  and (_20186_, _20185_, _07125_);
  and (_20187_, _20186_, _20181_);
  and (_20188_, _20187_, _20178_);
  and (_20189_, _10289_, _07812_);
  or (_20190_, _20189_, _20143_);
  and (_20191_, _20190_, _06402_);
  or (_20192_, _20191_, _20188_);
  and (_20193_, _20192_, _07132_);
  or (_20194_, _20143_, _08339_);
  and (_20196_, _20183_, _06306_);
  and (_20197_, _20196_, _20194_);
  or (_20198_, _20197_, _20193_);
  and (_20199_, _20198_, _07130_);
  and (_20200_, _20152_, _06411_);
  and (_20201_, _20200_, _20194_);
  or (_20202_, _20201_, _06303_);
  or (_20203_, _20202_, _20199_);
  and (_20204_, _15026_, _07812_);
  or (_20205_, _20143_, _08819_);
  or (_20207_, _20205_, _20204_);
  and (_20208_, _20207_, _08824_);
  and (_20209_, _20208_, _20203_);
  nor (_20210_, _10288_, _11214_);
  or (_20211_, _20210_, _20143_);
  and (_20212_, _20211_, _06396_);
  or (_20213_, _20212_, _06433_);
  or (_20214_, _20213_, _20209_);
  or (_20215_, _20148_, _06829_);
  and (_20216_, _20215_, _06444_);
  and (_20218_, _20216_, _20214_);
  and (_20219_, _15087_, _07812_);
  or (_20220_, _20219_, _20143_);
  and (_20221_, _20220_, _06440_);
  or (_20222_, _20221_, _01321_);
  or (_20223_, _20222_, _20218_);
  or (_20224_, _01317_, \oc8051_golden_model_1.TMOD [4]);
  and (_20225_, _20224_, _43100_);
  and (_43624_, _20225_, _20223_);
  and (_20226_, _11214_, \oc8051_golden_model_1.TMOD [5]);
  and (_20228_, _15119_, _07812_);
  or (_20229_, _20228_, _20226_);
  or (_20230_, _20229_, _06161_);
  and (_20231_, _07812_, \oc8051_golden_model_1.ACC [5]);
  or (_20232_, _20231_, _20226_);
  and (_20233_, _20232_, _07056_);
  and (_20234_, _07057_, \oc8051_golden_model_1.TMOD [5]);
  or (_20235_, _20234_, _06160_);
  or (_20236_, _20235_, _20233_);
  and (_20237_, _20236_, _07075_);
  and (_20239_, _20237_, _20230_);
  and (_20240_, _08101_, _07812_);
  or (_20241_, _20240_, _20226_);
  and (_20242_, _20241_, _06217_);
  or (_20243_, _20242_, _20239_);
  and (_20244_, _20243_, _06229_);
  and (_20245_, _20232_, _06220_);
  or (_20246_, _20245_, _09842_);
  or (_20247_, _20246_, _20244_);
  or (_20248_, _20241_, _06132_);
  and (_20250_, _20248_, _20247_);
  or (_20251_, _20250_, _06116_);
  and (_20252_, _09208_, _07812_);
  or (_20253_, _20226_, _06117_);
  or (_20254_, _20253_, _20252_);
  and (_20255_, _20254_, _06114_);
  and (_20256_, _20255_, _20251_);
  and (_20257_, _15203_, _07812_);
  or (_20258_, _20257_, _20226_);
  and (_20259_, _20258_, _05787_);
  or (_20261_, _20259_, _11136_);
  or (_20262_, _20261_, _20256_);
  and (_20263_, _15219_, _07812_);
  or (_20264_, _20226_, _07127_);
  or (_20265_, _20264_, _20263_);
  and (_20266_, _08736_, _07812_);
  or (_20267_, _20266_, _20226_);
  or (_20268_, _20267_, _06111_);
  and (_20269_, _20268_, _07125_);
  and (_20270_, _20269_, _20265_);
  and (_20272_, _20270_, _20262_);
  and (_20273_, _12325_, _07812_);
  or (_20274_, _20273_, _20226_);
  and (_20275_, _20274_, _06402_);
  or (_20276_, _20275_, _20272_);
  and (_20277_, _20276_, _07132_);
  or (_20278_, _20226_, _08104_);
  and (_20279_, _20267_, _06306_);
  and (_20280_, _20279_, _20278_);
  or (_20281_, _20280_, _20277_);
  and (_20283_, _20281_, _07130_);
  and (_20284_, _20232_, _06411_);
  and (_20285_, _20284_, _20278_);
  or (_20286_, _20285_, _06303_);
  or (_20287_, _20286_, _20283_);
  and (_20288_, _15216_, _07812_);
  or (_20289_, _20226_, _08819_);
  or (_20290_, _20289_, _20288_);
  and (_20291_, _20290_, _08824_);
  and (_20292_, _20291_, _20287_);
  nor (_20294_, _10269_, _11214_);
  or (_20295_, _20294_, _20226_);
  and (_20296_, _20295_, _06396_);
  or (_20297_, _20296_, _06433_);
  or (_20298_, _20297_, _20292_);
  or (_20299_, _20229_, _06829_);
  and (_20300_, _20299_, _06444_);
  and (_20301_, _20300_, _20298_);
  and (_20302_, _15275_, _07812_);
  or (_20303_, _20302_, _20226_);
  and (_20305_, _20303_, _06440_);
  or (_20306_, _20305_, _01321_);
  or (_20307_, _20306_, _20301_);
  or (_20308_, _01317_, \oc8051_golden_model_1.TMOD [5]);
  and (_20309_, _20308_, _43100_);
  and (_43625_, _20309_, _20307_);
  and (_20310_, _11214_, \oc8051_golden_model_1.TMOD [6]);
  and (_20311_, _15300_, _07812_);
  or (_20312_, _20311_, _20310_);
  or (_20313_, _20312_, _06161_);
  and (_20315_, _07812_, \oc8051_golden_model_1.ACC [6]);
  or (_20316_, _20315_, _20310_);
  and (_20317_, _20316_, _07056_);
  and (_20318_, _07057_, \oc8051_golden_model_1.TMOD [6]);
  or (_20319_, _20318_, _06160_);
  or (_20320_, _20319_, _20317_);
  and (_20321_, _20320_, _07075_);
  and (_20322_, _20321_, _20313_);
  and (_20323_, _08012_, _07812_);
  or (_20324_, _20323_, _20310_);
  and (_20326_, _20324_, _06217_);
  or (_20327_, _20326_, _20322_);
  and (_20328_, _20327_, _06229_);
  and (_20329_, _20316_, _06220_);
  or (_20330_, _20329_, _09842_);
  or (_20331_, _20330_, _20328_);
  or (_20332_, _20324_, _06132_);
  and (_20333_, _20332_, _20331_);
  or (_20334_, _20333_, _06116_);
  and (_20335_, _09207_, _07812_);
  or (_20337_, _20310_, _06117_);
  or (_20338_, _20337_, _20335_);
  and (_20339_, _20338_, _06114_);
  and (_20340_, _20339_, _20334_);
  and (_20341_, _15395_, _07812_);
  or (_20342_, _20341_, _20310_);
  and (_20343_, _20342_, _05787_);
  or (_20344_, _20343_, _11136_);
  or (_20345_, _20344_, _20340_);
  and (_20346_, _15413_, _07812_);
  or (_20348_, _20310_, _07127_);
  or (_20349_, _20348_, _20346_);
  and (_20350_, _15402_, _07812_);
  or (_20351_, _20350_, _20310_);
  or (_20352_, _20351_, _06111_);
  and (_20353_, _20352_, _07125_);
  and (_20354_, _20353_, _20349_);
  and (_20355_, _20354_, _20345_);
  and (_20356_, _10295_, _07812_);
  or (_20357_, _20356_, _20310_);
  and (_20359_, _20357_, _06402_);
  or (_20360_, _20359_, _20355_);
  and (_20361_, _20360_, _07132_);
  or (_20362_, _20310_, _08015_);
  and (_20363_, _20351_, _06306_);
  and (_20364_, _20363_, _20362_);
  or (_20365_, _20364_, _20361_);
  and (_20366_, _20365_, _07130_);
  and (_20367_, _20316_, _06411_);
  and (_20368_, _20367_, _20362_);
  or (_20370_, _20368_, _06303_);
  or (_20371_, _20370_, _20366_);
  and (_20372_, _15410_, _07812_);
  or (_20373_, _20310_, _08819_);
  or (_20374_, _20373_, _20372_);
  and (_20375_, _20374_, _08824_);
  and (_20376_, _20375_, _20371_);
  nor (_20377_, _10294_, _11214_);
  or (_20378_, _20377_, _20310_);
  and (_20379_, _20378_, _06396_);
  or (_20381_, _20379_, _06433_);
  or (_20382_, _20381_, _20376_);
  or (_20383_, _20312_, _06829_);
  and (_20384_, _20383_, _06444_);
  and (_20385_, _20384_, _20382_);
  and (_20386_, _15478_, _07812_);
  or (_20387_, _20386_, _20310_);
  and (_20388_, _20387_, _06440_);
  or (_20389_, _20388_, _01321_);
  or (_20390_, _20389_, _20385_);
  or (_20392_, _01317_, \oc8051_golden_model_1.TMOD [6]);
  and (_20393_, _20392_, _43100_);
  and (_43626_, _20393_, _20390_);
  not (_20394_, \oc8051_golden_model_1.DPL [0]);
  nor (_20395_, _01317_, _20394_);
  nand (_20396_, _10276_, _07849_);
  nor (_20397_, _07849_, _20394_);
  nor (_20398_, _20397_, _07130_);
  nand (_20399_, _20398_, _20396_);
  and (_20400_, _07849_, _07049_);
  or (_20402_, _20400_, _20397_);
  or (_20403_, _20402_, _06132_);
  and (_20404_, _07849_, \oc8051_golden_model_1.ACC [0]);
  or (_20405_, _20404_, _20397_);
  or (_20406_, _20405_, _06229_);
  nor (_20407_, _08211_, _11371_);
  or (_20408_, _20407_, _20397_);
  or (_20409_, _20408_, _06161_);
  and (_20410_, _20405_, _07056_);
  nor (_20411_, _07056_, _20394_);
  or (_20413_, _20411_, _06160_);
  or (_20414_, _20413_, _20410_);
  and (_20415_, _20414_, _07075_);
  and (_20416_, _20415_, _20409_);
  and (_20417_, _20402_, _06217_);
  or (_20418_, _20417_, _06220_);
  or (_20419_, _20418_, _20416_);
  and (_20420_, _20419_, _20406_);
  or (_20421_, _20420_, _11311_);
  nand (_20422_, _11311_, \oc8051_golden_model_1.DPL [0]);
  and (_20424_, _20422_, _11296_);
  and (_20425_, _20424_, _20421_);
  nor (_20426_, _06758_, _11296_);
  or (_20427_, _20426_, _09842_);
  or (_20428_, _20427_, _20425_);
  and (_20429_, _20428_, _20403_);
  or (_20430_, _20429_, _06116_);
  and (_20431_, _09160_, _07849_);
  or (_20432_, _20397_, _06117_);
  or (_20433_, _20432_, _20431_);
  and (_20435_, _20433_, _20430_);
  or (_20436_, _20435_, _05787_);
  and (_20437_, _14260_, _07849_);
  or (_20438_, _20437_, _20397_);
  or (_20439_, _20438_, _06114_);
  and (_20440_, _20439_, _06111_);
  and (_20441_, _20440_, _20436_);
  and (_20442_, _07849_, _08708_);
  or (_20443_, _20442_, _20397_);
  and (_20444_, _20443_, _06110_);
  or (_20446_, _20444_, _06297_);
  or (_20447_, _20446_, _20441_);
  and (_20448_, _14275_, _07849_);
  or (_20449_, _20448_, _20397_);
  or (_20450_, _20449_, _07127_);
  and (_20451_, _20450_, _07125_);
  and (_20452_, _20451_, _20447_);
  nor (_20453_, _12321_, _11371_);
  or (_20454_, _20453_, _20397_);
  and (_20455_, _20396_, _06402_);
  and (_20457_, _20455_, _20454_);
  or (_20458_, _20457_, _20452_);
  and (_20459_, _20458_, _07132_);
  nand (_20460_, _20443_, _06306_);
  nor (_20461_, _20460_, _20407_);
  or (_20462_, _20461_, _06411_);
  or (_20463_, _20462_, _20459_);
  and (_20464_, _20463_, _20399_);
  or (_20465_, _20464_, _06303_);
  and (_20466_, _14167_, _07849_);
  or (_20468_, _20397_, _08819_);
  or (_20469_, _20468_, _20466_);
  and (_20470_, _20469_, _08824_);
  and (_20471_, _20470_, _20465_);
  and (_20472_, _20454_, _06396_);
  or (_20473_, _20472_, _19287_);
  or (_20474_, _20473_, _20471_);
  or (_20475_, _20408_, _06630_);
  and (_20476_, _20475_, _01317_);
  and (_20477_, _20476_, _20474_);
  or (_20479_, _20477_, _20395_);
  and (_43628_, _20479_, _43100_);
  not (_20480_, \oc8051_golden_model_1.DPL [1]);
  nor (_20481_, _01317_, _20480_);
  and (_20482_, _09115_, _07849_);
  nor (_20483_, _07849_, _20480_);
  or (_20484_, _20483_, _20482_);
  and (_20485_, _20484_, _06116_);
  or (_20486_, _07849_, \oc8051_golden_model_1.DPL [1]);
  and (_20487_, _14363_, _07849_);
  not (_20489_, _20487_);
  and (_20490_, _20489_, _20486_);
  or (_20491_, _20490_, _06161_);
  and (_20492_, _07849_, \oc8051_golden_model_1.ACC [1]);
  or (_20493_, _20492_, _20483_);
  and (_20494_, _20493_, _07056_);
  nor (_20495_, _07056_, _20480_);
  or (_20496_, _20495_, _06160_);
  or (_20497_, _20496_, _20494_);
  and (_20498_, _20497_, _07075_);
  and (_20500_, _20498_, _20491_);
  and (_20501_, _07849_, _07306_);
  or (_20502_, _20501_, _20483_);
  and (_20503_, _20502_, _06217_);
  or (_20504_, _20503_, _06220_);
  or (_20505_, _20504_, _20500_);
  or (_20506_, _20493_, _06229_);
  and (_20507_, _20506_, _11312_);
  and (_20508_, _20507_, _20505_);
  nor (_20509_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_20511_, _20509_, _11316_);
  and (_20512_, _20511_, _11311_);
  or (_20513_, _20512_, _20508_);
  and (_20514_, _20513_, _11296_);
  nor (_20515_, _06945_, _11296_);
  or (_20516_, _20515_, _09842_);
  or (_20517_, _20516_, _20514_);
  or (_20518_, _20502_, _06132_);
  and (_20519_, _20518_, _06117_);
  and (_20520_, _20519_, _20517_);
  or (_20522_, _20520_, _20485_);
  and (_20523_, _20522_, _06114_);
  or (_20524_, _14442_, _11371_);
  and (_20525_, _20486_, _05787_);
  and (_20526_, _20525_, _20524_);
  or (_20527_, _20526_, _20523_);
  and (_20528_, _20527_, _06298_);
  or (_20529_, _14346_, _11371_);
  and (_20530_, _20529_, _06297_);
  nand (_20531_, _07849_, _06945_);
  and (_20533_, _20531_, _06110_);
  or (_20534_, _20533_, _20530_);
  and (_20535_, _20534_, _20486_);
  or (_20536_, _20535_, _06402_);
  or (_20537_, _20536_, _20528_);
  nor (_20538_, _10277_, _11371_);
  or (_20539_, _20538_, _20483_);
  nand (_20540_, _10275_, _07849_);
  and (_20541_, _20540_, _20539_);
  or (_20542_, _20541_, _07125_);
  and (_20544_, _20542_, _07132_);
  and (_20545_, _20544_, _20537_);
  or (_20546_, _14344_, _11371_);
  and (_20547_, _20486_, _06306_);
  and (_20548_, _20547_, _20546_);
  or (_20549_, _20548_, _06411_);
  or (_20550_, _20549_, _20545_);
  nor (_20551_, _20483_, _07130_);
  nand (_20552_, _20551_, _20540_);
  and (_20553_, _20552_, _08819_);
  and (_20555_, _20553_, _20550_);
  or (_20556_, _20531_, _08176_);
  and (_20557_, _20486_, _06303_);
  and (_20558_, _20557_, _20556_);
  or (_20559_, _20558_, _06396_);
  or (_20560_, _20559_, _20555_);
  or (_20561_, _20539_, _08824_);
  and (_20562_, _20561_, _06829_);
  and (_20563_, _20562_, _20560_);
  and (_20564_, _20490_, _06433_);
  or (_20566_, _20564_, _06440_);
  or (_20567_, _20566_, _20563_);
  or (_20568_, _20483_, _06444_);
  or (_20569_, _20568_, _20487_);
  and (_20570_, _20569_, _01317_);
  and (_20571_, _20570_, _20567_);
  or (_20572_, _20571_, _20481_);
  and (_43629_, _20572_, _43100_);
  not (_20573_, \oc8051_golden_model_1.DPL [2]);
  nor (_20574_, _01317_, _20573_);
  nor (_20576_, _07849_, _20573_);
  or (_20577_, _20576_, _08248_);
  and (_20578_, _07849_, _08768_);
  or (_20579_, _20578_, _20576_);
  and (_20580_, _20579_, _06306_);
  and (_20581_, _20580_, _20577_);
  and (_20582_, _07849_, _07708_);
  or (_20583_, _20582_, _20576_);
  or (_20584_, _20583_, _07075_);
  and (_20585_, _14542_, _07849_);
  or (_20587_, _20585_, _20576_);
  and (_20588_, _20587_, _06160_);
  nor (_20589_, _07056_, _20573_);
  and (_20590_, _07849_, \oc8051_golden_model_1.ACC [2]);
  or (_20591_, _20590_, _20576_);
  and (_20592_, _20591_, _07056_);
  or (_20593_, _20592_, _20589_);
  and (_20594_, _20593_, _06161_);
  or (_20595_, _20594_, _06217_);
  or (_20596_, _20595_, _20588_);
  and (_20598_, _20596_, _20584_);
  or (_20599_, _20598_, _06220_);
  or (_20600_, _20591_, _06229_);
  and (_20601_, _20600_, _11312_);
  and (_20602_, _20601_, _20599_);
  nor (_20603_, _11316_, \oc8051_golden_model_1.DPL [2]);
  nor (_20604_, _20603_, _11317_);
  and (_20605_, _20604_, _11311_);
  or (_20606_, _20605_, _20602_);
  and (_20607_, _20606_, _11296_);
  nor (_20609_, _06521_, _11296_);
  or (_20610_, _20609_, _09842_);
  or (_20611_, _20610_, _20607_);
  or (_20612_, _20583_, _06132_);
  and (_20613_, _20612_, _20611_);
  or (_20614_, _20613_, _06116_);
  and (_20615_, _09211_, _07849_);
  or (_20616_, _20576_, _06117_);
  or (_20617_, _20616_, _20615_);
  and (_20618_, _20617_, _06114_);
  and (_20620_, _20618_, _20614_);
  and (_20621_, _14630_, _07849_);
  or (_20622_, _20621_, _20576_);
  and (_20623_, _20622_, _05787_);
  or (_20624_, _20623_, _11136_);
  or (_20625_, _20624_, _20620_);
  and (_20626_, _14646_, _07849_);
  or (_20627_, _20576_, _07127_);
  or (_20628_, _20627_, _20626_);
  or (_20629_, _20579_, _06111_);
  and (_20631_, _20629_, _07125_);
  and (_20632_, _20631_, _20628_);
  and (_20633_, _20632_, _20625_);
  and (_20634_, _10282_, _07849_);
  or (_20635_, _20634_, _20576_);
  and (_20636_, _20635_, _06402_);
  or (_20637_, _20636_, _20633_);
  and (_20638_, _20637_, _07132_);
  or (_20639_, _20638_, _20581_);
  and (_20640_, _20639_, _07130_);
  and (_20642_, _20591_, _06411_);
  and (_20643_, _20642_, _20577_);
  or (_20644_, _20643_, _06303_);
  or (_20645_, _20644_, _20640_);
  and (_20646_, _14643_, _07849_);
  or (_20647_, _20576_, _08819_);
  or (_20648_, _20647_, _20646_);
  and (_20649_, _20648_, _08824_);
  and (_20650_, _20649_, _20645_);
  nor (_20651_, _10281_, _11371_);
  or (_20653_, _20651_, _20576_);
  and (_20654_, _20653_, _06396_);
  or (_20655_, _20654_, _20650_);
  and (_20656_, _20655_, _06829_);
  and (_20657_, _20587_, _06433_);
  or (_20658_, _20657_, _06440_);
  or (_20659_, _20658_, _20656_);
  and (_20660_, _14710_, _07849_);
  or (_20661_, _20576_, _06444_);
  or (_20662_, _20661_, _20660_);
  and (_20664_, _20662_, _01317_);
  and (_20665_, _20664_, _20659_);
  or (_20666_, _20665_, _20574_);
  and (_43630_, _20666_, _43100_);
  and (_20667_, _11371_, \oc8051_golden_model_1.DPL [3]);
  or (_20668_, _20667_, _08140_);
  and (_20669_, _07849_, _08712_);
  or (_20670_, _20669_, _20667_);
  and (_20671_, _20670_, _06306_);
  and (_20672_, _20671_, _20668_);
  and (_20674_, _14738_, _07849_);
  or (_20675_, _20674_, _20667_);
  or (_20676_, _20675_, _06161_);
  and (_20677_, _07849_, \oc8051_golden_model_1.ACC [3]);
  or (_20678_, _20677_, _20667_);
  and (_20679_, _20678_, _07056_);
  and (_20680_, _07057_, \oc8051_golden_model_1.DPL [3]);
  or (_20681_, _20680_, _06160_);
  or (_20682_, _20681_, _20679_);
  and (_20683_, _20682_, _07075_);
  and (_20685_, _20683_, _20676_);
  and (_20686_, _07849_, _07544_);
  or (_20687_, _20686_, _20667_);
  and (_20688_, _20687_, _06217_);
  or (_20689_, _20688_, _06220_);
  or (_20690_, _20689_, _20685_);
  or (_20691_, _20678_, _06229_);
  and (_20692_, _20691_, _11312_);
  and (_20693_, _20692_, _20690_);
  nor (_20694_, _11317_, \oc8051_golden_model_1.DPL [3]);
  nor (_20696_, _20694_, _11318_);
  and (_20697_, _20696_, _11311_);
  or (_20698_, _20697_, _20693_);
  and (_20699_, _20698_, _11296_);
  nor (_20700_, _06389_, _11296_);
  or (_20701_, _20700_, _09842_);
  or (_20702_, _20701_, _20699_);
  or (_20703_, _20687_, _06132_);
  and (_20704_, _20703_, _20702_);
  or (_20705_, _20704_, _06116_);
  and (_20707_, _09210_, _07849_);
  or (_20708_, _20667_, _06117_);
  or (_20709_, _20708_, _20707_);
  and (_20710_, _20709_, _06114_);
  and (_20711_, _20710_, _20705_);
  and (_20712_, _14825_, _07849_);
  or (_20713_, _20712_, _20667_);
  and (_20714_, _20713_, _05787_);
  or (_20715_, _20714_, _11136_);
  or (_20716_, _20715_, _20711_);
  and (_20718_, _14727_, _07849_);
  or (_20719_, _20667_, _07127_);
  or (_20720_, _20719_, _20718_);
  or (_20721_, _20670_, _06111_);
  and (_20722_, _20721_, _07125_);
  and (_20723_, _20722_, _20720_);
  and (_20724_, _20723_, _20716_);
  and (_20725_, _12318_, _07849_);
  or (_20726_, _20725_, _20667_);
  and (_20727_, _20726_, _06402_);
  or (_20729_, _20727_, _20724_);
  and (_20730_, _20729_, _07132_);
  or (_20731_, _20730_, _20672_);
  and (_20732_, _20731_, _07130_);
  and (_20733_, _20678_, _06411_);
  and (_20734_, _20733_, _20668_);
  or (_20735_, _20734_, _06303_);
  or (_20736_, _20735_, _20732_);
  and (_20737_, _14724_, _07849_);
  or (_20738_, _20667_, _08819_);
  or (_20740_, _20738_, _20737_);
  and (_20741_, _20740_, _08824_);
  and (_20742_, _20741_, _20736_);
  nor (_20743_, _10273_, _11371_);
  or (_20744_, _20743_, _20667_);
  and (_20745_, _20744_, _06396_);
  or (_20746_, _20745_, _06433_);
  or (_20747_, _20746_, _20742_);
  or (_20748_, _20675_, _06829_);
  and (_20749_, _20748_, _06444_);
  and (_20751_, _20749_, _20747_);
  and (_20752_, _14897_, _07849_);
  or (_20753_, _20752_, _20667_);
  and (_20754_, _20753_, _06440_);
  or (_20755_, _20754_, _01321_);
  or (_20756_, _20755_, _20751_);
  or (_20757_, _01317_, \oc8051_golden_model_1.DPL [3]);
  and (_20758_, _20757_, _43100_);
  and (_43631_, _20758_, _20756_);
  and (_20759_, _11371_, \oc8051_golden_model_1.DPL [4]);
  and (_20760_, _08336_, _07849_);
  or (_20761_, _20760_, _20759_);
  or (_20762_, _20761_, _06132_);
  and (_20763_, _14928_, _07849_);
  or (_20764_, _20763_, _20759_);
  or (_20765_, _20764_, _06161_);
  and (_20766_, _07849_, \oc8051_golden_model_1.ACC [4]);
  or (_20767_, _20766_, _20759_);
  and (_20768_, _20767_, _07056_);
  and (_20769_, _07057_, \oc8051_golden_model_1.DPL [4]);
  or (_20771_, _20769_, _06160_);
  or (_20772_, _20771_, _20768_);
  and (_20773_, _20772_, _07075_);
  and (_20774_, _20773_, _20765_);
  and (_20775_, _20761_, _06217_);
  or (_20776_, _20775_, _06220_);
  or (_20777_, _20776_, _20774_);
  or (_20778_, _20767_, _06229_);
  and (_20779_, _20778_, _11312_);
  and (_20780_, _20779_, _20777_);
  nor (_20783_, _11318_, \oc8051_golden_model_1.DPL [4]);
  nor (_20784_, _20783_, _11319_);
  and (_20785_, _20784_, _11311_);
  or (_20786_, _20785_, _20780_);
  and (_20787_, _20786_, _11296_);
  nor (_20788_, _08670_, _11296_);
  or (_20789_, _20788_, _09842_);
  or (_20790_, _20789_, _20787_);
  and (_20791_, _20790_, _20762_);
  or (_20792_, _20791_, _06116_);
  and (_20794_, _09209_, _07849_);
  or (_20795_, _20759_, _06117_);
  or (_20796_, _20795_, _20794_);
  and (_20797_, _20796_, _06114_);
  and (_20798_, _20797_, _20792_);
  and (_20799_, _15013_, _07849_);
  or (_20800_, _20799_, _20759_);
  and (_20801_, _20800_, _05787_);
  or (_20802_, _20801_, _20798_);
  or (_20803_, _20802_, _11136_);
  and (_20804_, _15029_, _07849_);
  or (_20805_, _20759_, _07127_);
  or (_20806_, _20805_, _20804_);
  and (_20807_, _08715_, _07849_);
  or (_20808_, _20807_, _20759_);
  or (_20809_, _20808_, _06111_);
  and (_20810_, _20809_, _07125_);
  and (_20811_, _20810_, _20806_);
  and (_20812_, _20811_, _20803_);
  and (_20813_, _10289_, _07849_);
  or (_20815_, _20813_, _20759_);
  and (_20816_, _20815_, _06402_);
  or (_20817_, _20816_, _20812_);
  and (_20818_, _20817_, _07132_);
  or (_20819_, _20759_, _08339_);
  and (_20820_, _20808_, _06306_);
  and (_20821_, _20820_, _20819_);
  or (_20822_, _20821_, _20818_);
  and (_20823_, _20822_, _07130_);
  and (_20824_, _20767_, _06411_);
  and (_20827_, _20824_, _20819_);
  or (_20828_, _20827_, _06303_);
  or (_20829_, _20828_, _20823_);
  and (_20830_, _15026_, _07849_);
  or (_20831_, _20759_, _08819_);
  or (_20832_, _20831_, _20830_);
  and (_20833_, _20832_, _08824_);
  and (_20834_, _20833_, _20829_);
  nor (_20835_, _10288_, _11371_);
  or (_20836_, _20835_, _20759_);
  and (_20837_, _20836_, _06396_);
  or (_20838_, _20837_, _06433_);
  or (_20839_, _20838_, _20834_);
  or (_20840_, _20764_, _06829_);
  and (_20841_, _20840_, _06444_);
  and (_20842_, _20841_, _20839_);
  and (_20843_, _15087_, _07849_);
  or (_20844_, _20843_, _20759_);
  and (_20845_, _20844_, _06440_);
  or (_20846_, _20845_, _01321_);
  or (_20848_, _20846_, _20842_);
  or (_20849_, _01317_, \oc8051_golden_model_1.DPL [4]);
  and (_20850_, _20849_, _43100_);
  and (_43632_, _20850_, _20848_);
  and (_20851_, _11371_, \oc8051_golden_model_1.DPL [5]);
  and (_20852_, _08101_, _07849_);
  or (_20853_, _20852_, _20851_);
  or (_20854_, _20853_, _06132_);
  and (_20855_, _15119_, _07849_);
  or (_20856_, _20855_, _20851_);
  or (_20859_, _20856_, _06161_);
  and (_20860_, _07849_, \oc8051_golden_model_1.ACC [5]);
  or (_20861_, _20860_, _20851_);
  and (_20862_, _20861_, _07056_);
  and (_20863_, _07057_, \oc8051_golden_model_1.DPL [5]);
  or (_20864_, _20863_, _06160_);
  or (_20865_, _20864_, _20862_);
  and (_20866_, _20865_, _07075_);
  and (_20867_, _20866_, _20859_);
  and (_20868_, _20853_, _06217_);
  or (_20870_, _20868_, _06220_);
  or (_20871_, _20870_, _20867_);
  or (_20872_, _20861_, _06229_);
  and (_20873_, _20872_, _11312_);
  and (_20874_, _20873_, _20871_);
  nor (_20875_, _11319_, \oc8051_golden_model_1.DPL [5]);
  nor (_20876_, _20875_, _11320_);
  and (_20877_, _20876_, _11311_);
  or (_20878_, _20877_, _20874_);
  and (_20879_, _20878_, _11296_);
  nor (_20881_, _08701_, _11296_);
  or (_20882_, _20881_, _09842_);
  or (_20883_, _20882_, _20879_);
  and (_20884_, _20883_, _20854_);
  or (_20885_, _20884_, _06116_);
  and (_20886_, _09208_, _07849_);
  or (_20887_, _20851_, _06117_);
  or (_20888_, _20887_, _20886_);
  and (_20889_, _20888_, _06114_);
  and (_20890_, _20889_, _20885_);
  and (_20892_, _15203_, _07849_);
  or (_20893_, _20892_, _20851_);
  and (_20894_, _20893_, _05787_);
  or (_20895_, _20894_, _20890_);
  or (_20896_, _20895_, _11136_);
  and (_20897_, _15219_, _07849_);
  or (_20898_, _20851_, _07127_);
  or (_20899_, _20898_, _20897_);
  and (_20900_, _08736_, _07849_);
  or (_20901_, _20900_, _20851_);
  or (_20902_, _20901_, _06111_);
  and (_20903_, _20902_, _07125_);
  and (_20904_, _20903_, _20899_);
  and (_20905_, _20904_, _20896_);
  and (_20906_, _12325_, _07849_);
  or (_20907_, _20906_, _20851_);
  and (_20908_, _20907_, _06402_);
  or (_20909_, _20908_, _20905_);
  and (_20910_, _20909_, _07132_);
  or (_20911_, _20851_, _08104_);
  and (_20914_, _20901_, _06306_);
  and (_20915_, _20914_, _20911_);
  or (_20916_, _20915_, _20910_);
  and (_20917_, _20916_, _07130_);
  and (_20918_, _20861_, _06411_);
  and (_20919_, _20918_, _20911_);
  or (_20920_, _20919_, _06303_);
  or (_20921_, _20920_, _20917_);
  and (_20922_, _15216_, _07849_);
  or (_20923_, _20851_, _08819_);
  or (_20925_, _20923_, _20922_);
  and (_20926_, _20925_, _08824_);
  and (_20927_, _20926_, _20921_);
  nor (_20928_, _10269_, _11371_);
  or (_20929_, _20928_, _20851_);
  and (_20930_, _20929_, _06396_);
  or (_20931_, _20930_, _06433_);
  or (_20932_, _20931_, _20927_);
  or (_20933_, _20856_, _06829_);
  and (_20934_, _20933_, _06444_);
  and (_20936_, _20934_, _20932_);
  and (_20937_, _15275_, _07849_);
  or (_20938_, _20937_, _20851_);
  and (_20939_, _20938_, _06440_);
  or (_20940_, _20939_, _01321_);
  or (_20941_, _20940_, _20936_);
  or (_20942_, _01317_, \oc8051_golden_model_1.DPL [5]);
  and (_20943_, _20942_, _43100_);
  and (_43633_, _20943_, _20941_);
  and (_20944_, _11371_, \oc8051_golden_model_1.DPL [6]);
  and (_20946_, _08012_, _07849_);
  or (_20947_, _20946_, _20944_);
  or (_20948_, _20947_, _06132_);
  and (_20949_, _15300_, _07849_);
  or (_20950_, _20949_, _20944_);
  or (_20951_, _20950_, _06161_);
  and (_20952_, _07849_, \oc8051_golden_model_1.ACC [6]);
  or (_20953_, _20952_, _20944_);
  and (_20954_, _20953_, _07056_);
  and (_20955_, _07057_, \oc8051_golden_model_1.DPL [6]);
  or (_20957_, _20955_, _06160_);
  or (_20958_, _20957_, _20954_);
  and (_20959_, _20958_, _07075_);
  and (_20960_, _20959_, _20951_);
  and (_20961_, _20947_, _06217_);
  or (_20962_, _20961_, _06220_);
  or (_20963_, _20962_, _20960_);
  or (_20964_, _20953_, _06229_);
  and (_20965_, _20964_, _11312_);
  and (_20966_, _20965_, _20963_);
  nor (_20968_, _11320_, \oc8051_golden_model_1.DPL [6]);
  nor (_20969_, _20968_, _11321_);
  and (_20970_, _20969_, _11311_);
  or (_20971_, _20970_, _20966_);
  and (_20972_, _20971_, _11296_);
  nor (_20973_, _08638_, _11296_);
  or (_20974_, _20973_, _09842_);
  or (_20975_, _20974_, _20972_);
  and (_20976_, _20975_, _20948_);
  or (_20977_, _20976_, _06116_);
  and (_20979_, _09207_, _07849_);
  or (_20980_, _20944_, _06117_);
  or (_20981_, _20980_, _20979_);
  and (_20982_, _20981_, _06114_);
  and (_20983_, _20982_, _20977_);
  and (_20984_, _15395_, _07849_);
  or (_20985_, _20984_, _20944_);
  and (_20986_, _20985_, _05787_);
  or (_20987_, _20986_, _20983_);
  or (_20988_, _20987_, _11136_);
  and (_20990_, _15413_, _07849_);
  or (_20991_, _20944_, _07127_);
  or (_20992_, _20991_, _20990_);
  and (_20993_, _15402_, _07849_);
  or (_20994_, _20993_, _20944_);
  or (_20995_, _20994_, _06111_);
  and (_20996_, _20995_, _07125_);
  and (_20997_, _20996_, _20992_);
  and (_20998_, _20997_, _20988_);
  and (_20999_, _10295_, _07849_);
  or (_21001_, _20999_, _20944_);
  and (_21002_, _21001_, _06402_);
  or (_21003_, _21002_, _20998_);
  and (_21004_, _21003_, _07132_);
  or (_21005_, _20944_, _08015_);
  and (_21006_, _20994_, _06306_);
  and (_21007_, _21006_, _21005_);
  or (_21008_, _21007_, _21004_);
  and (_21009_, _21008_, _07130_);
  and (_21010_, _20953_, _06411_);
  and (_21012_, _21010_, _21005_);
  or (_21013_, _21012_, _06303_);
  or (_21014_, _21013_, _21009_);
  and (_21015_, _15410_, _07849_);
  or (_21016_, _20944_, _08819_);
  or (_21017_, _21016_, _21015_);
  and (_21018_, _21017_, _08824_);
  and (_21019_, _21018_, _21014_);
  nor (_21020_, _10294_, _11371_);
  or (_21021_, _21020_, _20944_);
  and (_21023_, _21021_, _06396_);
  or (_21024_, _21023_, _06433_);
  or (_21025_, _21024_, _21019_);
  or (_21026_, _20950_, _06829_);
  and (_21027_, _21026_, _06444_);
  and (_21028_, _21027_, _21025_);
  and (_21029_, _15478_, _07849_);
  or (_21030_, _21029_, _20944_);
  and (_21031_, _21030_, _06440_);
  or (_21032_, _21031_, _01321_);
  or (_21033_, _21032_, _21028_);
  or (_21034_, _01317_, \oc8051_golden_model_1.DPL [6]);
  and (_21035_, _21034_, _43100_);
  and (_43634_, _21035_, _21033_);
  nor (_21036_, _01317_, _12434_);
  nor (_21037_, _11390_, _12434_);
  and (_21038_, _11390_, \oc8051_golden_model_1.ACC [0]);
  and (_21039_, _21038_, _08211_);
  or (_21040_, _21039_, _21037_);
  or (_21041_, _21040_, _07130_);
  nor (_21044_, _08211_, _11468_);
  or (_21045_, _21044_, _21037_);
  or (_21046_, _21045_, _06161_);
  or (_21047_, _21038_, _21037_);
  and (_21048_, _21047_, _07056_);
  nor (_21049_, _07056_, _12434_);
  or (_21050_, _21049_, _06160_);
  or (_21051_, _21050_, _21048_);
  and (_21052_, _21051_, _07075_);
  and (_21053_, _21052_, _21046_);
  and (_21055_, _07852_, _07049_);
  or (_21056_, _21055_, _21037_);
  and (_21057_, _21056_, _06217_);
  or (_21058_, _21057_, _06220_);
  or (_21059_, _21058_, _21053_);
  or (_21060_, _21047_, _06229_);
  and (_21061_, _21060_, _11312_);
  and (_21062_, _21061_, _21059_);
  nor (_21063_, _11323_, \oc8051_golden_model_1.DPH [0]);
  nor (_21064_, _21063_, _11412_);
  and (_21066_, _21064_, _11311_);
  or (_21067_, _21066_, _21062_);
  and (_21068_, _21067_, _11296_);
  nor (_21069_, _11296_, _06107_);
  or (_21070_, _21069_, _09842_);
  or (_21071_, _21070_, _21068_);
  or (_21072_, _21056_, _06132_);
  and (_21073_, _21072_, _21071_);
  or (_21074_, _21073_, _06116_);
  and (_21075_, _09160_, _11390_);
  or (_21077_, _21037_, _06117_);
  or (_21078_, _21077_, _21075_);
  and (_21079_, _21078_, _21074_);
  or (_21080_, _21079_, _05787_);
  and (_21081_, _14260_, _11390_);
  or (_21082_, _21081_, _21037_);
  or (_21083_, _21082_, _06114_);
  and (_21084_, _21083_, _06111_);
  and (_21085_, _21084_, _21080_);
  and (_21086_, _11390_, _08708_);
  or (_21088_, _21086_, _21037_);
  and (_21089_, _21088_, _06110_);
  or (_21090_, _21089_, _06297_);
  or (_21091_, _21090_, _21085_);
  and (_21092_, _14275_, _07852_);
  or (_21093_, _21037_, _07127_);
  or (_21094_, _21093_, _21092_);
  and (_21095_, _21094_, _07125_);
  and (_21096_, _21095_, _21091_);
  nor (_21097_, _12321_, _11468_);
  or (_21099_, _21097_, _21037_);
  nor (_21100_, _21039_, _07125_);
  and (_21101_, _21100_, _21099_);
  or (_21102_, _21101_, _21096_);
  and (_21103_, _21102_, _07132_);
  nand (_21104_, _21088_, _06306_);
  nor (_21105_, _21104_, _21044_);
  or (_21106_, _21105_, _06411_);
  or (_21107_, _21106_, _21103_);
  and (_21108_, _21107_, _21041_);
  or (_21110_, _21108_, _06303_);
  and (_21111_, _14167_, _07852_);
  or (_21112_, _21037_, _08819_);
  or (_21113_, _21112_, _21111_);
  and (_21114_, _21113_, _08824_);
  and (_21115_, _21114_, _21110_);
  and (_21116_, _21099_, _06396_);
  or (_21117_, _21116_, _19287_);
  or (_21118_, _21117_, _21115_);
  or (_21119_, _21045_, _06630_);
  and (_21121_, _21119_, _01317_);
  and (_21122_, _21121_, _21118_);
  or (_21123_, _21122_, _21036_);
  and (_43636_, _21123_, _43100_);
  not (_21124_, \oc8051_golden_model_1.DPH [1]);
  nor (_21125_, _11390_, _21124_);
  nor (_21126_, _10277_, _11468_);
  or (_21127_, _21126_, _21125_);
  or (_21128_, _21127_, _08824_);
  or (_21129_, _14442_, _11468_);
  or (_21131_, _11390_, \oc8051_golden_model_1.DPH [1]);
  and (_21132_, _21131_, _05787_);
  and (_21133_, _21132_, _21129_);
  and (_21134_, _09115_, _11390_);
  or (_21135_, _21134_, _21125_);
  and (_21136_, _21135_, _06116_);
  and (_21137_, _14363_, _07852_);
  not (_21138_, _21137_);
  and (_21139_, _21138_, _21131_);
  or (_21140_, _21139_, _06161_);
  and (_21142_, _11390_, \oc8051_golden_model_1.ACC [1]);
  or (_21143_, _21142_, _21125_);
  and (_21144_, _21143_, _07056_);
  nor (_21145_, _07056_, _21124_);
  or (_21146_, _21145_, _06160_);
  or (_21147_, _21146_, _21144_);
  and (_21148_, _21147_, _07075_);
  and (_21149_, _21148_, _21140_);
  and (_21150_, _07852_, _07306_);
  or (_21151_, _21150_, _21125_);
  and (_21153_, _21151_, _06217_);
  or (_21154_, _21153_, _06220_);
  or (_21155_, _21154_, _21149_);
  or (_21156_, _21143_, _06229_);
  and (_21157_, _21156_, _11312_);
  and (_21158_, _21157_, _21155_);
  nor (_21159_, _11412_, \oc8051_golden_model_1.DPH [1]);
  nor (_21160_, _21159_, _11413_);
  and (_21161_, _21160_, _11311_);
  or (_21162_, _21161_, _21158_);
  and (_21164_, _21162_, _11296_);
  nor (_21165_, _06912_, _11296_);
  or (_21166_, _21165_, _09842_);
  or (_21167_, _21166_, _21164_);
  or (_21168_, _21151_, _06132_);
  and (_21169_, _21168_, _06117_);
  and (_21170_, _21169_, _21167_);
  or (_21171_, _21170_, _21136_);
  and (_21172_, _21171_, _06114_);
  or (_21173_, _21172_, _21133_);
  and (_21175_, _21173_, _06298_);
  or (_21176_, _14346_, _11468_);
  and (_21177_, _21176_, _06297_);
  nand (_21178_, _07852_, _06945_);
  and (_21179_, _21178_, _06110_);
  or (_21180_, _21179_, _21177_);
  and (_21181_, _21180_, _21131_);
  or (_21182_, _21181_, _06402_);
  or (_21183_, _21182_, _21175_);
  nand (_21184_, _10275_, _07852_);
  and (_21186_, _21184_, _21127_);
  or (_21187_, _21186_, _07125_);
  and (_21188_, _21187_, _07132_);
  and (_21189_, _21188_, _21183_);
  or (_21190_, _14344_, _11468_);
  and (_21191_, _21131_, _06306_);
  and (_21192_, _21191_, _21190_);
  or (_21193_, _21192_, _06411_);
  or (_21194_, _21193_, _21189_);
  nor (_21195_, _21125_, _07130_);
  nand (_21197_, _21195_, _21184_);
  and (_21198_, _21197_, _08819_);
  and (_21199_, _21198_, _21194_);
  or (_21200_, _21178_, _08176_);
  and (_21201_, _21131_, _06303_);
  and (_21202_, _21201_, _21200_);
  or (_21203_, _21202_, _06396_);
  or (_21204_, _21203_, _21199_);
  and (_21205_, _21204_, _21128_);
  or (_21206_, _21205_, _06433_);
  or (_21207_, _21139_, _06829_);
  and (_21208_, _21207_, _06444_);
  and (_21209_, _21208_, _21206_);
  or (_21210_, _21137_, _21125_);
  and (_21211_, _21210_, _06440_);
  or (_21212_, _21211_, _01321_);
  or (_21213_, _21212_, _21209_);
  or (_21214_, _01317_, \oc8051_golden_model_1.DPH [1]);
  and (_21215_, _21214_, _43100_);
  and (_43637_, _21215_, _21213_);
  and (_21218_, _01321_, \oc8051_golden_model_1.DPH [2]);
  and (_21219_, _11468_, \oc8051_golden_model_1.DPH [2]);
  and (_21220_, _07852_, _07708_);
  or (_21221_, _21220_, _21219_);
  or (_21222_, _21221_, _06132_);
  and (_21223_, _14542_, _07852_);
  or (_21224_, _21223_, _21219_);
  or (_21225_, _21224_, _06161_);
  and (_21226_, _11390_, \oc8051_golden_model_1.ACC [2]);
  or (_21227_, _21226_, _21219_);
  and (_21229_, _21227_, _07056_);
  and (_21230_, _07057_, \oc8051_golden_model_1.DPH [2]);
  or (_21231_, _21230_, _06160_);
  or (_21232_, _21231_, _21229_);
  and (_21233_, _21232_, _07075_);
  and (_21234_, _21233_, _21225_);
  and (_21235_, _21221_, _06217_);
  or (_21236_, _21235_, _06220_);
  or (_21237_, _21236_, _21234_);
  or (_21238_, _21227_, _06229_);
  and (_21240_, _21238_, _11312_);
  and (_21241_, _21240_, _21237_);
  or (_21242_, _11413_, \oc8051_golden_model_1.DPH [2]);
  nor (_21243_, _11414_, _11312_);
  and (_21244_, _21243_, _21242_);
  or (_21245_, _21244_, _21241_);
  and (_21246_, _21245_, _11296_);
  nor (_21247_, _06625_, _11296_);
  or (_21248_, _21247_, _09842_);
  or (_21249_, _21248_, _21246_);
  and (_21251_, _21249_, _21222_);
  or (_21252_, _21251_, _06116_);
  or (_21253_, _21219_, _06117_);
  and (_21254_, _09211_, _11390_);
  or (_21255_, _21254_, _21253_);
  and (_21256_, _21255_, _06114_);
  and (_21257_, _21256_, _21252_);
  and (_21258_, _14630_, _11390_);
  or (_21259_, _21258_, _21219_);
  and (_21260_, _21259_, _05787_);
  or (_21262_, _21260_, _21257_);
  or (_21263_, _21262_, _11136_);
  and (_21264_, _14646_, _07852_);
  or (_21265_, _21219_, _07127_);
  or (_21266_, _21265_, _21264_);
  and (_21267_, _11390_, _08768_);
  or (_21268_, _21267_, _21219_);
  or (_21269_, _21268_, _06111_);
  and (_21270_, _21269_, _07125_);
  and (_21271_, _21270_, _21266_);
  and (_21273_, _21271_, _21263_);
  and (_21274_, _10282_, _11390_);
  or (_21275_, _21274_, _21219_);
  and (_21276_, _21275_, _06402_);
  or (_21277_, _21276_, _21273_);
  and (_21278_, _21277_, _07132_);
  or (_21279_, _21219_, _08248_);
  and (_21280_, _21268_, _06306_);
  and (_21281_, _21280_, _21279_);
  or (_21282_, _21281_, _21278_);
  and (_21284_, _21282_, _07130_);
  and (_21285_, _21227_, _06411_);
  and (_21286_, _21285_, _21279_);
  or (_21287_, _21286_, _06303_);
  or (_21288_, _21287_, _21284_);
  and (_21289_, _14643_, _07852_);
  or (_21290_, _21219_, _08819_);
  or (_21291_, _21290_, _21289_);
  and (_21292_, _21291_, _08824_);
  and (_21293_, _21292_, _21288_);
  nor (_21295_, _10281_, _11468_);
  or (_21296_, _21295_, _21219_);
  and (_21297_, _21296_, _06396_);
  or (_21298_, _21297_, _21293_);
  and (_21299_, _21298_, _06829_);
  and (_21300_, _21224_, _06433_);
  or (_21301_, _21300_, _06440_);
  or (_21302_, _21301_, _21299_);
  and (_21303_, _14710_, _07852_);
  or (_21304_, _21219_, _06444_);
  or (_21306_, _21304_, _21303_);
  and (_21307_, _21306_, _01317_);
  and (_21308_, _21307_, _21302_);
  or (_21309_, _21308_, _21218_);
  and (_43638_, _21309_, _43100_);
  and (_21310_, _11468_, \oc8051_golden_model_1.DPH [3]);
  or (_21311_, _21310_, _08140_);
  and (_21312_, _11390_, _08712_);
  or (_21313_, _21312_, _21310_);
  and (_21314_, _21313_, _06306_);
  and (_21316_, _21314_, _21311_);
  and (_21317_, _14738_, _07852_);
  or (_21318_, _21317_, _21310_);
  or (_21319_, _21318_, _06161_);
  and (_21320_, _11390_, \oc8051_golden_model_1.ACC [3]);
  or (_21321_, _21320_, _21310_);
  and (_21322_, _21321_, _07056_);
  and (_21323_, _07057_, \oc8051_golden_model_1.DPH [3]);
  or (_21324_, _21323_, _06160_);
  or (_21325_, _21324_, _21322_);
  and (_21327_, _21325_, _07075_);
  and (_21328_, _21327_, _21319_);
  and (_21329_, _07852_, _07544_);
  or (_21330_, _21329_, _21310_);
  and (_21331_, _21330_, _06217_);
  or (_21332_, _21331_, _06220_);
  or (_21333_, _21332_, _21328_);
  or (_21334_, _21321_, _06229_);
  and (_21335_, _21334_, _11312_);
  and (_21336_, _21335_, _21333_);
  or (_21338_, _11414_, \oc8051_golden_model_1.DPH [3]);
  nor (_21339_, _11415_, _11312_);
  and (_21340_, _21339_, _21338_);
  or (_21341_, _21340_, _21336_);
  and (_21342_, _21341_, _11296_);
  nor (_21343_, _11296_, _06070_);
  or (_21344_, _21343_, _09842_);
  or (_21345_, _21344_, _21342_);
  or (_21346_, _21330_, _06132_);
  and (_21347_, _21346_, _21345_);
  or (_21349_, _21347_, _06116_);
  and (_21350_, _09210_, _11390_);
  or (_21351_, _21310_, _06117_);
  or (_21352_, _21351_, _21350_);
  and (_21353_, _21352_, _06114_);
  and (_21354_, _21353_, _21349_);
  and (_21355_, _14825_, _07852_);
  or (_21356_, _21355_, _21310_);
  and (_21357_, _21356_, _05787_);
  or (_21358_, _21357_, _11136_);
  or (_21360_, _21358_, _21354_);
  and (_21361_, _14727_, _07852_);
  or (_21362_, _21310_, _07127_);
  or (_21363_, _21362_, _21361_);
  or (_21364_, _21313_, _06111_);
  and (_21365_, _21364_, _07125_);
  and (_21366_, _21365_, _21363_);
  and (_21367_, _21366_, _21360_);
  and (_21368_, _12318_, _11390_);
  or (_21369_, _21368_, _21310_);
  and (_21371_, _21369_, _06402_);
  or (_21372_, _21371_, _21367_);
  and (_21373_, _21372_, _07132_);
  or (_21374_, _21373_, _21316_);
  and (_21375_, _21374_, _07130_);
  and (_21376_, _21321_, _06411_);
  and (_21377_, _21376_, _21311_);
  or (_21378_, _21377_, _06303_);
  or (_21379_, _21378_, _21375_);
  and (_21380_, _14724_, _07852_);
  or (_21382_, _21310_, _08819_);
  or (_21383_, _21382_, _21380_);
  and (_21384_, _21383_, _08824_);
  and (_21385_, _21384_, _21379_);
  nor (_21386_, _10273_, _11468_);
  or (_21387_, _21386_, _21310_);
  and (_21388_, _21387_, _06396_);
  or (_21389_, _21388_, _06433_);
  or (_21390_, _21389_, _21385_);
  or (_21391_, _21318_, _06829_);
  and (_21393_, _21391_, _06444_);
  and (_21394_, _21393_, _21390_);
  and (_21395_, _14897_, _07852_);
  or (_21396_, _21395_, _21310_);
  and (_21397_, _21396_, _06440_);
  or (_21398_, _21397_, _01321_);
  or (_21399_, _21398_, _21394_);
  or (_21400_, _01317_, \oc8051_golden_model_1.DPH [3]);
  and (_21401_, _21400_, _43100_);
  and (_43640_, _21401_, _21399_);
  not (_21402_, \oc8051_golden_model_1.DPH [4]);
  nor (_21403_, _11390_, _21402_);
  and (_21404_, _08336_, _07852_);
  or (_21405_, _21404_, _21403_);
  or (_21406_, _21405_, _06132_);
  and (_21407_, _14928_, _07852_);
  or (_21408_, _21407_, _21403_);
  or (_21409_, _21408_, _06161_);
  and (_21410_, _11390_, \oc8051_golden_model_1.ACC [4]);
  or (_21411_, _21410_, _21403_);
  and (_21414_, _21411_, _07056_);
  nor (_21415_, _07056_, _21402_);
  or (_21416_, _21415_, _06160_);
  or (_21417_, _21416_, _21414_);
  and (_21418_, _21417_, _07075_);
  and (_21419_, _21418_, _21409_);
  and (_21420_, _21405_, _06217_);
  or (_21421_, _21420_, _06220_);
  or (_21422_, _21421_, _21419_);
  or (_21423_, _21411_, _06229_);
  and (_21425_, _21423_, _11312_);
  and (_21426_, _21425_, _21422_);
  or (_21427_, _11415_, \oc8051_golden_model_1.DPH [4]);
  nor (_21428_, _11416_, _11312_);
  and (_21429_, _21428_, _21427_);
  or (_21430_, _21429_, _21426_);
  and (_21431_, _21430_, _11296_);
  nor (_21432_, _06876_, _11296_);
  or (_21433_, _21432_, _09842_);
  or (_21434_, _21433_, _21431_);
  and (_21436_, _21434_, _21406_);
  or (_21437_, _21436_, _06116_);
  or (_21438_, _21403_, _06117_);
  and (_21439_, _09209_, _11390_);
  or (_21440_, _21439_, _21438_);
  and (_21441_, _21440_, _06114_);
  and (_21442_, _21441_, _21437_);
  and (_21443_, _15013_, _11390_);
  or (_21444_, _21443_, _21403_);
  and (_21445_, _21444_, _05787_);
  or (_21447_, _21445_, _21442_);
  or (_21448_, _21447_, _11136_);
  and (_21449_, _15029_, _07852_);
  or (_21450_, _21403_, _07127_);
  or (_21451_, _21450_, _21449_);
  and (_21452_, _08715_, _11390_);
  or (_21453_, _21452_, _21403_);
  or (_21454_, _21453_, _06111_);
  and (_21455_, _21454_, _07125_);
  and (_21456_, _21455_, _21451_);
  and (_21458_, _21456_, _21448_);
  and (_21459_, _10289_, _11390_);
  or (_21460_, _21459_, _21403_);
  and (_21461_, _21460_, _06402_);
  or (_21462_, _21461_, _21458_);
  and (_21463_, _21462_, _07132_);
  or (_21464_, _21403_, _08339_);
  and (_21465_, _21453_, _06306_);
  and (_21466_, _21465_, _21464_);
  or (_21467_, _21466_, _21463_);
  and (_21469_, _21467_, _07130_);
  and (_21470_, _21411_, _06411_);
  and (_21471_, _21470_, _21464_);
  or (_21472_, _21471_, _06303_);
  or (_21473_, _21472_, _21469_);
  and (_21474_, _15026_, _07852_);
  or (_21475_, _21403_, _08819_);
  or (_21476_, _21475_, _21474_);
  and (_21477_, _21476_, _08824_);
  and (_21478_, _21477_, _21473_);
  nor (_21480_, _10288_, _11468_);
  or (_21481_, _21480_, _21403_);
  and (_21482_, _21481_, _06396_);
  or (_21483_, _21482_, _06433_);
  or (_21484_, _21483_, _21478_);
  or (_21485_, _21408_, _06829_);
  and (_21486_, _21485_, _06444_);
  and (_21487_, _21486_, _21484_);
  and (_21488_, _15087_, _07852_);
  or (_21489_, _21488_, _21403_);
  and (_21491_, _21489_, _06440_);
  or (_21492_, _21491_, _01321_);
  or (_21493_, _21492_, _21487_);
  or (_21494_, _01317_, \oc8051_golden_model_1.DPH [4]);
  and (_21495_, _21494_, _43100_);
  and (_43641_, _21495_, _21493_);
  and (_21496_, _11468_, \oc8051_golden_model_1.DPH [5]);
  and (_21497_, _08101_, _07852_);
  or (_21498_, _21497_, _21496_);
  or (_21499_, _21498_, _06132_);
  and (_21501_, _15119_, _07852_);
  or (_21502_, _21501_, _21496_);
  or (_21503_, _21502_, _06161_);
  and (_21504_, _11390_, \oc8051_golden_model_1.ACC [5]);
  or (_21505_, _21504_, _21496_);
  and (_21506_, _21505_, _07056_);
  and (_21507_, _07057_, \oc8051_golden_model_1.DPH [5]);
  or (_21508_, _21507_, _06160_);
  or (_21509_, _21508_, _21506_);
  and (_21510_, _21509_, _07075_);
  and (_21512_, _21510_, _21503_);
  and (_21513_, _21498_, _06217_);
  or (_21514_, _21513_, _06220_);
  or (_21515_, _21514_, _21512_);
  or (_21516_, _21505_, _06229_);
  and (_21517_, _21516_, _11312_);
  and (_21518_, _21517_, _21515_);
  or (_21519_, _11416_, \oc8051_golden_model_1.DPH [5]);
  nor (_21520_, _11417_, _11312_);
  and (_21521_, _21520_, _21519_);
  or (_21523_, _21521_, _21518_);
  and (_21524_, _21523_, _11296_);
  nor (_21525_, _06477_, _11296_);
  or (_21526_, _21525_, _09842_);
  or (_21527_, _21526_, _21524_);
  and (_21528_, _21527_, _21499_);
  or (_21529_, _21528_, _06116_);
  or (_21530_, _21496_, _06117_);
  and (_21531_, _09208_, _11390_);
  or (_21532_, _21531_, _21530_);
  and (_21534_, _21532_, _06114_);
  and (_21535_, _21534_, _21529_);
  and (_21536_, _15203_, _11390_);
  or (_21537_, _21536_, _21496_);
  and (_21538_, _21537_, _05787_);
  or (_21539_, _21538_, _21535_);
  or (_21540_, _21539_, _11136_);
  and (_21541_, _15219_, _07852_);
  or (_21542_, _21496_, _07127_);
  or (_21543_, _21542_, _21541_);
  and (_21545_, _08736_, _11390_);
  or (_21546_, _21545_, _21496_);
  or (_21547_, _21546_, _06111_);
  and (_21548_, _21547_, _07125_);
  and (_21549_, _21548_, _21543_);
  and (_21550_, _21549_, _21540_);
  and (_21551_, _12325_, _11390_);
  or (_21552_, _21551_, _21496_);
  and (_21553_, _21552_, _06402_);
  or (_21554_, _21553_, _21550_);
  and (_21556_, _21554_, _07132_);
  or (_21557_, _21496_, _08104_);
  and (_21558_, _21546_, _06306_);
  and (_21559_, _21558_, _21557_);
  or (_21560_, _21559_, _21556_);
  and (_21561_, _21560_, _07130_);
  and (_21562_, _21505_, _06411_);
  and (_21563_, _21562_, _21557_);
  or (_21564_, _21563_, _06303_);
  or (_21565_, _21564_, _21561_);
  and (_21567_, _15216_, _07852_);
  or (_21568_, _21496_, _08819_);
  or (_21569_, _21568_, _21567_);
  and (_21570_, _21569_, _08824_);
  and (_21571_, _21570_, _21565_);
  nor (_21572_, _10269_, _11468_);
  or (_21573_, _21572_, _21496_);
  and (_21574_, _21573_, _06396_);
  or (_21575_, _21574_, _06433_);
  or (_21576_, _21575_, _21571_);
  or (_21578_, _21502_, _06829_);
  and (_21579_, _21578_, _06444_);
  and (_21580_, _21579_, _21576_);
  and (_21581_, _15275_, _07852_);
  or (_21582_, _21581_, _21496_);
  and (_21583_, _21582_, _06440_);
  or (_21584_, _21583_, _01321_);
  or (_21585_, _21584_, _21580_);
  or (_21586_, _01317_, \oc8051_golden_model_1.DPH [5]);
  and (_21587_, _21586_, _43100_);
  and (_43642_, _21587_, _21585_);
  not (_21589_, \oc8051_golden_model_1.DPH [6]);
  nor (_21590_, _11390_, _21589_);
  and (_21591_, _08012_, _07852_);
  or (_21592_, _21591_, _21590_);
  or (_21593_, _21592_, _06132_);
  and (_21594_, _15300_, _07852_);
  or (_21595_, _21594_, _21590_);
  or (_21596_, _21595_, _06161_);
  and (_21597_, _11390_, \oc8051_golden_model_1.ACC [6]);
  or (_21599_, _21597_, _21590_);
  and (_21600_, _21599_, _07056_);
  nor (_21601_, _07056_, _21589_);
  or (_21602_, _21601_, _06160_);
  or (_21603_, _21602_, _21600_);
  and (_21604_, _21603_, _07075_);
  and (_21605_, _21604_, _21596_);
  and (_21606_, _21592_, _06217_);
  or (_21607_, _21606_, _06220_);
  or (_21608_, _21607_, _21605_);
  or (_21610_, _21599_, _06229_);
  and (_21611_, _21610_, _11312_);
  and (_21612_, _21611_, _21608_);
  or (_21613_, _11417_, \oc8051_golden_model_1.DPH [6]);
  nor (_21614_, _11418_, _11312_);
  and (_21615_, _21614_, _21613_);
  or (_21616_, _21615_, _21612_);
  and (_21617_, _21616_, _11296_);
  nor (_21618_, _11296_, _06203_);
  or (_21619_, _21618_, _09842_);
  or (_21621_, _21619_, _21617_);
  and (_21622_, _21621_, _21593_);
  or (_21623_, _21622_, _06116_);
  or (_21624_, _21590_, _06117_);
  and (_21625_, _09207_, _11390_);
  or (_21626_, _21625_, _21624_);
  and (_21627_, _21626_, _06114_);
  and (_21628_, _21627_, _21623_);
  and (_21629_, _15395_, _11390_);
  or (_21630_, _21629_, _21590_);
  and (_21632_, _21630_, _05787_);
  or (_21633_, _21632_, _21628_);
  or (_21634_, _21633_, _11136_);
  and (_21635_, _15413_, _07852_);
  or (_21636_, _21590_, _07127_);
  or (_21637_, _21636_, _21635_);
  and (_21638_, _15402_, _11390_);
  or (_21639_, _21638_, _21590_);
  or (_21640_, _21639_, _06111_);
  and (_21641_, _21640_, _07125_);
  and (_21643_, _21641_, _21637_);
  and (_21644_, _21643_, _21634_);
  and (_21645_, _10295_, _11390_);
  or (_21646_, _21645_, _21590_);
  and (_21647_, _21646_, _06402_);
  or (_21648_, _21647_, _21644_);
  and (_21649_, _21648_, _07132_);
  or (_21650_, _21590_, _08015_);
  and (_21651_, _21639_, _06306_);
  and (_21652_, _21651_, _21650_);
  or (_21654_, _21652_, _21649_);
  and (_21655_, _21654_, _07130_);
  and (_21656_, _21599_, _06411_);
  and (_21657_, _21656_, _21650_);
  or (_21658_, _21657_, _06303_);
  or (_21659_, _21658_, _21655_);
  and (_21660_, _15410_, _07852_);
  or (_21661_, _21590_, _08819_);
  or (_21662_, _21661_, _21660_);
  and (_21663_, _21662_, _08824_);
  and (_21665_, _21663_, _21659_);
  nor (_21666_, _10294_, _11468_);
  or (_21667_, _21666_, _21590_);
  and (_21668_, _21667_, _06396_);
  or (_21669_, _21668_, _06433_);
  or (_21670_, _21669_, _21665_);
  or (_21671_, _21595_, _06829_);
  and (_21672_, _21671_, _06444_);
  and (_21673_, _21672_, _21670_);
  and (_21674_, _15478_, _07852_);
  or (_21676_, _21674_, _21590_);
  and (_21677_, _21676_, _06440_);
  or (_21678_, _21677_, _01321_);
  or (_21679_, _21678_, _21673_);
  or (_21680_, _01317_, \oc8051_golden_model_1.DPH [6]);
  and (_21681_, _21680_, _43100_);
  and (_43643_, _21681_, _21679_);
  not (_21682_, \oc8051_golden_model_1.TL1 [0]);
  nor (_21683_, _01317_, _21682_);
  nand (_21684_, _10276_, _07837_);
  nor (_21686_, _07837_, _21682_);
  nor (_21687_, _21686_, _07130_);
  nand (_21688_, _21687_, _21684_);
  nor (_21689_, _08211_, _11484_);
  or (_21690_, _21689_, _21686_);
  or (_21691_, _21690_, _06161_);
  and (_21692_, _07837_, \oc8051_golden_model_1.ACC [0]);
  or (_21693_, _21692_, _21686_);
  and (_21694_, _21693_, _07056_);
  nor (_21695_, _07056_, _21682_);
  or (_21697_, _21695_, _06160_);
  or (_21698_, _21697_, _21694_);
  and (_21699_, _21698_, _07075_);
  and (_21700_, _21699_, _21691_);
  and (_21701_, _07837_, _07049_);
  or (_21702_, _21701_, _21686_);
  and (_21703_, _21702_, _06217_);
  or (_21704_, _21703_, _21700_);
  and (_21705_, _21704_, _06229_);
  and (_21706_, _21693_, _06220_);
  or (_21708_, _21706_, _09842_);
  or (_21709_, _21708_, _21705_);
  or (_21710_, _21702_, _06132_);
  and (_21711_, _21710_, _21709_);
  or (_21712_, _21711_, _06116_);
  and (_21713_, _09160_, _07837_);
  or (_21714_, _21686_, _06117_);
  or (_21715_, _21714_, _21713_);
  and (_21716_, _21715_, _21712_);
  or (_21717_, _21716_, _05787_);
  and (_21719_, _14260_, _07837_);
  or (_21720_, _21686_, _06114_);
  or (_21721_, _21720_, _21719_);
  and (_21722_, _21721_, _06111_);
  and (_21723_, _21722_, _21717_);
  and (_21724_, _07837_, _08708_);
  or (_21725_, _21724_, _21686_);
  and (_21726_, _21725_, _06110_);
  or (_21727_, _21726_, _06297_);
  or (_21728_, _21727_, _21723_);
  and (_21730_, _14275_, _07837_);
  or (_21731_, _21730_, _21686_);
  or (_21732_, _21731_, _07127_);
  and (_21733_, _21732_, _07125_);
  and (_21734_, _21733_, _21728_);
  nor (_21735_, _12321_, _11484_);
  or (_21736_, _21735_, _21686_);
  and (_21737_, _21684_, _06402_);
  and (_21738_, _21737_, _21736_);
  or (_21739_, _21738_, _21734_);
  and (_21741_, _21739_, _07132_);
  nand (_21742_, _21725_, _06306_);
  nor (_21743_, _21742_, _21689_);
  or (_21744_, _21743_, _06411_);
  or (_21745_, _21744_, _21741_);
  and (_21746_, _21745_, _21688_);
  or (_21747_, _21746_, _06303_);
  and (_21748_, _14167_, _07837_);
  or (_21749_, _21686_, _08819_);
  or (_21750_, _21749_, _21748_);
  and (_21751_, _21750_, _08824_);
  and (_21752_, _21751_, _21747_);
  and (_21753_, _21736_, _06396_);
  or (_21754_, _21753_, _19287_);
  or (_21755_, _21754_, _21752_);
  or (_21756_, _21690_, _06630_);
  and (_21757_, _21756_, _01317_);
  and (_21758_, _21757_, _21755_);
  or (_21759_, _21758_, _21683_);
  and (_43645_, _21759_, _43100_);
  not (_21762_, \oc8051_golden_model_1.TL1 [1]);
  nor (_21763_, _01317_, _21762_);
  and (_21764_, _09115_, _07837_);
  nor (_21765_, _07837_, _21762_);
  or (_21766_, _21765_, _06117_);
  or (_21767_, _21766_, _21764_);
  and (_21768_, _07837_, _07306_);
  or (_21769_, _21768_, _21765_);
  or (_21770_, _21769_, _06132_);
  or (_21771_, _07837_, \oc8051_golden_model_1.TL1 [1]);
  and (_21773_, _14363_, _07837_);
  not (_21774_, _21773_);
  and (_21775_, _21774_, _21771_);
  or (_21776_, _21775_, _06161_);
  and (_21777_, _07837_, \oc8051_golden_model_1.ACC [1]);
  or (_21778_, _21777_, _21765_);
  and (_21779_, _21778_, _07056_);
  nor (_21780_, _07056_, _21762_);
  or (_21781_, _21780_, _06160_);
  or (_21782_, _21781_, _21779_);
  and (_21784_, _21782_, _07075_);
  and (_21785_, _21784_, _21776_);
  and (_21786_, _21769_, _06217_);
  or (_21787_, _21786_, _21785_);
  and (_21788_, _21787_, _06229_);
  and (_21789_, _21778_, _06220_);
  or (_21790_, _21789_, _09842_);
  or (_21791_, _21790_, _21788_);
  and (_21792_, _21791_, _21770_);
  or (_21793_, _21792_, _06116_);
  and (_21795_, _21793_, _06114_);
  and (_21796_, _21795_, _21767_);
  or (_21797_, _14442_, _11484_);
  and (_21798_, _21771_, _05787_);
  and (_21799_, _21798_, _21797_);
  or (_21800_, _21799_, _21796_);
  and (_21801_, _21800_, _06298_);
  or (_21802_, _14346_, _11484_);
  and (_21803_, _21802_, _06297_);
  nand (_21804_, _07837_, _06945_);
  and (_21806_, _21804_, _06110_);
  or (_21807_, _21806_, _21803_);
  and (_21808_, _21807_, _21771_);
  or (_21809_, _21808_, _06402_);
  or (_21810_, _21809_, _21801_);
  nor (_21811_, _10277_, _11484_);
  or (_21812_, _21811_, _21765_);
  nand (_21813_, _10275_, _07837_);
  and (_21814_, _21813_, _21812_);
  or (_21815_, _21814_, _07125_);
  and (_21817_, _21815_, _07132_);
  and (_21818_, _21817_, _21810_);
  or (_21819_, _14344_, _11484_);
  and (_21820_, _21771_, _06306_);
  and (_21821_, _21820_, _21819_);
  or (_21822_, _21821_, _06411_);
  or (_21823_, _21822_, _21818_);
  nor (_21824_, _21765_, _07130_);
  nand (_21825_, _21824_, _21813_);
  and (_21826_, _21825_, _08819_);
  and (_21828_, _21826_, _21823_);
  or (_21829_, _21804_, _08176_);
  and (_21830_, _21771_, _06303_);
  and (_21831_, _21830_, _21829_);
  or (_21832_, _21831_, _06396_);
  or (_21833_, _21832_, _21828_);
  or (_21834_, _21812_, _08824_);
  and (_21835_, _21834_, _06829_);
  and (_21836_, _21835_, _21833_);
  and (_21837_, _21775_, _06433_);
  or (_21839_, _21837_, _06440_);
  or (_21840_, _21839_, _21836_);
  or (_21841_, _21765_, _06444_);
  or (_21842_, _21841_, _21773_);
  and (_21843_, _21842_, _01317_);
  and (_21844_, _21843_, _21840_);
  or (_21845_, _21844_, _21763_);
  and (_43646_, _21845_, _43100_);
  and (_21846_, _01321_, \oc8051_golden_model_1.TL1 [2]);
  and (_21847_, _11484_, \oc8051_golden_model_1.TL1 [2]);
  or (_21849_, _21847_, _08248_);
  and (_21850_, _07837_, _08768_);
  or (_21851_, _21850_, _21847_);
  and (_21852_, _21851_, _06306_);
  and (_21853_, _21852_, _21849_);
  and (_21854_, _09211_, _07837_);
  or (_21855_, _21854_, _21847_);
  and (_21856_, _21855_, _06116_);
  and (_21857_, _14542_, _07837_);
  or (_21858_, _21857_, _21847_);
  or (_21859_, _21858_, _06161_);
  and (_21860_, _07837_, \oc8051_golden_model_1.ACC [2]);
  or (_21861_, _21860_, _21847_);
  and (_21862_, _21861_, _07056_);
  and (_21863_, _07057_, \oc8051_golden_model_1.TL1 [2]);
  or (_21864_, _21863_, _06160_);
  or (_21865_, _21864_, _21862_);
  and (_21866_, _21865_, _07075_);
  and (_21867_, _21866_, _21859_);
  and (_21868_, _07837_, _07708_);
  or (_21871_, _21868_, _21847_);
  and (_21872_, _21871_, _06217_);
  or (_21873_, _21872_, _21867_);
  and (_21874_, _21873_, _06229_);
  and (_21875_, _21861_, _06220_);
  or (_21876_, _21875_, _09842_);
  or (_21877_, _21876_, _21874_);
  or (_21878_, _21871_, _06132_);
  and (_21879_, _21878_, _06117_);
  and (_21880_, _21879_, _21877_);
  or (_21882_, _21880_, _05787_);
  or (_21883_, _21882_, _21856_);
  and (_21884_, _14630_, _07837_);
  or (_21885_, _21884_, _21847_);
  or (_21886_, _21885_, _06114_);
  and (_21887_, _21886_, _06111_);
  and (_21888_, _21887_, _21883_);
  and (_21889_, _21851_, _06110_);
  or (_21890_, _21889_, _06297_);
  or (_21891_, _21890_, _21888_);
  and (_21893_, _14646_, _07837_);
  or (_21894_, _21893_, _21847_);
  or (_21895_, _21894_, _07127_);
  and (_21896_, _21895_, _07125_);
  and (_21897_, _21896_, _21891_);
  and (_21898_, _10282_, _07837_);
  or (_21899_, _21898_, _21847_);
  and (_21900_, _21899_, _06402_);
  or (_21901_, _21900_, _21897_);
  and (_21902_, _21901_, _07132_);
  or (_21904_, _21902_, _21853_);
  and (_21905_, _21904_, _07130_);
  and (_21906_, _21861_, _06411_);
  and (_21907_, _21906_, _21849_);
  or (_21908_, _21907_, _06303_);
  or (_21909_, _21908_, _21905_);
  and (_21910_, _14643_, _07837_);
  or (_21911_, _21847_, _08819_);
  or (_21912_, _21911_, _21910_);
  and (_21913_, _21912_, _08824_);
  and (_21915_, _21913_, _21909_);
  nor (_21916_, _10281_, _11484_);
  or (_21917_, _21916_, _21847_);
  and (_21918_, _21917_, _06396_);
  or (_21919_, _21918_, _21915_);
  and (_21920_, _21919_, _06829_);
  and (_21921_, _21858_, _06433_);
  or (_21922_, _21921_, _06440_);
  or (_21923_, _21922_, _21920_);
  and (_21924_, _14710_, _07837_);
  or (_21926_, _21847_, _06444_);
  or (_21927_, _21926_, _21924_);
  and (_21928_, _21927_, _01317_);
  and (_21929_, _21928_, _21923_);
  or (_21930_, _21929_, _21846_);
  and (_43647_, _21930_, _43100_);
  and (_21931_, _11484_, \oc8051_golden_model_1.TL1 [3]);
  and (_21932_, _14738_, _07837_);
  or (_21933_, _21932_, _21931_);
  or (_21934_, _21933_, _06161_);
  and (_21936_, _07837_, \oc8051_golden_model_1.ACC [3]);
  or (_21937_, _21936_, _21931_);
  and (_21938_, _21937_, _07056_);
  and (_21939_, _07057_, \oc8051_golden_model_1.TL1 [3]);
  or (_21940_, _21939_, _06160_);
  or (_21941_, _21940_, _21938_);
  and (_21942_, _21941_, _07075_);
  and (_21943_, _21942_, _21934_);
  and (_21944_, _07837_, _07544_);
  or (_21945_, _21944_, _21931_);
  and (_21947_, _21945_, _06217_);
  or (_21948_, _21947_, _21943_);
  and (_21949_, _21948_, _06229_);
  and (_21950_, _21937_, _06220_);
  or (_21951_, _21950_, _09842_);
  or (_21952_, _21951_, _21949_);
  or (_21953_, _21945_, _06132_);
  and (_21954_, _21953_, _21952_);
  or (_21955_, _21954_, _06116_);
  and (_21956_, _09210_, _07837_);
  or (_21958_, _21931_, _06117_);
  or (_21959_, _21958_, _21956_);
  and (_21960_, _21959_, _06114_);
  and (_21961_, _21960_, _21955_);
  and (_21962_, _14825_, _07837_);
  or (_21963_, _21962_, _21931_);
  and (_21964_, _21963_, _05787_);
  or (_21965_, _21964_, _11136_);
  or (_21966_, _21965_, _21961_);
  and (_21967_, _14727_, _07837_);
  or (_21969_, _21931_, _07127_);
  or (_21970_, _21969_, _21967_);
  and (_21971_, _07837_, _08712_);
  or (_21972_, _21971_, _21931_);
  or (_21973_, _21972_, _06111_);
  and (_21974_, _21973_, _07125_);
  and (_21975_, _21974_, _21970_);
  and (_21976_, _21975_, _21966_);
  and (_21977_, _12318_, _07837_);
  or (_21978_, _21977_, _21931_);
  and (_21980_, _21978_, _06402_);
  or (_21981_, _21980_, _21976_);
  and (_21982_, _21981_, _07132_);
  or (_21983_, _21931_, _08140_);
  and (_21984_, _21972_, _06306_);
  and (_21985_, _21984_, _21983_);
  or (_21986_, _21985_, _21982_);
  and (_21987_, _21986_, _07130_);
  and (_21988_, _21937_, _06411_);
  and (_21989_, _21988_, _21983_);
  or (_21991_, _21989_, _06303_);
  or (_21992_, _21991_, _21987_);
  and (_21993_, _14724_, _07837_);
  or (_21994_, _21931_, _08819_);
  or (_21995_, _21994_, _21993_);
  and (_21996_, _21995_, _08824_);
  and (_21997_, _21996_, _21992_);
  nor (_21998_, _10273_, _11484_);
  or (_21999_, _21998_, _21931_);
  and (_22000_, _21999_, _06396_);
  or (_22002_, _22000_, _06433_);
  or (_22003_, _22002_, _21997_);
  or (_22004_, _21933_, _06829_);
  and (_22005_, _22004_, _06444_);
  and (_22006_, _22005_, _22003_);
  and (_22007_, _14897_, _07837_);
  or (_22008_, _22007_, _21931_);
  and (_22009_, _22008_, _06440_);
  or (_22010_, _22009_, _01321_);
  or (_22011_, _22010_, _22006_);
  or (_22013_, _01317_, \oc8051_golden_model_1.TL1 [3]);
  and (_22014_, _22013_, _43100_);
  and (_43648_, _22014_, _22011_);
  and (_22015_, _11484_, \oc8051_golden_model_1.TL1 [4]);
  and (_22016_, _14928_, _07837_);
  or (_22017_, _22016_, _22015_);
  or (_22018_, _22017_, _06161_);
  and (_22019_, _07837_, \oc8051_golden_model_1.ACC [4]);
  or (_22020_, _22019_, _22015_);
  and (_22021_, _22020_, _07056_);
  and (_22023_, _07057_, \oc8051_golden_model_1.TL1 [4]);
  or (_22024_, _22023_, _06160_);
  or (_22025_, _22024_, _22021_);
  and (_22026_, _22025_, _07075_);
  and (_22027_, _22026_, _22018_);
  and (_22028_, _08336_, _07837_);
  or (_22029_, _22028_, _22015_);
  and (_22030_, _22029_, _06217_);
  or (_22031_, _22030_, _22027_);
  and (_22032_, _22031_, _06229_);
  and (_22034_, _22020_, _06220_);
  or (_22035_, _22034_, _09842_);
  or (_22036_, _22035_, _22032_);
  or (_22037_, _22029_, _06132_);
  and (_22038_, _22037_, _22036_);
  or (_22039_, _22038_, _06116_);
  and (_22040_, _09209_, _07837_);
  or (_22041_, _22015_, _06117_);
  or (_22042_, _22041_, _22040_);
  and (_22043_, _22042_, _06114_);
  and (_22045_, _22043_, _22039_);
  and (_22046_, _15013_, _07837_);
  or (_22047_, _22046_, _22015_);
  and (_22048_, _22047_, _05787_);
  or (_22049_, _22048_, _22045_);
  or (_22050_, _22049_, _11136_);
  and (_22051_, _15029_, _07837_);
  or (_22052_, _22015_, _07127_);
  or (_22053_, _22052_, _22051_);
  and (_22054_, _08715_, _07837_);
  or (_22056_, _22054_, _22015_);
  or (_22057_, _22056_, _06111_);
  and (_22058_, _22057_, _07125_);
  and (_22059_, _22058_, _22053_);
  and (_22060_, _22059_, _22050_);
  and (_22061_, _10289_, _07837_);
  or (_22062_, _22061_, _22015_);
  and (_22063_, _22062_, _06402_);
  or (_22064_, _22063_, _22060_);
  and (_22065_, _22064_, _07132_);
  or (_22067_, _22015_, _08339_);
  and (_22068_, _22056_, _06306_);
  and (_22069_, _22068_, _22067_);
  or (_22070_, _22069_, _22065_);
  and (_22071_, _22070_, _07130_);
  and (_22072_, _22020_, _06411_);
  and (_22073_, _22072_, _22067_);
  or (_22074_, _22073_, _06303_);
  or (_22075_, _22074_, _22071_);
  and (_22076_, _15026_, _07837_);
  or (_22078_, _22015_, _08819_);
  or (_22079_, _22078_, _22076_);
  and (_22080_, _22079_, _08824_);
  and (_22081_, _22080_, _22075_);
  nor (_22082_, _10288_, _11484_);
  or (_22083_, _22082_, _22015_);
  and (_22084_, _22083_, _06396_);
  or (_22085_, _22084_, _06433_);
  or (_22086_, _22085_, _22081_);
  or (_22087_, _22017_, _06829_);
  and (_22089_, _22087_, _06444_);
  and (_22090_, _22089_, _22086_);
  and (_22091_, _15087_, _07837_);
  or (_22092_, _22091_, _22015_);
  and (_22093_, _22092_, _06440_);
  or (_22094_, _22093_, _01321_);
  or (_22095_, _22094_, _22090_);
  or (_22096_, _01317_, \oc8051_golden_model_1.TL1 [4]);
  and (_22097_, _22096_, _43100_);
  and (_43649_, _22097_, _22095_);
  and (_22099_, _11484_, \oc8051_golden_model_1.TL1 [5]);
  or (_22100_, _22099_, _08104_);
  and (_22101_, _08736_, _07837_);
  or (_22102_, _22101_, _22099_);
  and (_22103_, _22102_, _06306_);
  and (_22104_, _22103_, _22100_);
  and (_22105_, _15119_, _07837_);
  or (_22106_, _22105_, _22099_);
  or (_22107_, _22106_, _06161_);
  and (_22108_, _07837_, \oc8051_golden_model_1.ACC [5]);
  or (_22110_, _22108_, _22099_);
  and (_22111_, _22110_, _07056_);
  and (_22112_, _07057_, \oc8051_golden_model_1.TL1 [5]);
  or (_22113_, _22112_, _06160_);
  or (_22114_, _22113_, _22111_);
  and (_22115_, _22114_, _07075_);
  and (_22116_, _22115_, _22107_);
  and (_22117_, _08101_, _07837_);
  or (_22118_, _22117_, _22099_);
  and (_22119_, _22118_, _06217_);
  or (_22121_, _22119_, _22116_);
  and (_22122_, _22121_, _06229_);
  and (_22123_, _22110_, _06220_);
  or (_22124_, _22123_, _09842_);
  or (_22125_, _22124_, _22122_);
  or (_22126_, _22118_, _06132_);
  and (_22127_, _22126_, _22125_);
  or (_22128_, _22127_, _06116_);
  and (_22129_, _09208_, _07837_);
  or (_22130_, _22099_, _06117_);
  or (_22132_, _22130_, _22129_);
  and (_22133_, _22132_, _06114_);
  and (_22134_, _22133_, _22128_);
  and (_22135_, _15203_, _07837_);
  or (_22136_, _22135_, _22099_);
  and (_22137_, _22136_, _05787_);
  or (_22138_, _22137_, _11136_);
  or (_22139_, _22138_, _22134_);
  and (_22140_, _15219_, _07837_);
  or (_22141_, _22099_, _07127_);
  or (_22143_, _22141_, _22140_);
  or (_22144_, _22102_, _06111_);
  and (_22145_, _22144_, _07125_);
  and (_22146_, _22145_, _22143_);
  and (_22147_, _22146_, _22139_);
  and (_22148_, _12325_, _07837_);
  or (_22149_, _22148_, _22099_);
  and (_22150_, _22149_, _06402_);
  or (_22151_, _22150_, _22147_);
  and (_22152_, _22151_, _07132_);
  or (_22154_, _22152_, _22104_);
  and (_22155_, _22154_, _07130_);
  and (_22156_, _22110_, _06411_);
  and (_22157_, _22156_, _22100_);
  or (_22158_, _22157_, _06303_);
  or (_22159_, _22158_, _22155_);
  and (_22160_, _15216_, _07837_);
  or (_22161_, _22099_, _08819_);
  or (_22162_, _22161_, _22160_);
  and (_22163_, _22162_, _08824_);
  and (_22165_, _22163_, _22159_);
  nor (_22166_, _10269_, _11484_);
  or (_22167_, _22166_, _22099_);
  and (_22168_, _22167_, _06396_);
  or (_22169_, _22168_, _06433_);
  or (_22170_, _22169_, _22165_);
  or (_22171_, _22106_, _06829_);
  and (_22172_, _22171_, _06444_);
  and (_22173_, _22172_, _22170_);
  and (_22174_, _15275_, _07837_);
  or (_22176_, _22174_, _22099_);
  and (_22177_, _22176_, _06440_);
  or (_22178_, _22177_, _01321_);
  or (_22179_, _22178_, _22173_);
  or (_22180_, _01317_, \oc8051_golden_model_1.TL1 [5]);
  and (_22181_, _22180_, _43100_);
  and (_43650_, _22181_, _22179_);
  and (_22182_, _11484_, \oc8051_golden_model_1.TL1 [6]);
  or (_22183_, _22182_, _08015_);
  and (_22184_, _15402_, _07837_);
  or (_22186_, _22184_, _22182_);
  and (_22187_, _22186_, _06306_);
  and (_22188_, _22187_, _22183_);
  and (_22189_, _15300_, _07837_);
  or (_22190_, _22189_, _22182_);
  or (_22191_, _22190_, _06161_);
  and (_22192_, _07837_, \oc8051_golden_model_1.ACC [6]);
  or (_22193_, _22192_, _22182_);
  and (_22194_, _22193_, _07056_);
  and (_22195_, _07057_, \oc8051_golden_model_1.TL1 [6]);
  or (_22197_, _22195_, _06160_);
  or (_22198_, _22197_, _22194_);
  and (_22199_, _22198_, _07075_);
  and (_22200_, _22199_, _22191_);
  and (_22201_, _08012_, _07837_);
  or (_22202_, _22201_, _22182_);
  and (_22203_, _22202_, _06217_);
  or (_22204_, _22203_, _22200_);
  and (_22205_, _22204_, _06229_);
  and (_22206_, _22193_, _06220_);
  or (_22208_, _22206_, _09842_);
  or (_22209_, _22208_, _22205_);
  or (_22210_, _22202_, _06132_);
  and (_22211_, _22210_, _22209_);
  or (_22212_, _22211_, _06116_);
  and (_22213_, _09207_, _07837_);
  or (_22214_, _22182_, _06117_);
  or (_22215_, _22214_, _22213_);
  and (_22216_, _22215_, _06114_);
  and (_22217_, _22216_, _22212_);
  and (_22220_, _15395_, _07837_);
  or (_22221_, _22220_, _22182_);
  and (_22222_, _22221_, _05787_);
  or (_22223_, _22222_, _11136_);
  or (_22224_, _22223_, _22217_);
  and (_22225_, _15413_, _07837_);
  or (_22226_, _22182_, _07127_);
  or (_22227_, _22226_, _22225_);
  or (_22228_, _22186_, _06111_);
  and (_22229_, _22228_, _07125_);
  and (_22231_, _22229_, _22227_);
  and (_22232_, _22231_, _22224_);
  and (_22233_, _10295_, _07837_);
  or (_22234_, _22233_, _22182_);
  and (_22235_, _22234_, _06402_);
  or (_22236_, _22235_, _22232_);
  and (_22237_, _22236_, _07132_);
  or (_22238_, _22237_, _22188_);
  and (_22239_, _22238_, _07130_);
  and (_22240_, _22193_, _06411_);
  and (_22242_, _22240_, _22183_);
  or (_22243_, _22242_, _06303_);
  or (_22244_, _22243_, _22239_);
  and (_22245_, _15410_, _07837_);
  or (_22246_, _22182_, _08819_);
  or (_22247_, _22246_, _22245_);
  and (_22248_, _22247_, _08824_);
  and (_22249_, _22248_, _22244_);
  nor (_22250_, _10294_, _11484_);
  or (_22251_, _22250_, _22182_);
  and (_22253_, _22251_, _06396_);
  or (_22254_, _22253_, _06433_);
  or (_22255_, _22254_, _22249_);
  or (_22256_, _22190_, _06829_);
  and (_22257_, _22256_, _06444_);
  and (_22258_, _22257_, _22255_);
  and (_22259_, _15478_, _07837_);
  or (_22260_, _22259_, _22182_);
  and (_22261_, _22260_, _06440_);
  or (_22262_, _22261_, _01321_);
  or (_22264_, _22262_, _22258_);
  or (_22265_, _01317_, \oc8051_golden_model_1.TL1 [6]);
  and (_22266_, _22265_, _43100_);
  and (_43651_, _22266_, _22264_);
  not (_22267_, \oc8051_golden_model_1.TL0 [0]);
  nor (_22268_, _01317_, _22267_);
  nand (_22269_, _10276_, _07803_);
  nor (_22270_, _07803_, _22267_);
  nor (_22271_, _22270_, _07130_);
  nand (_22272_, _22271_, _22269_);
  and (_22274_, _07803_, _07049_);
  or (_22275_, _22274_, _22270_);
  or (_22276_, _22275_, _06132_);
  nor (_22277_, _08211_, _11561_);
  or (_22278_, _22277_, _22270_);
  or (_22279_, _22278_, _06161_);
  and (_22280_, _07803_, \oc8051_golden_model_1.ACC [0]);
  or (_22281_, _22280_, _22270_);
  and (_22282_, _22281_, _07056_);
  nor (_22283_, _07056_, _22267_);
  or (_22285_, _22283_, _06160_);
  or (_22286_, _22285_, _22282_);
  and (_22287_, _22286_, _07075_);
  and (_22288_, _22287_, _22279_);
  and (_22289_, _22275_, _06217_);
  or (_22290_, _22289_, _22288_);
  and (_22291_, _22290_, _06229_);
  and (_22292_, _22281_, _06220_);
  or (_22293_, _22292_, _09842_);
  or (_22294_, _22293_, _22291_);
  and (_22296_, _22294_, _22276_);
  or (_22297_, _22296_, _06116_);
  and (_22298_, _09160_, _07803_);
  or (_22299_, _22270_, _06117_);
  or (_22300_, _22299_, _22298_);
  and (_22301_, _22300_, _22297_);
  or (_22302_, _22301_, _05787_);
  and (_22303_, _14260_, _07803_);
  or (_22304_, _22303_, _22270_);
  or (_22305_, _22304_, _06114_);
  and (_22306_, _22305_, _06111_);
  and (_22307_, _22306_, _22302_);
  and (_22308_, _07803_, _08708_);
  or (_22309_, _22308_, _22270_);
  and (_22310_, _22309_, _06110_);
  or (_22311_, _22310_, _06297_);
  or (_22312_, _22311_, _22307_);
  and (_22313_, _14275_, _07803_);
  or (_22314_, _22270_, _07127_);
  or (_22315_, _22314_, _22313_);
  and (_22318_, _22315_, _07125_);
  and (_22319_, _22318_, _22312_);
  nor (_22320_, _12321_, _11561_);
  or (_22321_, _22320_, _22270_);
  and (_22322_, _22269_, _06402_);
  and (_22323_, _22322_, _22321_);
  or (_22324_, _22323_, _22319_);
  and (_22325_, _22324_, _07132_);
  nand (_22326_, _22309_, _06306_);
  nor (_22327_, _22326_, _22277_);
  or (_22329_, _22327_, _06411_);
  or (_22330_, _22329_, _22325_);
  and (_22331_, _22330_, _22272_);
  or (_22332_, _22331_, _06303_);
  and (_22333_, _14167_, _07803_);
  or (_22334_, _22333_, _22270_);
  or (_22335_, _22334_, _08819_);
  and (_22336_, _22335_, _08824_);
  and (_22337_, _22336_, _22332_);
  and (_22338_, _22321_, _06396_);
  or (_22340_, _22338_, _19287_);
  or (_22341_, _22340_, _22337_);
  or (_22342_, _22278_, _06630_);
  and (_22343_, _22342_, _01317_);
  and (_22344_, _22343_, _22341_);
  or (_22345_, _22344_, _22268_);
  and (_43653_, _22345_, _43100_);
  and (_22346_, _11561_, \oc8051_golden_model_1.TL0 [1]);
  nor (_22347_, _10277_, _11561_);
  or (_22348_, _22347_, _22346_);
  or (_22350_, _22348_, _08824_);
  or (_22351_, _14442_, _11561_);
  or (_22352_, _07803_, \oc8051_golden_model_1.TL0 [1]);
  and (_22353_, _22352_, _05787_);
  and (_22354_, _22353_, _22351_);
  and (_22355_, _09115_, _07803_);
  or (_22356_, _22346_, _06117_);
  or (_22357_, _22356_, _22355_);
  and (_22358_, _14363_, _07803_);
  not (_22359_, _22358_);
  and (_22361_, _22359_, _22352_);
  or (_22362_, _22361_, _06161_);
  and (_22363_, _07803_, \oc8051_golden_model_1.ACC [1]);
  or (_22364_, _22363_, _22346_);
  and (_22365_, _22364_, _07056_);
  and (_22366_, _07057_, \oc8051_golden_model_1.TL0 [1]);
  or (_22367_, _22366_, _06160_);
  or (_22368_, _22367_, _22365_);
  and (_22369_, _22368_, _07075_);
  and (_22370_, _22369_, _22362_);
  and (_22372_, _07803_, _07306_);
  or (_22373_, _22372_, _22346_);
  and (_22374_, _22373_, _06217_);
  or (_22375_, _22374_, _22370_);
  and (_22376_, _22375_, _06229_);
  and (_22377_, _22364_, _06220_);
  or (_22378_, _22377_, _09842_);
  or (_22379_, _22378_, _22376_);
  or (_22380_, _22373_, _06132_);
  and (_22381_, _22380_, _22379_);
  or (_22383_, _22381_, _06116_);
  and (_22384_, _22383_, _06114_);
  and (_22385_, _22384_, _22357_);
  or (_22386_, _22385_, _22354_);
  and (_22387_, _22386_, _06298_);
  or (_22388_, _14346_, _11561_);
  and (_22389_, _22388_, _06297_);
  nand (_22390_, _07803_, _06945_);
  and (_22391_, _22390_, _06110_);
  or (_22392_, _22391_, _22389_);
  and (_22394_, _22392_, _22352_);
  or (_22395_, _22394_, _06402_);
  or (_22396_, _22395_, _22387_);
  nand (_22397_, _10275_, _07803_);
  and (_22398_, _22397_, _22348_);
  or (_22399_, _22398_, _07125_);
  and (_22400_, _22399_, _07132_);
  and (_22401_, _22400_, _22396_);
  or (_22402_, _14344_, _11561_);
  and (_22403_, _22352_, _06306_);
  and (_22405_, _22403_, _22402_);
  or (_22406_, _22405_, _06411_);
  or (_22407_, _22406_, _22401_);
  nor (_22408_, _22346_, _07130_);
  nand (_22409_, _22408_, _22397_);
  and (_22410_, _22409_, _08819_);
  and (_22411_, _22410_, _22407_);
  or (_22412_, _22390_, _08176_);
  and (_22413_, _22352_, _06303_);
  and (_22414_, _22413_, _22412_);
  or (_22416_, _22414_, _06396_);
  or (_22417_, _22416_, _22411_);
  and (_22418_, _22417_, _22350_);
  or (_22419_, _22418_, _06433_);
  or (_22420_, _22361_, _06829_);
  and (_22421_, _22420_, _06444_);
  and (_22422_, _22421_, _22419_);
  or (_22423_, _22358_, _22346_);
  and (_22424_, _22423_, _06440_);
  or (_22425_, _22424_, _01321_);
  or (_22427_, _22425_, _22422_);
  or (_22428_, _01317_, \oc8051_golden_model_1.TL0 [1]);
  and (_22429_, _22428_, _43100_);
  and (_43654_, _22429_, _22427_);
  and (_22430_, _01321_, \oc8051_golden_model_1.TL0 [2]);
  and (_22431_, _11561_, \oc8051_golden_model_1.TL0 [2]);
  and (_22432_, _09211_, _07803_);
  or (_22433_, _22432_, _22431_);
  and (_22434_, _22433_, _06116_);
  and (_22435_, _14542_, _07803_);
  or (_22437_, _22435_, _22431_);
  or (_22438_, _22437_, _06161_);
  and (_22439_, _07803_, \oc8051_golden_model_1.ACC [2]);
  or (_22440_, _22439_, _22431_);
  and (_22441_, _22440_, _07056_);
  and (_22442_, _07057_, \oc8051_golden_model_1.TL0 [2]);
  or (_22443_, _22442_, _06160_);
  or (_22444_, _22443_, _22441_);
  and (_22445_, _22444_, _07075_);
  and (_22446_, _22445_, _22438_);
  and (_22448_, _07803_, _07708_);
  or (_22449_, _22448_, _22431_);
  and (_22450_, _22449_, _06217_);
  or (_22451_, _22450_, _22446_);
  and (_22452_, _22451_, _06229_);
  and (_22453_, _22440_, _06220_);
  or (_22454_, _22453_, _09842_);
  or (_22455_, _22454_, _22452_);
  or (_22456_, _22449_, _06132_);
  and (_22457_, _22456_, _06117_);
  and (_22459_, _22457_, _22455_);
  or (_22460_, _22459_, _05787_);
  or (_22461_, _22460_, _22434_);
  and (_22462_, _14630_, _07803_);
  or (_22463_, _22431_, _06114_);
  or (_22464_, _22463_, _22462_);
  and (_22465_, _22464_, _06111_);
  and (_22466_, _22465_, _22461_);
  and (_22467_, _07803_, _08768_);
  or (_22468_, _22467_, _22431_);
  and (_22470_, _22468_, _06110_);
  or (_22471_, _22470_, _06297_);
  or (_22472_, _22471_, _22466_);
  and (_22473_, _14646_, _07803_);
  or (_22474_, _22473_, _22431_);
  or (_22475_, _22474_, _07127_);
  and (_22476_, _22475_, _07125_);
  and (_22477_, _22476_, _22472_);
  and (_22478_, _10282_, _07803_);
  or (_22479_, _22478_, _22431_);
  and (_22481_, _22479_, _06402_);
  or (_22482_, _22481_, _22477_);
  and (_22483_, _22482_, _07132_);
  or (_22484_, _22431_, _08248_);
  and (_22485_, _22468_, _06306_);
  and (_22486_, _22485_, _22484_);
  or (_22487_, _22486_, _22483_);
  and (_22488_, _22487_, _07130_);
  and (_22489_, _22440_, _06411_);
  and (_22490_, _22489_, _22484_);
  or (_22492_, _22490_, _06303_);
  or (_22493_, _22492_, _22488_);
  and (_22494_, _14643_, _07803_);
  or (_22495_, _22431_, _08819_);
  or (_22496_, _22495_, _22494_);
  and (_22497_, _22496_, _08824_);
  and (_22498_, _22497_, _22493_);
  nor (_22499_, _10281_, _11561_);
  or (_22500_, _22499_, _22431_);
  and (_22501_, _22500_, _06396_);
  or (_22503_, _22501_, _22498_);
  and (_22504_, _22503_, _06829_);
  and (_22505_, _22437_, _06433_);
  or (_22506_, _22505_, _06440_);
  or (_22507_, _22506_, _22504_);
  and (_22508_, _14710_, _07803_);
  or (_22509_, _22431_, _06444_);
  or (_22510_, _22509_, _22508_);
  and (_22511_, _22510_, _01317_);
  and (_22512_, _22511_, _22507_);
  or (_22514_, _22512_, _22430_);
  and (_43655_, _22514_, _43100_);
  and (_22515_, _11561_, \oc8051_golden_model_1.TL0 [3]);
  or (_22516_, _22515_, _08140_);
  and (_22517_, _07803_, _08712_);
  or (_22518_, _22517_, _22515_);
  and (_22519_, _22518_, _06306_);
  and (_22520_, _22519_, _22516_);
  and (_22521_, _14738_, _07803_);
  or (_22522_, _22521_, _22515_);
  or (_22524_, _22522_, _06161_);
  and (_22525_, _07803_, \oc8051_golden_model_1.ACC [3]);
  or (_22526_, _22525_, _22515_);
  and (_22527_, _22526_, _07056_);
  and (_22528_, _07057_, \oc8051_golden_model_1.TL0 [3]);
  or (_22529_, _22528_, _06160_);
  or (_22530_, _22529_, _22527_);
  and (_22531_, _22530_, _07075_);
  and (_22532_, _22531_, _22524_);
  and (_22533_, _07803_, _07544_);
  or (_22535_, _22533_, _22515_);
  and (_22536_, _22535_, _06217_);
  or (_22537_, _22536_, _22532_);
  and (_22538_, _22537_, _06229_);
  and (_22539_, _22526_, _06220_);
  or (_22540_, _22539_, _09842_);
  or (_22541_, _22540_, _22538_);
  or (_22542_, _22535_, _06132_);
  and (_22543_, _22542_, _06117_);
  and (_22544_, _22543_, _22541_);
  and (_22546_, _09210_, _07803_);
  or (_22547_, _22546_, _22515_);
  and (_22548_, _22547_, _06116_);
  or (_22549_, _22548_, _05787_);
  or (_22550_, _22549_, _22544_);
  and (_22551_, _14825_, _07803_);
  or (_22552_, _22551_, _22515_);
  or (_22553_, _22552_, _06114_);
  and (_22554_, _22553_, _06111_);
  and (_22555_, _22554_, _22550_);
  and (_22557_, _22518_, _06110_);
  or (_22558_, _22557_, _06297_);
  or (_22559_, _22558_, _22555_);
  and (_22560_, _14727_, _07803_);
  or (_22561_, _22515_, _07127_);
  or (_22562_, _22561_, _22560_);
  and (_22563_, _22562_, _07125_);
  and (_22564_, _22563_, _22559_);
  and (_22565_, _12318_, _07803_);
  or (_22566_, _22565_, _22515_);
  and (_22568_, _22566_, _06402_);
  or (_22569_, _22568_, _22564_);
  and (_22570_, _22569_, _07132_);
  or (_22571_, _22570_, _22520_);
  and (_22572_, _22571_, _07130_);
  and (_22573_, _22526_, _06411_);
  and (_22574_, _22573_, _22516_);
  or (_22575_, _22574_, _06303_);
  or (_22576_, _22575_, _22572_);
  and (_22577_, _14724_, _07803_);
  or (_22579_, _22515_, _08819_);
  or (_22580_, _22579_, _22577_);
  and (_22581_, _22580_, _08824_);
  and (_22582_, _22581_, _22576_);
  nor (_22583_, _10273_, _11561_);
  or (_22584_, _22583_, _22515_);
  and (_22585_, _22584_, _06396_);
  or (_22586_, _22585_, _06433_);
  or (_22587_, _22586_, _22582_);
  or (_22588_, _22522_, _06829_);
  and (_22590_, _22588_, _06444_);
  and (_22591_, _22590_, _22587_);
  and (_22592_, _14897_, _07803_);
  or (_22593_, _22592_, _22515_);
  and (_22594_, _22593_, _06440_);
  or (_22595_, _22594_, _01321_);
  or (_22596_, _22595_, _22591_);
  or (_22597_, _01317_, \oc8051_golden_model_1.TL0 [3]);
  and (_22598_, _22597_, _43100_);
  and (_43656_, _22598_, _22596_);
  and (_22599_, _11561_, \oc8051_golden_model_1.TL0 [4]);
  and (_22600_, _08336_, _07803_);
  or (_22601_, _22600_, _22599_);
  or (_22602_, _22601_, _06132_);
  and (_22603_, _14928_, _07803_);
  or (_22604_, _22603_, _22599_);
  or (_22605_, _22604_, _06161_);
  and (_22606_, _07803_, \oc8051_golden_model_1.ACC [4]);
  or (_22607_, _22606_, _22599_);
  and (_22608_, _22607_, _07056_);
  and (_22611_, _07057_, \oc8051_golden_model_1.TL0 [4]);
  or (_22612_, _22611_, _06160_);
  or (_22613_, _22612_, _22608_);
  and (_22614_, _22613_, _07075_);
  and (_22615_, _22614_, _22605_);
  and (_22616_, _22601_, _06217_);
  or (_22617_, _22616_, _22615_);
  and (_22618_, _22617_, _06229_);
  and (_22619_, _22607_, _06220_);
  or (_22620_, _22619_, _09842_);
  or (_22622_, _22620_, _22618_);
  and (_22623_, _22622_, _22602_);
  or (_22624_, _22623_, _06116_);
  and (_22625_, _09209_, _07803_);
  or (_22626_, _22599_, _06117_);
  or (_22627_, _22626_, _22625_);
  and (_22628_, _22627_, _06114_);
  and (_22629_, _22628_, _22624_);
  and (_22630_, _15013_, _07803_);
  or (_22631_, _22630_, _22599_);
  and (_22633_, _22631_, _05787_);
  or (_22634_, _22633_, _22629_);
  or (_22635_, _22634_, _11136_);
  and (_22636_, _15029_, _07803_);
  or (_22637_, _22599_, _07127_);
  or (_22638_, _22637_, _22636_);
  and (_22639_, _08715_, _07803_);
  or (_22640_, _22639_, _22599_);
  or (_22641_, _22640_, _06111_);
  and (_22642_, _22641_, _07125_);
  and (_22644_, _22642_, _22638_);
  and (_22645_, _22644_, _22635_);
  and (_22646_, _10289_, _07803_);
  or (_22647_, _22646_, _22599_);
  and (_22648_, _22647_, _06402_);
  or (_22649_, _22648_, _22645_);
  and (_22650_, _22649_, _07132_);
  or (_22651_, _22599_, _08339_);
  and (_22652_, _22640_, _06306_);
  and (_22653_, _22652_, _22651_);
  or (_22655_, _22653_, _22650_);
  and (_22656_, _22655_, _07130_);
  and (_22657_, _22607_, _06411_);
  and (_22658_, _22657_, _22651_);
  or (_22659_, _22658_, _06303_);
  or (_22660_, _22659_, _22656_);
  and (_22661_, _15026_, _07803_);
  or (_22662_, _22599_, _08819_);
  or (_22663_, _22662_, _22661_);
  and (_22664_, _22663_, _08824_);
  and (_22666_, _22664_, _22660_);
  nor (_22667_, _10288_, _11561_);
  or (_22668_, _22667_, _22599_);
  and (_22669_, _22668_, _06396_);
  or (_22670_, _22669_, _06433_);
  or (_22671_, _22670_, _22666_);
  or (_22672_, _22604_, _06829_);
  and (_22673_, _22672_, _06444_);
  and (_22674_, _22673_, _22671_);
  and (_22675_, _15087_, _07803_);
  or (_22677_, _22675_, _22599_);
  and (_22678_, _22677_, _06440_);
  or (_22679_, _22678_, _01321_);
  or (_22680_, _22679_, _22674_);
  or (_22681_, _01317_, \oc8051_golden_model_1.TL0 [4]);
  and (_22682_, _22681_, _43100_);
  and (_43657_, _22682_, _22680_);
  and (_22683_, _11561_, \oc8051_golden_model_1.TL0 [5]);
  or (_22684_, _22683_, _08104_);
  and (_22685_, _08736_, _07803_);
  or (_22687_, _22685_, _22683_);
  and (_22688_, _22687_, _06306_);
  and (_22689_, _22688_, _22684_);
  and (_22690_, _15119_, _07803_);
  or (_22691_, _22690_, _22683_);
  or (_22692_, _22691_, _06161_);
  and (_22693_, _07803_, \oc8051_golden_model_1.ACC [5]);
  or (_22694_, _22693_, _22683_);
  and (_22695_, _22694_, _07056_);
  and (_22696_, _07057_, \oc8051_golden_model_1.TL0 [5]);
  or (_22698_, _22696_, _06160_);
  or (_22699_, _22698_, _22695_);
  and (_22700_, _22699_, _07075_);
  and (_22701_, _22700_, _22692_);
  and (_22702_, _08101_, _07803_);
  or (_22703_, _22702_, _22683_);
  and (_22704_, _22703_, _06217_);
  or (_22705_, _22704_, _22701_);
  and (_22706_, _22705_, _06229_);
  and (_22707_, _22694_, _06220_);
  or (_22708_, _22707_, _09842_);
  or (_22709_, _22708_, _22706_);
  or (_22710_, _22703_, _06132_);
  and (_22711_, _22710_, _22709_);
  or (_22712_, _22711_, _06116_);
  and (_22713_, _09208_, _07803_);
  or (_22714_, _22683_, _06117_);
  or (_22715_, _22714_, _22713_);
  and (_22716_, _22715_, _06114_);
  and (_22717_, _22716_, _22712_);
  and (_22720_, _15203_, _07803_);
  or (_22721_, _22720_, _22683_);
  and (_22722_, _22721_, _05787_);
  or (_22723_, _22722_, _11136_);
  or (_22724_, _22723_, _22717_);
  and (_22725_, _15219_, _07803_);
  or (_22726_, _22683_, _07127_);
  or (_22727_, _22726_, _22725_);
  or (_22728_, _22687_, _06111_);
  and (_22729_, _22728_, _07125_);
  and (_22731_, _22729_, _22727_);
  and (_22732_, _22731_, _22724_);
  and (_22733_, _12325_, _07803_);
  or (_22734_, _22733_, _22683_);
  and (_22735_, _22734_, _06402_);
  or (_22736_, _22735_, _22732_);
  and (_22737_, _22736_, _07132_);
  or (_22738_, _22737_, _22689_);
  and (_22739_, _22738_, _07130_);
  and (_22740_, _22694_, _06411_);
  and (_22742_, _22740_, _22684_);
  or (_22743_, _22742_, _06303_);
  or (_22744_, _22743_, _22739_);
  and (_22745_, _15216_, _07803_);
  or (_22746_, _22683_, _08819_);
  or (_22747_, _22746_, _22745_);
  and (_22748_, _22747_, _08824_);
  and (_22749_, _22748_, _22744_);
  nor (_22750_, _10269_, _11561_);
  or (_22751_, _22750_, _22683_);
  and (_22753_, _22751_, _06396_);
  or (_22754_, _22753_, _06433_);
  or (_22755_, _22754_, _22749_);
  or (_22756_, _22691_, _06829_);
  and (_22757_, _22756_, _06444_);
  and (_22758_, _22757_, _22755_);
  and (_22759_, _15275_, _07803_);
  or (_22760_, _22759_, _22683_);
  and (_22761_, _22760_, _06440_);
  or (_22762_, _22761_, _01321_);
  or (_22764_, _22762_, _22758_);
  or (_22765_, _01317_, \oc8051_golden_model_1.TL0 [5]);
  and (_22766_, _22765_, _43100_);
  and (_43659_, _22766_, _22764_);
  and (_22767_, _11561_, \oc8051_golden_model_1.TL0 [6]);
  or (_22768_, _22767_, _08015_);
  and (_22769_, _15402_, _07803_);
  or (_22770_, _22769_, _22767_);
  and (_22771_, _22770_, _06306_);
  and (_22772_, _22771_, _22768_);
  and (_22774_, _15300_, _07803_);
  or (_22775_, _22774_, _22767_);
  or (_22776_, _22775_, _06161_);
  and (_22777_, _07803_, \oc8051_golden_model_1.ACC [6]);
  or (_22778_, _22777_, _22767_);
  and (_22779_, _22778_, _07056_);
  and (_22780_, _07057_, \oc8051_golden_model_1.TL0 [6]);
  or (_22781_, _22780_, _06160_);
  or (_22782_, _22781_, _22779_);
  and (_22783_, _22782_, _07075_);
  and (_22785_, _22783_, _22776_);
  and (_22786_, _08012_, _07803_);
  or (_22787_, _22786_, _22767_);
  and (_22788_, _22787_, _06217_);
  or (_22789_, _22788_, _22785_);
  and (_22790_, _22789_, _06229_);
  and (_22791_, _22778_, _06220_);
  or (_22792_, _22791_, _09842_);
  or (_22793_, _22792_, _22790_);
  or (_22794_, _22787_, _06132_);
  and (_22796_, _22794_, _22793_);
  or (_22797_, _22796_, _06116_);
  and (_22798_, _09207_, _07803_);
  or (_22799_, _22767_, _06117_);
  or (_22800_, _22799_, _22798_);
  and (_22801_, _22800_, _06114_);
  and (_22802_, _22801_, _22797_);
  and (_22803_, _15395_, _07803_);
  or (_22804_, _22803_, _22767_);
  and (_22805_, _22804_, _05787_);
  or (_22807_, _22805_, _11136_);
  or (_22808_, _22807_, _22802_);
  and (_22809_, _15413_, _07803_);
  or (_22810_, _22767_, _07127_);
  or (_22811_, _22810_, _22809_);
  or (_22812_, _22770_, _06111_);
  and (_22813_, _22812_, _07125_);
  and (_22814_, _22813_, _22811_);
  and (_22815_, _22814_, _22808_);
  and (_22816_, _10295_, _07803_);
  or (_22818_, _22816_, _22767_);
  and (_22819_, _22818_, _06402_);
  or (_22820_, _22819_, _22815_);
  and (_22821_, _22820_, _07132_);
  or (_22822_, _22821_, _22772_);
  and (_22823_, _22822_, _07130_);
  and (_22824_, _22778_, _06411_);
  and (_22825_, _22824_, _22768_);
  or (_22826_, _22825_, _06303_);
  or (_22827_, _22826_, _22823_);
  and (_22829_, _15410_, _07803_);
  or (_22830_, _22767_, _08819_);
  or (_22831_, _22830_, _22829_);
  and (_22832_, _22831_, _08824_);
  and (_22833_, _22832_, _22827_);
  nor (_22834_, _10294_, _11561_);
  or (_22835_, _22834_, _22767_);
  and (_22836_, _22835_, _06396_);
  or (_22837_, _22836_, _06433_);
  or (_22838_, _22837_, _22833_);
  or (_22840_, _22775_, _06829_);
  and (_22841_, _22840_, _06444_);
  and (_22842_, _22841_, _22838_);
  and (_22843_, _15478_, _07803_);
  or (_22844_, _22843_, _22767_);
  and (_22845_, _22844_, _06440_);
  or (_22846_, _22845_, _01321_);
  or (_22847_, _22846_, _22842_);
  or (_22848_, _01317_, \oc8051_golden_model_1.TL0 [6]);
  and (_22849_, _22848_, _43100_);
  and (_43660_, _22849_, _22847_);
  not (_22851_, \oc8051_golden_model_1.TCON [0]);
  nor (_22852_, _01317_, _22851_);
  nand (_22853_, _10276_, _07788_);
  nor (_22854_, _07788_, _22851_);
  nor (_22855_, _22854_, _07130_);
  nand (_22856_, _22855_, _22853_);
  and (_22857_, _07788_, _07049_);
  or (_22858_, _22857_, _22854_);
  or (_22859_, _22858_, _06132_);
  nor (_22861_, _08211_, _11639_);
  or (_22862_, _22861_, _22854_);
  or (_22863_, _22862_, _06161_);
  and (_22864_, _07788_, \oc8051_golden_model_1.ACC [0]);
  or (_22865_, _22864_, _22854_);
  and (_22866_, _22865_, _07056_);
  nor (_22867_, _07056_, _22851_);
  or (_22868_, _22867_, _06160_);
  or (_22869_, _22868_, _22866_);
  and (_22870_, _22869_, _06157_);
  and (_22872_, _22870_, _22863_);
  nor (_22873_, _08407_, _22851_);
  and (_22874_, _14169_, _08407_);
  or (_22875_, _22874_, _22873_);
  and (_22876_, _22875_, _06156_);
  or (_22877_, _22876_, _22872_);
  and (_22878_, _22877_, _07075_);
  and (_22879_, _22858_, _06217_);
  or (_22880_, _22879_, _06220_);
  or (_22881_, _22880_, _22878_);
  or (_22883_, _22865_, _06229_);
  and (_22884_, _22883_, _06153_);
  and (_22885_, _22884_, _22881_);
  and (_22886_, _22854_, _06152_);
  or (_22887_, _22886_, _06145_);
  or (_22888_, _22887_, _22885_);
  or (_22889_, _22862_, _06146_);
  and (_22890_, _22889_, _06140_);
  and (_22891_, _22890_, _22888_);
  or (_22892_, _22873_, _14170_);
  and (_22894_, _22892_, _06139_);
  and (_22895_, _22894_, _22875_);
  or (_22896_, _22895_, _09842_);
  or (_22897_, _22896_, _22891_);
  and (_22898_, _22897_, _22859_);
  or (_22899_, _22898_, _06116_);
  and (_22900_, _09160_, _07788_);
  or (_22901_, _22854_, _06117_);
  or (_22902_, _22901_, _22900_);
  and (_22903_, _22902_, _06114_);
  and (_22905_, _22903_, _22899_);
  and (_22906_, _14260_, _07788_);
  or (_22907_, _22906_, _22854_);
  and (_22908_, _22907_, _05787_);
  or (_22909_, _22908_, _22905_);
  or (_22910_, _22909_, _11136_);
  and (_22911_, _14275_, _07788_);
  or (_22912_, _22854_, _07127_);
  or (_22913_, _22912_, _22911_);
  and (_22914_, _07788_, _08708_);
  or (_22916_, _22914_, _22854_);
  or (_22917_, _22916_, _06111_);
  and (_22918_, _22917_, _07125_);
  and (_22919_, _22918_, _22913_);
  and (_22920_, _22919_, _22910_);
  nor (_22921_, _12321_, _11639_);
  or (_22922_, _22921_, _22854_);
  and (_22923_, _22853_, _06402_);
  and (_22924_, _22923_, _22922_);
  or (_22925_, _22924_, _22920_);
  and (_22926_, _22925_, _07132_);
  nand (_22927_, _22916_, _06306_);
  nor (_22928_, _22927_, _22861_);
  or (_22929_, _22928_, _06411_);
  or (_22930_, _22929_, _22926_);
  and (_22931_, _22930_, _22856_);
  or (_22932_, _22931_, _06303_);
  and (_22933_, _14167_, _07788_);
  or (_22934_, _22854_, _08819_);
  or (_22935_, _22934_, _22933_);
  and (_22938_, _22935_, _08824_);
  and (_22939_, _22938_, _22932_);
  and (_22940_, _22922_, _06396_);
  or (_22941_, _22940_, _06433_);
  or (_22942_, _22941_, _22939_);
  or (_22943_, _22862_, _06829_);
  and (_22944_, _22943_, _22942_);
  or (_22945_, _22944_, _05748_);
  or (_22946_, _22854_, _05749_);
  and (_22947_, _22946_, _22945_);
  or (_22949_, _22947_, _06440_);
  or (_22950_, _22862_, _06444_);
  and (_22951_, _22950_, _01317_);
  and (_22952_, _22951_, _22949_);
  or (_22953_, _22952_, _22852_);
  and (_43661_, _22953_, _43100_);
  and (_22954_, _01321_, \oc8051_golden_model_1.TCON [1]);
  and (_22955_, _11639_, \oc8051_golden_model_1.TCON [1]);
  nor (_22956_, _10277_, _11639_);
  or (_22957_, _22956_, _22955_);
  or (_22959_, _22957_, _08824_);
  or (_22960_, _14442_, _11639_);
  or (_22961_, _07788_, \oc8051_golden_model_1.TCON [1]);
  and (_22962_, _22961_, _05787_);
  and (_22963_, _22962_, _22960_);
  and (_22964_, _07788_, _07306_);
  or (_22965_, _22964_, _22955_);
  or (_22966_, _22965_, _07075_);
  and (_22967_, _14363_, _07788_);
  not (_22968_, _22967_);
  and (_22970_, _22968_, _22961_);
  or (_22971_, _22970_, _06161_);
  and (_22972_, _07788_, \oc8051_golden_model_1.ACC [1]);
  or (_22973_, _22972_, _22955_);
  and (_22974_, _22973_, _07056_);
  and (_22975_, _07057_, \oc8051_golden_model_1.TCON [1]);
  or (_22976_, _22975_, _06160_);
  or (_22977_, _22976_, _22974_);
  and (_22978_, _22977_, _06157_);
  and (_22979_, _22978_, _22971_);
  and (_22981_, _11644_, \oc8051_golden_model_1.TCON [1]);
  and (_22982_, _14367_, _08407_);
  or (_22983_, _22982_, _22981_);
  and (_22984_, _22983_, _06156_);
  or (_22985_, _22984_, _06217_);
  or (_22986_, _22985_, _22979_);
  and (_22987_, _22986_, _22966_);
  or (_22988_, _22987_, _06220_);
  or (_22989_, _22973_, _06229_);
  and (_22990_, _22989_, _06153_);
  and (_22992_, _22990_, _22988_);
  and (_22993_, _14349_, _08407_);
  or (_22994_, _22993_, _22981_);
  and (_22995_, _22994_, _06152_);
  or (_22996_, _22995_, _06145_);
  or (_22997_, _22996_, _22992_);
  and (_22998_, _22982_, _14382_);
  or (_22999_, _22981_, _06146_);
  or (_23000_, _22999_, _22998_);
  and (_23001_, _23000_, _22997_);
  and (_23003_, _23001_, _06140_);
  and (_23004_, _14351_, _08407_);
  or (_23005_, _22981_, _23004_);
  and (_23006_, _23005_, _06139_);
  or (_23007_, _23006_, _09842_);
  or (_23008_, _23007_, _23003_);
  or (_23009_, _22965_, _06132_);
  and (_23010_, _23009_, _23008_);
  or (_23011_, _23010_, _06116_);
  and (_23012_, _09115_, _07788_);
  or (_23014_, _22955_, _06117_);
  or (_23015_, _23014_, _23012_);
  and (_23016_, _23015_, _06114_);
  and (_23017_, _23016_, _23011_);
  or (_23018_, _23017_, _22963_);
  and (_23019_, _23018_, _06298_);
  or (_23020_, _14346_, _11639_);
  and (_23021_, _23020_, _06297_);
  nand (_23022_, _07788_, _06945_);
  and (_23023_, _23022_, _06110_);
  or (_23025_, _23023_, _23021_);
  and (_23026_, _23025_, _22961_);
  or (_23027_, _23026_, _06402_);
  or (_23028_, _23027_, _23019_);
  and (_23029_, _10278_, _07788_);
  or (_23030_, _23029_, _22955_);
  or (_23031_, _23030_, _07125_);
  and (_23032_, _23031_, _07132_);
  and (_23033_, _23032_, _23028_);
  or (_23034_, _14344_, _11639_);
  and (_23036_, _22961_, _06306_);
  and (_23037_, _23036_, _23034_);
  or (_23038_, _23037_, _06411_);
  or (_23039_, _23038_, _23033_);
  and (_23040_, _22972_, _08176_);
  or (_23041_, _22955_, _07130_);
  or (_23042_, _23041_, _23040_);
  and (_23043_, _23042_, _08819_);
  and (_23044_, _23043_, _23039_);
  or (_23045_, _23022_, _08176_);
  and (_23046_, _22961_, _06303_);
  and (_23047_, _23046_, _23045_);
  or (_23048_, _23047_, _06396_);
  or (_23049_, _23048_, _23044_);
  and (_23050_, _23049_, _22959_);
  or (_23051_, _23050_, _06433_);
  or (_23052_, _22970_, _06829_);
  and (_23053_, _23052_, _05749_);
  and (_23054_, _23053_, _23051_);
  and (_23055_, _22994_, _05748_);
  or (_23057_, _23055_, _06440_);
  or (_23058_, _23057_, _23054_);
  or (_23059_, _22955_, _06444_);
  or (_23060_, _23059_, _22967_);
  and (_23061_, _23060_, _01317_);
  and (_23062_, _23061_, _23058_);
  or (_23063_, _23062_, _22954_);
  and (_43663_, _23063_, _43100_);
  and (_23064_, _01321_, \oc8051_golden_model_1.TCON [2]);
  and (_23065_, _11639_, \oc8051_golden_model_1.TCON [2]);
  and (_23067_, _07788_, _07708_);
  or (_23068_, _23067_, _23065_);
  or (_23069_, _23068_, _06132_);
  or (_23070_, _23068_, _07075_);
  and (_23071_, _14542_, _07788_);
  or (_23072_, _23071_, _23065_);
  or (_23073_, _23072_, _06161_);
  and (_23074_, _07788_, \oc8051_golden_model_1.ACC [2]);
  or (_23075_, _23074_, _23065_);
  and (_23076_, _23075_, _07056_);
  and (_23078_, _07057_, \oc8051_golden_model_1.TCON [2]);
  or (_23079_, _23078_, _06160_);
  or (_23080_, _23079_, _23076_);
  and (_23081_, _23080_, _06157_);
  and (_23082_, _23081_, _23073_);
  and (_23083_, _11644_, \oc8051_golden_model_1.TCON [2]);
  and (_23084_, _14538_, _08407_);
  or (_23085_, _23084_, _23083_);
  and (_23086_, _23085_, _06156_);
  or (_23087_, _23086_, _06217_);
  or (_23088_, _23087_, _23082_);
  and (_23089_, _23088_, _23070_);
  or (_23090_, _23089_, _06220_);
  or (_23091_, _23075_, _06229_);
  and (_23092_, _23091_, _06153_);
  and (_23093_, _23092_, _23090_);
  and (_23094_, _14536_, _08407_);
  or (_23095_, _23094_, _23083_);
  and (_23096_, _23095_, _06152_);
  or (_23097_, _23096_, _06145_);
  or (_23099_, _23097_, _23093_);
  and (_23100_, _23084_, _14569_);
  or (_23101_, _23083_, _06146_);
  or (_23102_, _23101_, _23100_);
  and (_23103_, _23102_, _06140_);
  and (_23104_, _23103_, _23099_);
  and (_23105_, _14583_, _08407_);
  or (_23106_, _23105_, _23083_);
  and (_23107_, _23106_, _06139_);
  or (_23108_, _23107_, _09842_);
  or (_23109_, _23108_, _23104_);
  and (_23110_, _23109_, _23069_);
  or (_23111_, _23110_, _06116_);
  and (_23112_, _09211_, _07788_);
  or (_23113_, _23065_, _06117_);
  or (_23114_, _23113_, _23112_);
  and (_23115_, _23114_, _06114_);
  and (_23116_, _23115_, _23111_);
  and (_23117_, _14630_, _07788_);
  or (_23118_, _23065_, _23117_);
  and (_23120_, _23118_, _05787_);
  or (_23121_, _23120_, _23116_);
  or (_23122_, _23121_, _11136_);
  and (_23123_, _14646_, _07788_);
  or (_23124_, _23065_, _07127_);
  or (_23125_, _23124_, _23123_);
  and (_23126_, _07788_, _08768_);
  or (_23127_, _23126_, _23065_);
  or (_23128_, _23127_, _06111_);
  and (_23129_, _23128_, _07125_);
  and (_23131_, _23129_, _23125_);
  and (_23132_, _23131_, _23122_);
  and (_23133_, _10282_, _07788_);
  or (_23134_, _23133_, _23065_);
  and (_23135_, _23134_, _06402_);
  or (_23136_, _23135_, _23132_);
  and (_23137_, _23136_, _07132_);
  or (_23138_, _23065_, _08248_);
  and (_23139_, _23127_, _06306_);
  and (_23140_, _23139_, _23138_);
  or (_23141_, _23140_, _23137_);
  and (_23142_, _23141_, _07130_);
  and (_23143_, _23075_, _06411_);
  and (_23144_, _23143_, _23138_);
  or (_23145_, _23144_, _06303_);
  or (_23146_, _23145_, _23142_);
  and (_23147_, _14643_, _07788_);
  or (_23148_, _23065_, _08819_);
  or (_23149_, _23148_, _23147_);
  and (_23150_, _23149_, _08824_);
  and (_23152_, _23150_, _23146_);
  nor (_23153_, _10281_, _11639_);
  or (_23154_, _23153_, _23065_);
  and (_23155_, _23154_, _06396_);
  or (_23156_, _23155_, _06433_);
  or (_23157_, _23156_, _23152_);
  or (_23158_, _23072_, _06829_);
  and (_23159_, _23158_, _05749_);
  and (_23160_, _23159_, _23157_);
  and (_23161_, _23095_, _05748_);
  or (_23163_, _23161_, _06440_);
  or (_23164_, _23163_, _23160_);
  and (_23165_, _14710_, _07788_);
  or (_23166_, _23065_, _06444_);
  or (_23167_, _23166_, _23165_);
  and (_23168_, _23167_, _01317_);
  and (_23169_, _23168_, _23164_);
  or (_23170_, _23169_, _23064_);
  and (_43664_, _23170_, _43100_);
  and (_23171_, _01321_, \oc8051_golden_model_1.TCON [3]);
  and (_23172_, _11639_, \oc8051_golden_model_1.TCON [3]);
  and (_23173_, _07788_, _07544_);
  or (_23174_, _23173_, _23172_);
  or (_23175_, _23174_, _06132_);
  and (_23176_, _14738_, _07788_);
  or (_23177_, _23176_, _23172_);
  or (_23178_, _23177_, _06161_);
  and (_23179_, _07788_, \oc8051_golden_model_1.ACC [3]);
  or (_23180_, _23179_, _23172_);
  and (_23181_, _23180_, _07056_);
  and (_23182_, _07057_, \oc8051_golden_model_1.TCON [3]);
  or (_23183_, _23182_, _06160_);
  or (_23184_, _23183_, _23181_);
  and (_23185_, _23184_, _06157_);
  and (_23186_, _23185_, _23178_);
  and (_23187_, _11644_, \oc8051_golden_model_1.TCON [3]);
  and (_23188_, _14735_, _08407_);
  or (_23189_, _23188_, _23187_);
  and (_23190_, _23189_, _06156_);
  or (_23191_, _23190_, _06217_);
  or (_23194_, _23191_, _23186_);
  or (_23195_, _23174_, _07075_);
  and (_23196_, _23195_, _23194_);
  or (_23197_, _23196_, _06220_);
  or (_23198_, _23180_, _06229_);
  and (_23199_, _23198_, _06153_);
  and (_23200_, _23199_, _23197_);
  and (_23201_, _14731_, _08407_);
  or (_23202_, _23201_, _23187_);
  and (_23203_, _23202_, _06152_);
  or (_23204_, _23203_, _06145_);
  or (_23205_, _23204_, _23200_);
  or (_23206_, _23187_, _14764_);
  and (_23207_, _23206_, _23189_);
  or (_23208_, _23207_, _06146_);
  and (_23209_, _23208_, _06140_);
  and (_23210_, _23209_, _23205_);
  and (_23211_, _14732_, _08407_);
  or (_23212_, _23211_, _23187_);
  and (_23213_, _23212_, _06139_);
  or (_23215_, _23213_, _09842_);
  or (_23216_, _23215_, _23210_);
  and (_23217_, _23216_, _23175_);
  or (_23218_, _23217_, _06116_);
  and (_23219_, _09210_, _07788_);
  or (_23220_, _23172_, _06117_);
  or (_23221_, _23220_, _23219_);
  and (_23222_, _23221_, _06114_);
  and (_23223_, _23222_, _23218_);
  and (_23224_, _14825_, _07788_);
  or (_23226_, _23172_, _23224_);
  and (_23227_, _23226_, _05787_);
  or (_23228_, _23227_, _23223_);
  or (_23229_, _23228_, _11136_);
  and (_23230_, _14727_, _07788_);
  or (_23231_, _23172_, _07127_);
  or (_23232_, _23231_, _23230_);
  and (_23233_, _07788_, _08712_);
  or (_23234_, _23233_, _23172_);
  or (_23235_, _23234_, _06111_);
  and (_23236_, _23235_, _07125_);
  and (_23237_, _23236_, _23232_);
  and (_23238_, _23237_, _23229_);
  and (_23239_, _12318_, _07788_);
  or (_23240_, _23239_, _23172_);
  and (_23241_, _23240_, _06402_);
  or (_23242_, _23241_, _23238_);
  and (_23243_, _23242_, _07132_);
  or (_23244_, _23172_, _08140_);
  and (_23245_, _23234_, _06306_);
  and (_23247_, _23245_, _23244_);
  or (_23248_, _23247_, _23243_);
  and (_23249_, _23248_, _07130_);
  and (_23250_, _23180_, _06411_);
  and (_23251_, _23250_, _23244_);
  or (_23252_, _23251_, _06303_);
  or (_23253_, _23252_, _23249_);
  and (_23254_, _14724_, _07788_);
  or (_23255_, _23172_, _08819_);
  or (_23256_, _23255_, _23254_);
  and (_23258_, _23256_, _08824_);
  and (_23259_, _23258_, _23253_);
  nor (_23260_, _10273_, _11639_);
  or (_23261_, _23260_, _23172_);
  and (_23262_, _23261_, _06396_);
  or (_23263_, _23262_, _06433_);
  or (_23264_, _23263_, _23259_);
  or (_23265_, _23177_, _06829_);
  and (_23266_, _23265_, _05749_);
  and (_23267_, _23266_, _23264_);
  and (_23268_, _23202_, _05748_);
  or (_23269_, _23268_, _06440_);
  or (_23270_, _23269_, _23267_);
  and (_23271_, _14897_, _07788_);
  or (_23272_, _23172_, _06444_);
  or (_23273_, _23272_, _23271_);
  and (_23274_, _23273_, _01317_);
  and (_23275_, _23274_, _23270_);
  or (_23276_, _23275_, _23171_);
  and (_43665_, _23276_, _43100_);
  and (_23278_, _01321_, \oc8051_golden_model_1.TCON [4]);
  and (_23279_, _11639_, \oc8051_golden_model_1.TCON [4]);
  and (_23280_, _08336_, _07788_);
  or (_23281_, _23280_, _23279_);
  or (_23282_, _23281_, _06132_);
  and (_23283_, _11644_, \oc8051_golden_model_1.TCON [4]);
  and (_23284_, _14942_, _08407_);
  or (_23285_, _23284_, _23283_);
  and (_23286_, _23285_, _06152_);
  and (_23287_, _14928_, _07788_);
  or (_23289_, _23287_, _23279_);
  or (_23290_, _23289_, _06161_);
  and (_23291_, _07788_, \oc8051_golden_model_1.ACC [4]);
  or (_23292_, _23291_, _23279_);
  and (_23293_, _23292_, _07056_);
  and (_23294_, _07057_, \oc8051_golden_model_1.TCON [4]);
  or (_23295_, _23294_, _06160_);
  or (_23296_, _23295_, _23293_);
  and (_23297_, _23296_, _06157_);
  and (_23298_, _23297_, _23290_);
  and (_23299_, _14932_, _08407_);
  or (_23300_, _23299_, _23283_);
  and (_23301_, _23300_, _06156_);
  or (_23302_, _23301_, _06217_);
  or (_23303_, _23302_, _23298_);
  or (_23304_, _23281_, _07075_);
  and (_23305_, _23304_, _23303_);
  or (_23306_, _23305_, _06220_);
  or (_23307_, _23292_, _06229_);
  and (_23308_, _23307_, _06153_);
  and (_23310_, _23308_, _23306_);
  or (_23311_, _23310_, _23286_);
  and (_23312_, _23311_, _06146_);
  and (_23313_, _14950_, _08407_);
  or (_23314_, _23313_, _23283_);
  and (_23315_, _23314_, _06145_);
  or (_23316_, _23315_, _23312_);
  and (_23317_, _23316_, _06140_);
  and (_23318_, _14966_, _08407_);
  or (_23319_, _23318_, _23283_);
  and (_23321_, _23319_, _06139_);
  or (_23322_, _23321_, _09842_);
  or (_23323_, _23322_, _23317_);
  and (_23324_, _23323_, _23282_);
  or (_23325_, _23324_, _06116_);
  and (_23326_, _09209_, _07788_);
  or (_23327_, _23279_, _06117_);
  or (_23328_, _23327_, _23326_);
  and (_23329_, _23328_, _06114_);
  and (_23330_, _23329_, _23325_);
  and (_23331_, _15013_, _07788_);
  or (_23332_, _23331_, _23279_);
  and (_23333_, _23332_, _05787_);
  or (_23334_, _23333_, _11136_);
  or (_23335_, _23334_, _23330_);
  and (_23336_, _15029_, _07788_);
  or (_23337_, _23279_, _07127_);
  or (_23338_, _23337_, _23336_);
  and (_23339_, _08715_, _07788_);
  or (_23340_, _23339_, _23279_);
  or (_23342_, _23340_, _06111_);
  and (_23343_, _23342_, _07125_);
  and (_23344_, _23343_, _23338_);
  and (_23345_, _23344_, _23335_);
  and (_23346_, _10289_, _07788_);
  or (_23347_, _23346_, _23279_);
  and (_23348_, _23347_, _06402_);
  or (_23349_, _23348_, _23345_);
  and (_23350_, _23349_, _07132_);
  or (_23351_, _23279_, _08339_);
  and (_23353_, _23340_, _06306_);
  and (_23354_, _23353_, _23351_);
  or (_23355_, _23354_, _23350_);
  and (_23356_, _23355_, _07130_);
  and (_23357_, _23292_, _06411_);
  and (_23358_, _23357_, _23351_);
  or (_23359_, _23358_, _06303_);
  or (_23360_, _23359_, _23356_);
  and (_23361_, _15026_, _07788_);
  or (_23362_, _23279_, _08819_);
  or (_23363_, _23362_, _23361_);
  and (_23364_, _23363_, _08824_);
  and (_23365_, _23364_, _23360_);
  nor (_23366_, _10288_, _11639_);
  or (_23367_, _23366_, _23279_);
  and (_23368_, _23367_, _06396_);
  or (_23369_, _23368_, _06433_);
  or (_23370_, _23369_, _23365_);
  or (_23371_, _23289_, _06829_);
  and (_23372_, _23371_, _05749_);
  and (_23374_, _23372_, _23370_);
  and (_23375_, _23285_, _05748_);
  or (_23376_, _23375_, _06440_);
  or (_23377_, _23376_, _23374_);
  and (_23378_, _15087_, _07788_);
  or (_23379_, _23279_, _06444_);
  or (_23380_, _23379_, _23378_);
  and (_23381_, _23380_, _01317_);
  and (_23382_, _23381_, _23377_);
  or (_23383_, _23382_, _23278_);
  and (_43666_, _23383_, _43100_);
  and (_23385_, _01321_, \oc8051_golden_model_1.TCON [5]);
  and (_23386_, _11639_, \oc8051_golden_model_1.TCON [5]);
  and (_23387_, _15119_, _07788_);
  or (_23388_, _23387_, _23386_);
  or (_23389_, _23388_, _06161_);
  and (_23390_, _07788_, \oc8051_golden_model_1.ACC [5]);
  or (_23391_, _23390_, _23386_);
  and (_23392_, _23391_, _07056_);
  and (_23393_, _07057_, \oc8051_golden_model_1.TCON [5]);
  or (_23394_, _23393_, _06160_);
  or (_23395_, _23394_, _23392_);
  and (_23396_, _23395_, _06157_);
  and (_23397_, _23396_, _23389_);
  and (_23398_, _11644_, \oc8051_golden_model_1.TCON [5]);
  and (_23399_, _15123_, _08407_);
  or (_23400_, _23399_, _23398_);
  and (_23401_, _23400_, _06156_);
  or (_23402_, _23401_, _06217_);
  or (_23403_, _23402_, _23397_);
  and (_23405_, _08101_, _07788_);
  or (_23406_, _23405_, _23386_);
  or (_23407_, _23406_, _07075_);
  and (_23408_, _23407_, _23403_);
  or (_23409_, _23408_, _06220_);
  or (_23410_, _23391_, _06229_);
  and (_23411_, _23410_, _06153_);
  and (_23412_, _23411_, _23409_);
  and (_23413_, _15104_, _08407_);
  or (_23414_, _23413_, _23398_);
  and (_23416_, _23414_, _06152_);
  or (_23417_, _23416_, _06145_);
  or (_23418_, _23417_, _23412_);
  or (_23419_, _23398_, _15138_);
  and (_23420_, _23419_, _23400_);
  or (_23421_, _23420_, _06146_);
  and (_23422_, _23421_, _06140_);
  and (_23423_, _23422_, _23418_);
  and (_23424_, _15155_, _08407_);
  or (_23425_, _23424_, _23398_);
  and (_23426_, _23425_, _06139_);
  or (_23427_, _23426_, _09842_);
  or (_23428_, _23427_, _23423_);
  or (_23429_, _23406_, _06132_);
  and (_23430_, _23429_, _23428_);
  or (_23431_, _23430_, _06116_);
  and (_23432_, _09208_, _07788_);
  or (_23433_, _23386_, _06117_);
  or (_23434_, _23433_, _23432_);
  and (_23435_, _23434_, _06114_);
  and (_23437_, _23435_, _23431_);
  and (_23438_, _15203_, _07788_);
  or (_23439_, _23438_, _23386_);
  and (_23440_, _23439_, _05787_);
  or (_23441_, _23440_, _11136_);
  or (_23442_, _23441_, _23437_);
  and (_23443_, _15219_, _07788_);
  or (_23444_, _23386_, _07127_);
  or (_23445_, _23444_, _23443_);
  and (_23446_, _08736_, _07788_);
  or (_23448_, _23446_, _23386_);
  or (_23449_, _23448_, _06111_);
  and (_23450_, _23449_, _07125_);
  and (_23451_, _23450_, _23445_);
  and (_23452_, _23451_, _23442_);
  and (_23453_, _12325_, _07788_);
  or (_23454_, _23453_, _23386_);
  and (_23455_, _23454_, _06402_);
  or (_23456_, _23455_, _23452_);
  and (_23457_, _23456_, _07132_);
  or (_23458_, _23386_, _08104_);
  and (_23459_, _23448_, _06306_);
  and (_23460_, _23459_, _23458_);
  or (_23461_, _23460_, _23457_);
  and (_23462_, _23461_, _07130_);
  and (_23463_, _23391_, _06411_);
  and (_23464_, _23463_, _23458_);
  or (_23465_, _23464_, _06303_);
  or (_23466_, _23465_, _23462_);
  and (_23467_, _15216_, _07788_);
  or (_23469_, _23386_, _08819_);
  or (_23470_, _23469_, _23467_);
  and (_23471_, _23470_, _08824_);
  and (_23472_, _23471_, _23466_);
  nor (_23473_, _10269_, _11639_);
  or (_23474_, _23473_, _23386_);
  and (_23475_, _23474_, _06396_);
  or (_23476_, _23475_, _06433_);
  or (_23477_, _23476_, _23472_);
  or (_23478_, _23388_, _06829_);
  and (_23480_, _23478_, _05749_);
  and (_23481_, _23480_, _23477_);
  and (_23482_, _23414_, _05748_);
  or (_23483_, _23482_, _06440_);
  or (_23484_, _23483_, _23481_);
  and (_23485_, _15275_, _07788_);
  or (_23486_, _23386_, _06444_);
  or (_23487_, _23486_, _23485_);
  and (_23488_, _23487_, _01317_);
  and (_23489_, _23488_, _23484_);
  or (_23491_, _23489_, _23385_);
  and (_43667_, _23491_, _43100_);
  and (_23492_, _01321_, \oc8051_golden_model_1.TCON [6]);
  and (_23493_, _11639_, \oc8051_golden_model_1.TCON [6]);
  and (_23494_, _15300_, _07788_);
  or (_23495_, _23494_, _23493_);
  or (_23496_, _23495_, _06161_);
  and (_23497_, _07788_, \oc8051_golden_model_1.ACC [6]);
  or (_23498_, _23497_, _23493_);
  and (_23499_, _23498_, _07056_);
  and (_23500_, _07057_, \oc8051_golden_model_1.TCON [6]);
  or (_23501_, _23500_, _06160_);
  or (_23502_, _23501_, _23499_);
  and (_23503_, _23502_, _06157_);
  and (_23504_, _23503_, _23496_);
  and (_23505_, _11644_, \oc8051_golden_model_1.TCON [6]);
  and (_23506_, _15316_, _08407_);
  or (_23507_, _23506_, _23505_);
  and (_23508_, _23507_, _06156_);
  or (_23509_, _23508_, _06217_);
  or (_23511_, _23509_, _23504_);
  and (_23512_, _08012_, _07788_);
  or (_23513_, _23512_, _23493_);
  or (_23514_, _23513_, _07075_);
  and (_23515_, _23514_, _23511_);
  or (_23516_, _23515_, _06220_);
  or (_23517_, _23498_, _06229_);
  and (_23518_, _23517_, _06153_);
  and (_23519_, _23518_, _23516_);
  and (_23520_, _15297_, _08407_);
  or (_23522_, _23520_, _23505_);
  and (_23523_, _23522_, _06152_);
  or (_23524_, _23523_, _06145_);
  or (_23525_, _23524_, _23519_);
  or (_23526_, _23505_, _15331_);
  and (_23527_, _23526_, _23507_);
  or (_23528_, _23527_, _06146_);
  and (_23529_, _23528_, _06140_);
  and (_23530_, _23529_, _23525_);
  and (_23531_, _15348_, _08407_);
  or (_23533_, _23531_, _23505_);
  and (_23534_, _23533_, _06139_);
  or (_23535_, _23534_, _09842_);
  or (_23536_, _23535_, _23530_);
  or (_23537_, _23513_, _06132_);
  and (_23538_, _23537_, _23536_);
  or (_23539_, _23538_, _06116_);
  and (_23540_, _09207_, _07788_);
  or (_23541_, _23493_, _06117_);
  or (_23542_, _23541_, _23540_);
  and (_23543_, _23542_, _06114_);
  and (_23544_, _23543_, _23539_);
  and (_23545_, _15395_, _07788_);
  or (_23546_, _23545_, _23493_);
  and (_23547_, _23546_, _05787_);
  or (_23548_, _23547_, _11136_);
  or (_23549_, _23548_, _23544_);
  and (_23550_, _15413_, _07788_);
  or (_23551_, _23493_, _07127_);
  or (_23552_, _23551_, _23550_);
  and (_23554_, _15402_, _07788_);
  or (_23555_, _23554_, _23493_);
  or (_23556_, _23555_, _06111_);
  and (_23557_, _23556_, _07125_);
  and (_23558_, _23557_, _23552_);
  and (_23559_, _23558_, _23549_);
  and (_23560_, _10295_, _07788_);
  or (_23561_, _23560_, _23493_);
  and (_23562_, _23561_, _06402_);
  or (_23563_, _23562_, _23559_);
  and (_23565_, _23563_, _07132_);
  or (_23566_, _23493_, _08015_);
  and (_23567_, _23555_, _06306_);
  and (_23568_, _23567_, _23566_);
  or (_23569_, _23568_, _23565_);
  and (_23570_, _23569_, _07130_);
  and (_23571_, _23498_, _06411_);
  and (_23572_, _23571_, _23566_);
  or (_23573_, _23572_, _06303_);
  or (_23574_, _23573_, _23570_);
  and (_23575_, _15410_, _07788_);
  or (_23576_, _23493_, _08819_);
  or (_23577_, _23576_, _23575_);
  and (_23578_, _23577_, _08824_);
  and (_23579_, _23578_, _23574_);
  nor (_23580_, _10294_, _11639_);
  or (_23581_, _23580_, _23493_);
  and (_23582_, _23581_, _06396_);
  or (_23583_, _23582_, _06433_);
  or (_23584_, _23583_, _23579_);
  or (_23586_, _23495_, _06829_);
  and (_23587_, _23586_, _05749_);
  and (_23588_, _23587_, _23584_);
  and (_23589_, _23522_, _05748_);
  or (_23590_, _23589_, _06440_);
  or (_23591_, _23590_, _23588_);
  and (_23592_, _15478_, _07788_);
  or (_23593_, _23493_, _06444_);
  or (_23594_, _23593_, _23592_);
  and (_23595_, _23594_, _01317_);
  and (_23597_, _23595_, _23591_);
  or (_23598_, _23597_, _23492_);
  and (_43668_, _23598_, _43100_);
  not (_23599_, \oc8051_golden_model_1.TH1 [0]);
  nor (_23600_, _01317_, _23599_);
  nand (_23601_, _10276_, _07817_);
  nor (_23602_, _07817_, _23599_);
  nor (_23603_, _23602_, _07130_);
  nand (_23604_, _23603_, _23601_);
  nor (_23605_, _08211_, _11740_);
  or (_23607_, _23605_, _23602_);
  or (_23608_, _23607_, _06161_);
  and (_23609_, _07817_, \oc8051_golden_model_1.ACC [0]);
  or (_23610_, _23609_, _23602_);
  and (_23611_, _23610_, _07056_);
  nor (_23612_, _07056_, _23599_);
  or (_23613_, _23612_, _06160_);
  or (_23614_, _23613_, _23611_);
  and (_23615_, _23614_, _07075_);
  and (_23616_, _23615_, _23608_);
  and (_23618_, _07817_, _07049_);
  or (_23619_, _23618_, _23602_);
  and (_23620_, _23619_, _06217_);
  or (_23621_, _23620_, _23616_);
  and (_23622_, _23621_, _06229_);
  and (_23623_, _23610_, _06220_);
  or (_23624_, _23623_, _09842_);
  or (_23625_, _23624_, _23622_);
  or (_23626_, _23619_, _06132_);
  and (_23627_, _23626_, _23625_);
  or (_23629_, _23627_, _06116_);
  and (_23630_, _09160_, _07817_);
  or (_23631_, _23602_, _06117_);
  or (_23632_, _23631_, _23630_);
  and (_23633_, _23632_, _23629_);
  or (_23634_, _23633_, _05787_);
  and (_23635_, _14260_, _07817_);
  or (_23636_, _23635_, _23602_);
  or (_23637_, _23636_, _06114_);
  and (_23638_, _23637_, _06111_);
  and (_23640_, _23638_, _23634_);
  and (_23641_, _07817_, _08708_);
  or (_23642_, _23641_, _23602_);
  and (_23643_, _23642_, _06110_);
  or (_23644_, _23643_, _06297_);
  or (_23645_, _23644_, _23640_);
  and (_23646_, _14275_, _07817_);
  or (_23647_, _23602_, _07127_);
  or (_23648_, _23647_, _23646_);
  and (_23649_, _23648_, _07125_);
  and (_23651_, _23649_, _23645_);
  nor (_23652_, _12321_, _11740_);
  or (_23653_, _23652_, _23602_);
  and (_23654_, _23601_, _06402_);
  and (_23655_, _23654_, _23653_);
  or (_23656_, _23655_, _23651_);
  and (_23657_, _23656_, _07132_);
  nand (_23658_, _23642_, _06306_);
  nor (_23659_, _23658_, _23605_);
  or (_23660_, _23659_, _06411_);
  or (_23662_, _23660_, _23657_);
  and (_23663_, _23662_, _23604_);
  or (_23664_, _23663_, _06303_);
  and (_23665_, _14167_, _07817_);
  or (_23666_, _23602_, _08819_);
  or (_23667_, _23666_, _23665_);
  and (_23668_, _23667_, _08824_);
  and (_23669_, _23668_, _23664_);
  and (_23670_, _23653_, _06396_);
  or (_23671_, _23670_, _19287_);
  or (_23673_, _23671_, _23669_);
  or (_23674_, _23607_, _06630_);
  and (_23675_, _23674_, _01317_);
  and (_23676_, _23675_, _23673_);
  or (_23677_, _23676_, _23600_);
  and (_43670_, _23677_, _43100_);
  not (_23678_, \oc8051_golden_model_1.TH1 [1]);
  nor (_23679_, _01317_, _23678_);
  or (_23680_, _14442_, _11740_);
  or (_23681_, _07817_, \oc8051_golden_model_1.TH1 [1]);
  and (_23682_, _23681_, _05787_);
  and (_23683_, _23682_, _23680_);
  nor (_23684_, _07817_, _23678_);
  and (_23685_, _07817_, _07306_);
  or (_23686_, _23685_, _23684_);
  or (_23687_, _23686_, _06132_);
  and (_23688_, _07817_, \oc8051_golden_model_1.ACC [1]);
  or (_23689_, _23688_, _23684_);
  and (_23690_, _23689_, _06220_);
  or (_23691_, _23690_, _09842_);
  and (_23692_, _14363_, _07817_);
  not (_23693_, _23692_);
  and (_23694_, _23693_, _23681_);
  and (_23695_, _23694_, _06160_);
  nor (_23696_, _07056_, _23678_);
  and (_23697_, _23689_, _07056_);
  or (_23698_, _23697_, _23696_);
  and (_23699_, _23698_, _06161_);
  or (_23700_, _23699_, _06217_);
  or (_23701_, _23700_, _23695_);
  or (_23703_, _23686_, _07075_);
  and (_23704_, _23703_, _06229_);
  and (_23705_, _23704_, _23701_);
  or (_23706_, _23705_, _23691_);
  and (_23707_, _23706_, _23687_);
  or (_23708_, _23707_, _06116_);
  and (_23709_, _23708_, _06114_);
  and (_23710_, _09115_, _07817_);
  or (_23711_, _23684_, _06117_);
  or (_23712_, _23711_, _23710_);
  and (_23714_, _23712_, _23709_);
  or (_23715_, _23714_, _23683_);
  and (_23716_, _23715_, _06298_);
  or (_23717_, _14346_, _11740_);
  and (_23718_, _23717_, _06297_);
  nand (_23719_, _07817_, _06945_);
  and (_23720_, _23719_, _06110_);
  or (_23721_, _23720_, _23718_);
  and (_23722_, _23721_, _23681_);
  or (_23723_, _23722_, _06402_);
  or (_23725_, _23723_, _23716_);
  nor (_23726_, _10277_, _11740_);
  or (_23727_, _23726_, _23684_);
  nand (_23728_, _10275_, _07817_);
  and (_23729_, _23728_, _23727_);
  or (_23730_, _23729_, _07125_);
  and (_23731_, _23730_, _07132_);
  and (_23732_, _23731_, _23725_);
  or (_23733_, _14344_, _11740_);
  and (_23734_, _23681_, _06306_);
  and (_23736_, _23734_, _23733_);
  or (_23737_, _23736_, _06411_);
  or (_23738_, _23737_, _23732_);
  nor (_23739_, _23684_, _07130_);
  nand (_23740_, _23739_, _23728_);
  and (_23741_, _23740_, _08819_);
  and (_23742_, _23741_, _23738_);
  or (_23743_, _23719_, _08176_);
  and (_23744_, _23681_, _06303_);
  and (_23745_, _23744_, _23743_);
  or (_23747_, _23745_, _06396_);
  or (_23748_, _23747_, _23742_);
  or (_23749_, _23727_, _08824_);
  and (_23750_, _23749_, _06829_);
  and (_23751_, _23750_, _23748_);
  and (_23752_, _23694_, _06433_);
  or (_23753_, _23752_, _06440_);
  or (_23754_, _23753_, _23751_);
  or (_23755_, _23684_, _06444_);
  or (_23756_, _23755_, _23692_);
  and (_23758_, _23756_, _01317_);
  and (_23759_, _23758_, _23754_);
  or (_23760_, _23759_, _23679_);
  and (_43671_, _23760_, _43100_);
  and (_23761_, _01321_, \oc8051_golden_model_1.TH1 [2]);
  and (_23762_, _11740_, \oc8051_golden_model_1.TH1 [2]);
  or (_23763_, _23762_, _08248_);
  and (_23764_, _07817_, _08768_);
  or (_23765_, _23764_, _23762_);
  and (_23766_, _23765_, _06306_);
  and (_23768_, _23766_, _23763_);
  and (_23769_, _09211_, _07817_);
  or (_23770_, _23769_, _23762_);
  and (_23771_, _23770_, _06116_);
  and (_23772_, _14542_, _07817_);
  or (_23773_, _23772_, _23762_);
  or (_23774_, _23773_, _06161_);
  and (_23775_, _07817_, \oc8051_golden_model_1.ACC [2]);
  or (_23776_, _23775_, _23762_);
  and (_23777_, _23776_, _07056_);
  and (_23779_, _07057_, \oc8051_golden_model_1.TH1 [2]);
  or (_23780_, _23779_, _06160_);
  or (_23781_, _23780_, _23777_);
  and (_23782_, _23781_, _07075_);
  and (_23783_, _23782_, _23774_);
  and (_23784_, _07817_, _07708_);
  or (_23785_, _23784_, _23762_);
  and (_23786_, _23785_, _06217_);
  or (_23787_, _23786_, _23783_);
  and (_23788_, _23787_, _06229_);
  and (_23790_, _23776_, _06220_);
  or (_23791_, _23790_, _09842_);
  or (_23792_, _23791_, _23788_);
  or (_23793_, _23785_, _06132_);
  and (_23794_, _23793_, _06117_);
  and (_23795_, _23794_, _23792_);
  or (_23796_, _23795_, _05787_);
  or (_23797_, _23796_, _23771_);
  and (_23798_, _14630_, _07817_);
  or (_23799_, _23798_, _23762_);
  or (_23801_, _23799_, _06114_);
  and (_23802_, _23801_, _06111_);
  and (_23803_, _23802_, _23797_);
  and (_23804_, _23765_, _06110_);
  or (_23805_, _23804_, _06297_);
  or (_23806_, _23805_, _23803_);
  and (_23807_, _14646_, _07817_);
  or (_23808_, _23762_, _07127_);
  or (_23809_, _23808_, _23807_);
  and (_23810_, _23809_, _07125_);
  and (_23812_, _23810_, _23806_);
  and (_23813_, _10282_, _07817_);
  or (_23814_, _23813_, _23762_);
  and (_23815_, _23814_, _06402_);
  or (_23816_, _23815_, _23812_);
  and (_23817_, _23816_, _07132_);
  or (_23818_, _23817_, _23768_);
  and (_23819_, _23818_, _07130_);
  and (_23820_, _23776_, _06411_);
  and (_23821_, _23820_, _23763_);
  or (_23823_, _23821_, _06303_);
  or (_23824_, _23823_, _23819_);
  and (_23825_, _14643_, _07817_);
  or (_23826_, _23762_, _08819_);
  or (_23827_, _23826_, _23825_);
  and (_23828_, _23827_, _08824_);
  and (_23829_, _23828_, _23824_);
  nor (_23830_, _10281_, _11740_);
  or (_23831_, _23830_, _23762_);
  and (_23832_, _23831_, _06396_);
  or (_23834_, _23832_, _23829_);
  and (_23835_, _23834_, _06829_);
  and (_23836_, _23773_, _06433_);
  or (_23837_, _23836_, _06440_);
  or (_23838_, _23837_, _23835_);
  and (_23839_, _14710_, _07817_);
  or (_23840_, _23762_, _06444_);
  or (_23841_, _23840_, _23839_);
  and (_23842_, _23841_, _01317_);
  and (_23843_, _23842_, _23838_);
  or (_23845_, _23843_, _23761_);
  and (_43672_, _23845_, _43100_);
  and (_23846_, _11740_, \oc8051_golden_model_1.TH1 [3]);
  and (_23847_, _14738_, _07817_);
  or (_23848_, _23847_, _23846_);
  or (_23849_, _23848_, _06161_);
  and (_23850_, _07817_, \oc8051_golden_model_1.ACC [3]);
  or (_23851_, _23850_, _23846_);
  and (_23852_, _23851_, _07056_);
  and (_23853_, _07057_, \oc8051_golden_model_1.TH1 [3]);
  or (_23855_, _23853_, _06160_);
  or (_23856_, _23855_, _23852_);
  and (_23857_, _23856_, _07075_);
  and (_23858_, _23857_, _23849_);
  and (_23859_, _07817_, _07544_);
  or (_23860_, _23859_, _23846_);
  and (_23861_, _23860_, _06217_);
  or (_23862_, _23861_, _23858_);
  and (_23863_, _23862_, _06229_);
  and (_23864_, _23851_, _06220_);
  or (_23866_, _23864_, _09842_);
  or (_23867_, _23866_, _23863_);
  or (_23868_, _23860_, _06132_);
  and (_23869_, _23868_, _06117_);
  and (_23870_, _23869_, _23867_);
  and (_23871_, _09210_, _07817_);
  or (_23872_, _23871_, _23846_);
  and (_23873_, _23872_, _06116_);
  or (_23874_, _23873_, _05787_);
  or (_23875_, _23874_, _23870_);
  and (_23877_, _14825_, _07817_);
  or (_23878_, _23846_, _06114_);
  or (_23879_, _23878_, _23877_);
  and (_23880_, _23879_, _06111_);
  and (_23881_, _23880_, _23875_);
  and (_23882_, _07817_, _08712_);
  or (_23883_, _23882_, _23846_);
  and (_23884_, _23883_, _06110_);
  or (_23885_, _23884_, _06297_);
  or (_23886_, _23885_, _23881_);
  and (_23887_, _14727_, _07817_);
  or (_23888_, _23887_, _23846_);
  or (_23889_, _23888_, _07127_);
  and (_23890_, _23889_, _07125_);
  and (_23891_, _23890_, _23886_);
  and (_23892_, _12318_, _07817_);
  or (_23893_, _23892_, _23846_);
  and (_23894_, _23893_, _06402_);
  or (_23895_, _23894_, _23891_);
  and (_23896_, _23895_, _07132_);
  or (_23899_, _23846_, _08140_);
  and (_23900_, _23883_, _06306_);
  and (_23901_, _23900_, _23899_);
  or (_23902_, _23901_, _23896_);
  and (_23903_, _23902_, _07130_);
  and (_23904_, _23851_, _06411_);
  and (_23905_, _23904_, _23899_);
  or (_23906_, _23905_, _06303_);
  or (_23907_, _23906_, _23903_);
  and (_23908_, _14724_, _07817_);
  or (_23910_, _23846_, _08819_);
  or (_23911_, _23910_, _23908_);
  and (_23912_, _23911_, _08824_);
  and (_23913_, _23912_, _23907_);
  nor (_23914_, _10273_, _11740_);
  or (_23915_, _23914_, _23846_);
  and (_23916_, _23915_, _06396_);
  or (_23917_, _23916_, _06433_);
  or (_23918_, _23917_, _23913_);
  or (_23919_, _23848_, _06829_);
  and (_23921_, _23919_, _06444_);
  and (_23922_, _23921_, _23918_);
  and (_23923_, _14897_, _07817_);
  or (_23924_, _23923_, _23846_);
  and (_23925_, _23924_, _06440_);
  or (_23926_, _23925_, _01321_);
  or (_23927_, _23926_, _23922_);
  or (_23928_, _01317_, \oc8051_golden_model_1.TH1 [3]);
  and (_23929_, _23928_, _43100_);
  and (_43673_, _23929_, _23927_);
  and (_23931_, _11740_, \oc8051_golden_model_1.TH1 [4]);
  and (_23932_, _14928_, _07817_);
  or (_23933_, _23932_, _23931_);
  or (_23934_, _23933_, _06161_);
  and (_23935_, _07817_, \oc8051_golden_model_1.ACC [4]);
  or (_23936_, _23935_, _23931_);
  and (_23937_, _23936_, _07056_);
  and (_23938_, _07057_, \oc8051_golden_model_1.TH1 [4]);
  or (_23939_, _23938_, _06160_);
  or (_23940_, _23939_, _23937_);
  and (_23942_, _23940_, _07075_);
  and (_23943_, _23942_, _23934_);
  and (_23944_, _08336_, _07817_);
  or (_23945_, _23944_, _23931_);
  and (_23946_, _23945_, _06217_);
  or (_23947_, _23946_, _23943_);
  and (_23948_, _23947_, _06229_);
  and (_23949_, _23936_, _06220_);
  or (_23950_, _23949_, _09842_);
  or (_23951_, _23950_, _23948_);
  or (_23953_, _23945_, _06132_);
  and (_23954_, _23953_, _23951_);
  or (_23955_, _23954_, _06116_);
  and (_23956_, _09209_, _07817_);
  or (_23957_, _23931_, _06117_);
  or (_23958_, _23957_, _23956_);
  and (_23959_, _23958_, _06114_);
  and (_23960_, _23959_, _23955_);
  and (_23961_, _15013_, _07817_);
  or (_23962_, _23961_, _23931_);
  and (_23964_, _23962_, _05787_);
  or (_23965_, _23964_, _23960_);
  or (_23966_, _23965_, _11136_);
  and (_23967_, _15029_, _07817_);
  or (_23968_, _23931_, _07127_);
  or (_23969_, _23968_, _23967_);
  and (_23970_, _08715_, _07817_);
  or (_23971_, _23970_, _23931_);
  or (_23972_, _23971_, _06111_);
  and (_23973_, _23972_, _07125_);
  and (_23975_, _23973_, _23969_);
  and (_23976_, _23975_, _23966_);
  and (_23977_, _10289_, _07817_);
  or (_23978_, _23977_, _23931_);
  and (_23979_, _23978_, _06402_);
  or (_23980_, _23979_, _23976_);
  and (_23981_, _23980_, _07132_);
  or (_23982_, _23931_, _08339_);
  and (_23983_, _23971_, _06306_);
  and (_23984_, _23983_, _23982_);
  or (_23986_, _23984_, _23981_);
  and (_23987_, _23986_, _07130_);
  and (_23988_, _23936_, _06411_);
  and (_23989_, _23988_, _23982_);
  or (_23990_, _23989_, _06303_);
  or (_23991_, _23990_, _23987_);
  and (_23992_, _15026_, _07817_);
  or (_23993_, _23931_, _08819_);
  or (_23994_, _23993_, _23992_);
  and (_23995_, _23994_, _08824_);
  and (_23997_, _23995_, _23991_);
  nor (_23998_, _10288_, _11740_);
  or (_23999_, _23998_, _23931_);
  and (_24000_, _23999_, _06396_);
  or (_24001_, _24000_, _06433_);
  or (_24002_, _24001_, _23997_);
  or (_24003_, _23933_, _06829_);
  and (_24004_, _24003_, _06444_);
  and (_24005_, _24004_, _24002_);
  and (_24006_, _15087_, _07817_);
  or (_24008_, _24006_, _23931_);
  and (_24009_, _24008_, _06440_);
  or (_24010_, _24009_, _01321_);
  or (_24011_, _24010_, _24005_);
  or (_24012_, _01317_, \oc8051_golden_model_1.TH1 [4]);
  and (_24013_, _24012_, _43100_);
  and (_43674_, _24013_, _24011_);
  and (_24014_, _11740_, \oc8051_golden_model_1.TH1 [5]);
  or (_24015_, _24014_, _08104_);
  and (_24016_, _08736_, _07817_);
  or (_24018_, _24016_, _24014_);
  and (_24019_, _24018_, _06306_);
  and (_24020_, _24019_, _24015_);
  and (_24021_, _15119_, _07817_);
  or (_24022_, _24021_, _24014_);
  or (_24023_, _24022_, _06161_);
  and (_24024_, _07817_, \oc8051_golden_model_1.ACC [5]);
  or (_24025_, _24024_, _24014_);
  and (_24026_, _24025_, _07056_);
  and (_24027_, _07057_, \oc8051_golden_model_1.TH1 [5]);
  or (_24029_, _24027_, _06160_);
  or (_24030_, _24029_, _24026_);
  and (_24031_, _24030_, _07075_);
  and (_24032_, _24031_, _24023_);
  and (_24033_, _08101_, _07817_);
  or (_24034_, _24033_, _24014_);
  and (_24035_, _24034_, _06217_);
  or (_24036_, _24035_, _24032_);
  and (_24037_, _24036_, _06229_);
  and (_24038_, _24025_, _06220_);
  or (_24040_, _24038_, _09842_);
  or (_24041_, _24040_, _24037_);
  or (_24042_, _24034_, _06132_);
  and (_24043_, _24042_, _24041_);
  or (_24044_, _24043_, _06116_);
  and (_24045_, _09208_, _07817_);
  or (_24046_, _24014_, _06117_);
  or (_24047_, _24046_, _24045_);
  and (_24048_, _24047_, _06114_);
  and (_24049_, _24048_, _24044_);
  and (_24051_, _15203_, _07817_);
  or (_24052_, _24051_, _24014_);
  and (_24053_, _24052_, _05787_);
  or (_24054_, _24053_, _11136_);
  or (_24055_, _24054_, _24049_);
  and (_24056_, _15219_, _07817_);
  or (_24057_, _24014_, _07127_);
  or (_24058_, _24057_, _24056_);
  or (_24059_, _24018_, _06111_);
  and (_24060_, _24059_, _07125_);
  and (_24062_, _24060_, _24058_);
  and (_24063_, _24062_, _24055_);
  and (_24064_, _12325_, _07817_);
  or (_24065_, _24064_, _24014_);
  and (_24066_, _24065_, _06402_);
  or (_24067_, _24066_, _24063_);
  and (_24068_, _24067_, _07132_);
  or (_24069_, _24068_, _24020_);
  and (_24070_, _24069_, _07130_);
  and (_24071_, _24025_, _06411_);
  and (_24072_, _24071_, _24015_);
  or (_24073_, _24072_, _06303_);
  or (_24074_, _24073_, _24070_);
  and (_24075_, _15216_, _07817_);
  or (_24076_, _24014_, _08819_);
  or (_24077_, _24076_, _24075_);
  and (_24078_, _24077_, _08824_);
  and (_24079_, _24078_, _24074_);
  nor (_24080_, _10269_, _11740_);
  or (_24081_, _24080_, _24014_);
  and (_24084_, _24081_, _06396_);
  or (_24085_, _24084_, _06433_);
  or (_24086_, _24085_, _24079_);
  or (_24087_, _24022_, _06829_);
  and (_24088_, _24087_, _06444_);
  and (_24089_, _24088_, _24086_);
  and (_24090_, _15275_, _07817_);
  or (_24091_, _24090_, _24014_);
  and (_24092_, _24091_, _06440_);
  or (_24093_, _24092_, _01321_);
  or (_24095_, _24093_, _24089_);
  or (_24096_, _01317_, \oc8051_golden_model_1.TH1 [5]);
  and (_24097_, _24096_, _43100_);
  and (_43675_, _24097_, _24095_);
  and (_24098_, _11740_, \oc8051_golden_model_1.TH1 [6]);
  and (_24099_, _15300_, _07817_);
  or (_24100_, _24099_, _24098_);
  or (_24101_, _24100_, _06161_);
  and (_24102_, _07817_, \oc8051_golden_model_1.ACC [6]);
  or (_24103_, _24102_, _24098_);
  and (_24105_, _24103_, _07056_);
  and (_24106_, _07057_, \oc8051_golden_model_1.TH1 [6]);
  or (_24107_, _24106_, _06160_);
  or (_24108_, _24107_, _24105_);
  and (_24109_, _24108_, _07075_);
  and (_24110_, _24109_, _24101_);
  and (_24111_, _08012_, _07817_);
  or (_24112_, _24111_, _24098_);
  and (_24113_, _24112_, _06217_);
  or (_24114_, _24113_, _24110_);
  and (_24116_, _24114_, _06229_);
  and (_24117_, _24103_, _06220_);
  or (_24118_, _24117_, _09842_);
  or (_24119_, _24118_, _24116_);
  or (_24120_, _24112_, _06132_);
  and (_24121_, _24120_, _24119_);
  or (_24122_, _24121_, _06116_);
  and (_24123_, _09207_, _07817_);
  or (_24124_, _24098_, _06117_);
  or (_24125_, _24124_, _24123_);
  and (_24127_, _24125_, _06114_);
  and (_24128_, _24127_, _24122_);
  and (_24129_, _15395_, _07817_);
  or (_24130_, _24129_, _24098_);
  and (_24131_, _24130_, _05787_);
  or (_24132_, _24131_, _11136_);
  or (_24133_, _24132_, _24128_);
  and (_24134_, _15413_, _07817_);
  or (_24135_, _24098_, _07127_);
  or (_24136_, _24135_, _24134_);
  and (_24138_, _15402_, _07817_);
  or (_24139_, _24138_, _24098_);
  or (_24140_, _24139_, _06111_);
  and (_24141_, _24140_, _07125_);
  and (_24142_, _24141_, _24136_);
  and (_24143_, _24142_, _24133_);
  and (_24144_, _10295_, _07817_);
  or (_24145_, _24144_, _24098_);
  and (_24146_, _24145_, _06402_);
  or (_24147_, _24146_, _24143_);
  and (_24149_, _24147_, _07132_);
  or (_24150_, _24098_, _08015_);
  and (_24151_, _24139_, _06306_);
  and (_24152_, _24151_, _24150_);
  or (_24153_, _24152_, _24149_);
  and (_24154_, _24153_, _07130_);
  and (_24155_, _24103_, _06411_);
  and (_24156_, _24155_, _24150_);
  or (_24157_, _24156_, _06303_);
  or (_24158_, _24157_, _24154_);
  and (_24160_, _15410_, _07817_);
  or (_24161_, _24098_, _08819_);
  or (_24162_, _24161_, _24160_);
  and (_24163_, _24162_, _08824_);
  and (_24164_, _24163_, _24158_);
  nor (_24165_, _10294_, _11740_);
  or (_24166_, _24165_, _24098_);
  and (_24167_, _24166_, _06396_);
  or (_24168_, _24167_, _06433_);
  or (_24169_, _24168_, _24164_);
  or (_24171_, _24100_, _06829_);
  and (_24172_, _24171_, _06444_);
  and (_24173_, _24172_, _24169_);
  and (_24174_, _15478_, _07817_);
  or (_24175_, _24174_, _24098_);
  and (_24176_, _24175_, _06440_);
  or (_24177_, _24176_, _01321_);
  or (_24178_, _24177_, _24173_);
  or (_24179_, _01317_, \oc8051_golden_model_1.TH1 [6]);
  and (_24180_, _24179_, _43100_);
  and (_43676_, _24180_, _24178_);
  not (_24182_, \oc8051_golden_model_1.TH0 [0]);
  nor (_24183_, _01317_, _24182_);
  nand (_24184_, _10276_, _07823_);
  nor (_24185_, _07823_, _24182_);
  nor (_24186_, _24185_, _07130_);
  nand (_24187_, _24186_, _24184_);
  and (_24188_, _07823_, \oc8051_golden_model_1.ACC [0]);
  or (_24189_, _24188_, _24185_);
  and (_24190_, _24189_, _06220_);
  or (_24192_, _24190_, _09842_);
  nor (_24193_, _08211_, _11817_);
  or (_24194_, _24193_, _24185_);
  and (_24195_, _24194_, _06160_);
  nor (_24196_, _07056_, _24182_);
  and (_24197_, _24189_, _07056_);
  or (_24198_, _24197_, _24196_);
  and (_24199_, _24198_, _06161_);
  or (_24200_, _24199_, _06217_);
  or (_24201_, _24200_, _24195_);
  and (_24203_, _24201_, _06229_);
  or (_24204_, _24203_, _24192_);
  and (_24205_, _07823_, _07049_);
  and (_24206_, _06132_, _07075_);
  or (_24207_, _24185_, _24206_);
  or (_24208_, _24207_, _24205_);
  and (_24209_, _24208_, _24204_);
  or (_24210_, _24209_, _06116_);
  and (_24211_, _09160_, _07823_);
  or (_24212_, _24185_, _06117_);
  or (_24214_, _24212_, _24211_);
  and (_24215_, _24214_, _24210_);
  or (_24216_, _24215_, _05787_);
  and (_24217_, _14260_, _07823_);
  or (_24218_, _24217_, _24185_);
  or (_24219_, _24218_, _06114_);
  and (_24220_, _24219_, _06111_);
  and (_24221_, _24220_, _24216_);
  and (_24222_, _07823_, _08708_);
  or (_24223_, _24222_, _24185_);
  and (_24225_, _24223_, _06110_);
  or (_24226_, _24225_, _06297_);
  or (_24227_, _24226_, _24221_);
  and (_24228_, _14275_, _07823_);
  or (_24229_, _24228_, _24185_);
  or (_24230_, _24229_, _07127_);
  and (_24231_, _24230_, _07125_);
  and (_24232_, _24231_, _24227_);
  nor (_24233_, _12321_, _11817_);
  or (_24234_, _24233_, _24185_);
  and (_24236_, _24184_, _06402_);
  and (_24237_, _24236_, _24234_);
  or (_24238_, _24237_, _24232_);
  and (_24239_, _24238_, _07132_);
  nand (_24240_, _24223_, _06306_);
  nor (_24241_, _24240_, _24193_);
  or (_24242_, _24241_, _06411_);
  or (_24243_, _24242_, _24239_);
  and (_24244_, _24243_, _24187_);
  or (_24245_, _24244_, _06303_);
  and (_24247_, _14167_, _07823_);
  or (_24248_, _24185_, _08819_);
  or (_24249_, _24248_, _24247_);
  and (_24250_, _24249_, _08824_);
  and (_24251_, _24250_, _24245_);
  and (_24252_, _24234_, _06396_);
  or (_24253_, _24252_, _19287_);
  or (_24254_, _24253_, _24251_);
  or (_24255_, _24194_, _06630_);
  and (_24256_, _24255_, _01317_);
  and (_24258_, _24256_, _24254_);
  or (_24259_, _24258_, _24183_);
  and (_43678_, _24259_, _43100_);
  not (_24260_, \oc8051_golden_model_1.TH0 [1]);
  nor (_24261_, _01317_, _24260_);
  or (_24262_, _14442_, _11817_);
  or (_24263_, _07823_, \oc8051_golden_model_1.TH0 [1]);
  and (_24264_, _24263_, _05787_);
  and (_24265_, _24264_, _24262_);
  and (_24266_, _09115_, _07823_);
  nor (_24268_, _07823_, _24260_);
  or (_24269_, _24268_, _06117_);
  or (_24270_, _24269_, _24266_);
  and (_24271_, _14363_, _07823_);
  not (_24272_, _24271_);
  and (_24273_, _24272_, _24263_);
  or (_24274_, _24273_, _06161_);
  and (_24275_, _07823_, \oc8051_golden_model_1.ACC [1]);
  or (_24276_, _24275_, _24268_);
  and (_24277_, _24276_, _07056_);
  nor (_24279_, _07056_, _24260_);
  or (_24280_, _24279_, _06160_);
  or (_24281_, _24280_, _24277_);
  and (_24282_, _24281_, _07075_);
  and (_24283_, _24282_, _24274_);
  and (_24284_, _07823_, _07306_);
  or (_24285_, _24284_, _24268_);
  and (_24286_, _24285_, _06217_);
  or (_24287_, _24286_, _24283_);
  and (_24288_, _24287_, _06229_);
  and (_24290_, _24276_, _06220_);
  or (_24291_, _24290_, _09842_);
  or (_24292_, _24291_, _24288_);
  or (_24293_, _24285_, _06132_);
  and (_24294_, _24293_, _24292_);
  or (_24295_, _24294_, _06116_);
  and (_24296_, _24295_, _06114_);
  and (_24297_, _24296_, _24270_);
  or (_24298_, _24297_, _24265_);
  and (_24299_, _24298_, _06298_);
  or (_24301_, _14346_, _11817_);
  and (_24302_, _24301_, _06297_);
  nand (_24303_, _07823_, _06945_);
  and (_24304_, _24303_, _06110_);
  or (_24305_, _24304_, _24302_);
  and (_24306_, _24305_, _24263_);
  or (_24307_, _24306_, _06402_);
  or (_24308_, _24307_, _24299_);
  nor (_24309_, _10277_, _11817_);
  or (_24310_, _24309_, _24268_);
  nand (_24312_, _10275_, _07823_);
  and (_24313_, _24312_, _24310_);
  or (_24314_, _24313_, _07125_);
  and (_24315_, _24314_, _07132_);
  and (_24316_, _24315_, _24308_);
  or (_24317_, _14344_, _11817_);
  and (_24318_, _24263_, _06306_);
  and (_24319_, _24318_, _24317_);
  or (_24320_, _24319_, _06411_);
  or (_24321_, _24320_, _24316_);
  nor (_24323_, _24268_, _07130_);
  nand (_24324_, _24323_, _24312_);
  and (_24325_, _24324_, _08819_);
  and (_24326_, _24325_, _24321_);
  or (_24327_, _24303_, _08176_);
  and (_24328_, _24263_, _06303_);
  and (_24329_, _24328_, _24327_);
  or (_24330_, _24329_, _06396_);
  or (_24331_, _24330_, _24326_);
  or (_24332_, _24310_, _08824_);
  and (_24334_, _24332_, _06829_);
  and (_24335_, _24334_, _24331_);
  and (_24336_, _24273_, _06433_);
  or (_24337_, _24336_, _06440_);
  or (_24338_, _24337_, _24335_);
  or (_24339_, _24268_, _06444_);
  or (_24340_, _24339_, _24271_);
  and (_24341_, _24340_, _01317_);
  and (_24342_, _24341_, _24338_);
  or (_24343_, _24342_, _24261_);
  and (_43679_, _24343_, _43100_);
  and (_24345_, _01321_, \oc8051_golden_model_1.TH0 [2]);
  and (_24346_, _11817_, \oc8051_golden_model_1.TH0 [2]);
  and (_24347_, _09211_, _07823_);
  or (_24348_, _24347_, _24346_);
  and (_24349_, _24348_, _06116_);
  and (_24350_, _14542_, _07823_);
  or (_24351_, _24350_, _24346_);
  or (_24352_, _24351_, _06161_);
  and (_24353_, _07823_, \oc8051_golden_model_1.ACC [2]);
  or (_24355_, _24353_, _24346_);
  and (_24356_, _24355_, _07056_);
  and (_24357_, _07057_, \oc8051_golden_model_1.TH0 [2]);
  or (_24358_, _24357_, _06160_);
  or (_24359_, _24358_, _24356_);
  and (_24360_, _24359_, _07075_);
  and (_24361_, _24360_, _24352_);
  and (_24362_, _07823_, _07708_);
  or (_24363_, _24362_, _24346_);
  and (_24364_, _24363_, _06217_);
  or (_24366_, _24364_, _24361_);
  and (_24367_, _24366_, _06229_);
  and (_24368_, _24355_, _06220_);
  or (_24369_, _24368_, _09842_);
  or (_24370_, _24369_, _24367_);
  or (_24371_, _24363_, _06132_);
  and (_24372_, _24371_, _06117_);
  and (_24373_, _24372_, _24370_);
  or (_24374_, _24373_, _05787_);
  or (_24375_, _24374_, _24349_);
  and (_24378_, _14630_, _07823_);
  or (_24379_, _24346_, _06114_);
  or (_24380_, _24379_, _24378_);
  and (_24381_, _24380_, _06111_);
  and (_24382_, _24381_, _24375_);
  and (_24383_, _07823_, _08768_);
  or (_24384_, _24383_, _24346_);
  and (_24385_, _24384_, _06110_);
  or (_24386_, _24385_, _06297_);
  or (_24387_, _24386_, _24382_);
  and (_24389_, _14646_, _07823_);
  or (_24390_, _24346_, _07127_);
  or (_24391_, _24390_, _24389_);
  and (_24392_, _24391_, _07125_);
  and (_24393_, _24392_, _24387_);
  and (_24394_, _10282_, _07823_);
  or (_24395_, _24394_, _24346_);
  and (_24396_, _24395_, _06402_);
  or (_24397_, _24396_, _24393_);
  and (_24398_, _24397_, _07132_);
  or (_24400_, _24346_, _08248_);
  and (_24401_, _24384_, _06306_);
  and (_24402_, _24401_, _24400_);
  or (_24403_, _24402_, _24398_);
  and (_24404_, _24403_, _07130_);
  and (_24405_, _24355_, _06411_);
  and (_24406_, _24405_, _24400_);
  or (_24407_, _24406_, _06303_);
  or (_24408_, _24407_, _24404_);
  and (_24409_, _14643_, _07823_);
  or (_24411_, _24346_, _08819_);
  or (_24412_, _24411_, _24409_);
  and (_24413_, _24412_, _08824_);
  and (_24414_, _24413_, _24408_);
  nor (_24415_, _10281_, _11817_);
  or (_24416_, _24415_, _24346_);
  and (_24417_, _24416_, _06396_);
  or (_24418_, _24417_, _24414_);
  and (_24419_, _24418_, _06829_);
  and (_24420_, _24351_, _06433_);
  or (_24422_, _24420_, _06440_);
  or (_24423_, _24422_, _24419_);
  and (_24424_, _14710_, _07823_);
  or (_24425_, _24346_, _06444_);
  or (_24426_, _24425_, _24424_);
  and (_24427_, _24426_, _01317_);
  and (_24428_, _24427_, _24423_);
  or (_24429_, _24428_, _24345_);
  and (_43680_, _24429_, _43100_);
  and (_24430_, _11817_, \oc8051_golden_model_1.TH0 [3]);
  and (_24432_, _14738_, _07823_);
  or (_24433_, _24432_, _24430_);
  or (_24434_, _24433_, _06161_);
  and (_24435_, _07823_, \oc8051_golden_model_1.ACC [3]);
  or (_24436_, _24435_, _24430_);
  and (_24437_, _24436_, _07056_);
  and (_24438_, _07057_, \oc8051_golden_model_1.TH0 [3]);
  or (_24439_, _24438_, _06160_);
  or (_24440_, _24439_, _24437_);
  and (_24441_, _24440_, _07075_);
  and (_24443_, _24441_, _24434_);
  and (_24444_, _07823_, _07544_);
  or (_24445_, _24444_, _24430_);
  and (_24446_, _24445_, _06217_);
  or (_24447_, _24446_, _24443_);
  and (_24448_, _24447_, _06229_);
  and (_24449_, _24436_, _06220_);
  or (_24450_, _24449_, _09842_);
  or (_24451_, _24450_, _24448_);
  or (_24452_, _24445_, _06132_);
  and (_24454_, _24452_, _24451_);
  or (_24455_, _24454_, _06116_);
  and (_24456_, _09210_, _07823_);
  or (_24457_, _24430_, _06117_);
  or (_24458_, _24457_, _24456_);
  and (_24459_, _24458_, _06114_);
  and (_24460_, _24459_, _24455_);
  and (_24461_, _14825_, _07823_);
  or (_24462_, _24461_, _24430_);
  and (_24463_, _24462_, _05787_);
  or (_24465_, _24463_, _11136_);
  or (_24466_, _24465_, _24460_);
  and (_24467_, _14727_, _07823_);
  or (_24468_, _24430_, _07127_);
  or (_24469_, _24468_, _24467_);
  and (_24470_, _07823_, _08712_);
  or (_24471_, _24470_, _24430_);
  or (_24472_, _24471_, _06111_);
  and (_24473_, _24472_, _07125_);
  and (_24474_, _24473_, _24469_);
  and (_24476_, _24474_, _24466_);
  and (_24477_, _12318_, _07823_);
  or (_24478_, _24477_, _24430_);
  and (_24479_, _24478_, _06402_);
  or (_24480_, _24479_, _24476_);
  and (_24481_, _24480_, _07132_);
  or (_24482_, _24430_, _08140_);
  and (_24483_, _24471_, _06306_);
  and (_24484_, _24483_, _24482_);
  or (_24485_, _24484_, _24481_);
  and (_24487_, _24485_, _07130_);
  and (_24488_, _24436_, _06411_);
  and (_24489_, _24488_, _24482_);
  or (_24490_, _24489_, _06303_);
  or (_24491_, _24490_, _24487_);
  and (_24492_, _14724_, _07823_);
  or (_24493_, _24430_, _08819_);
  or (_24494_, _24493_, _24492_);
  and (_24495_, _24494_, _08824_);
  and (_24496_, _24495_, _24491_);
  nor (_24498_, _10273_, _11817_);
  or (_24499_, _24498_, _24430_);
  and (_24500_, _24499_, _06396_);
  or (_24501_, _24500_, _06433_);
  or (_24502_, _24501_, _24496_);
  or (_24503_, _24433_, _06829_);
  and (_24504_, _24503_, _06444_);
  and (_24505_, _24504_, _24502_);
  and (_24506_, _14897_, _07823_);
  or (_24507_, _24506_, _24430_);
  and (_24509_, _24507_, _06440_);
  or (_24510_, _24509_, _01321_);
  or (_24511_, _24510_, _24505_);
  or (_24512_, _01317_, \oc8051_golden_model_1.TH0 [3]);
  and (_24513_, _24512_, _43100_);
  and (_43682_, _24513_, _24511_);
  and (_24514_, _11817_, \oc8051_golden_model_1.TH0 [4]);
  and (_24515_, _08336_, _07823_);
  or (_24516_, _24515_, _24514_);
  or (_24517_, _24516_, _06132_);
  and (_24519_, _14928_, _07823_);
  or (_24520_, _24519_, _24514_);
  or (_24521_, _24520_, _06161_);
  and (_24522_, _07823_, \oc8051_golden_model_1.ACC [4]);
  or (_24523_, _24522_, _24514_);
  and (_24524_, _24523_, _07056_);
  and (_24525_, _07057_, \oc8051_golden_model_1.TH0 [4]);
  or (_24526_, _24525_, _06160_);
  or (_24527_, _24526_, _24524_);
  and (_24528_, _24527_, _07075_);
  and (_24530_, _24528_, _24521_);
  and (_24531_, _24516_, _06217_);
  or (_24532_, _24531_, _24530_);
  and (_24533_, _24532_, _06229_);
  and (_24534_, _24523_, _06220_);
  or (_24535_, _24534_, _09842_);
  or (_24536_, _24535_, _24533_);
  and (_24537_, _24536_, _24517_);
  or (_24538_, _24537_, _06116_);
  and (_24539_, _09209_, _07823_);
  or (_24541_, _24514_, _06117_);
  or (_24542_, _24541_, _24539_);
  and (_24543_, _24542_, _06114_);
  and (_24544_, _24543_, _24538_);
  and (_24545_, _15013_, _07823_);
  or (_24546_, _24545_, _24514_);
  and (_24547_, _24546_, _05787_);
  or (_24548_, _24547_, _24544_);
  or (_24549_, _24548_, _11136_);
  and (_24550_, _15029_, _07823_);
  or (_24552_, _24514_, _07127_);
  or (_24553_, _24552_, _24550_);
  and (_24554_, _08715_, _07823_);
  or (_24555_, _24554_, _24514_);
  or (_24556_, _24555_, _06111_);
  and (_24557_, _24556_, _07125_);
  and (_24558_, _24557_, _24553_);
  and (_24559_, _24558_, _24549_);
  and (_24560_, _10289_, _07823_);
  or (_24561_, _24560_, _24514_);
  and (_24563_, _24561_, _06402_);
  or (_24564_, _24563_, _24559_);
  and (_24565_, _24564_, _07132_);
  or (_24566_, _24514_, _08339_);
  and (_24567_, _24555_, _06306_);
  and (_24568_, _24567_, _24566_);
  or (_24569_, _24568_, _24565_);
  and (_24570_, _24569_, _07130_);
  and (_24571_, _24523_, _06411_);
  and (_24572_, _24571_, _24566_);
  or (_24574_, _24572_, _06303_);
  or (_24575_, _24574_, _24570_);
  and (_24576_, _15026_, _07823_);
  or (_24577_, _24514_, _08819_);
  or (_24578_, _24577_, _24576_);
  and (_24579_, _24578_, _08824_);
  and (_24580_, _24579_, _24575_);
  nor (_24581_, _10288_, _11817_);
  or (_24582_, _24581_, _24514_);
  and (_24583_, _24582_, _06396_);
  or (_24585_, _24583_, _06433_);
  or (_24586_, _24585_, _24580_);
  or (_24587_, _24520_, _06829_);
  and (_24588_, _24587_, _06444_);
  and (_24589_, _24588_, _24586_);
  and (_24590_, _15087_, _07823_);
  or (_24591_, _24590_, _24514_);
  and (_24592_, _24591_, _06440_);
  or (_24593_, _24592_, _01321_);
  or (_24594_, _24593_, _24589_);
  or (_24596_, _01317_, \oc8051_golden_model_1.TH0 [4]);
  and (_24597_, _24596_, _43100_);
  and (_43683_, _24597_, _24594_);
  and (_24598_, _11817_, \oc8051_golden_model_1.TH0 [5]);
  and (_24599_, _15119_, _07823_);
  or (_24600_, _24599_, _24598_);
  or (_24601_, _24600_, _06161_);
  and (_24602_, _07823_, \oc8051_golden_model_1.ACC [5]);
  or (_24603_, _24602_, _24598_);
  and (_24604_, _24603_, _07056_);
  and (_24605_, _07057_, \oc8051_golden_model_1.TH0 [5]);
  or (_24606_, _24605_, _06160_);
  or (_24607_, _24606_, _24604_);
  and (_24608_, _24607_, _07075_);
  and (_24609_, _24608_, _24601_);
  and (_24610_, _08101_, _07823_);
  or (_24611_, _24610_, _24598_);
  and (_24612_, _24611_, _06217_);
  or (_24613_, _24612_, _24609_);
  and (_24614_, _24613_, _06229_);
  and (_24617_, _24603_, _06220_);
  or (_24618_, _24617_, _09842_);
  or (_24619_, _24618_, _24614_);
  or (_24620_, _24611_, _06132_);
  and (_24621_, _24620_, _24619_);
  or (_24622_, _24621_, _06116_);
  and (_24623_, _09208_, _07823_);
  or (_24624_, _24598_, _06117_);
  or (_24625_, _24624_, _24623_);
  and (_24626_, _24625_, _06114_);
  and (_24628_, _24626_, _24622_);
  and (_24629_, _15203_, _07823_);
  or (_24630_, _24629_, _24598_);
  and (_24631_, _24630_, _05787_);
  or (_24632_, _24631_, _11136_);
  or (_24633_, _24632_, _24628_);
  and (_24634_, _15219_, _07823_);
  or (_24635_, _24598_, _07127_);
  or (_24636_, _24635_, _24634_);
  and (_24637_, _08736_, _07823_);
  or (_24639_, _24637_, _24598_);
  or (_24640_, _24639_, _06111_);
  and (_24641_, _24640_, _07125_);
  and (_24642_, _24641_, _24636_);
  and (_24643_, _24642_, _24633_);
  and (_24644_, _12325_, _07823_);
  or (_24645_, _24644_, _24598_);
  and (_24646_, _24645_, _06402_);
  or (_24647_, _24646_, _24643_);
  and (_24648_, _24647_, _07132_);
  or (_24650_, _24598_, _08104_);
  and (_24651_, _24639_, _06306_);
  and (_24652_, _24651_, _24650_);
  or (_24653_, _24652_, _24648_);
  and (_24654_, _24653_, _07130_);
  and (_24655_, _24603_, _06411_);
  and (_24656_, _24655_, _24650_);
  or (_24657_, _24656_, _06303_);
  or (_24658_, _24657_, _24654_);
  and (_24659_, _15216_, _07823_);
  or (_24661_, _24598_, _08819_);
  or (_24662_, _24661_, _24659_);
  and (_24663_, _24662_, _08824_);
  and (_24664_, _24663_, _24658_);
  nor (_24665_, _10269_, _11817_);
  or (_24666_, _24665_, _24598_);
  and (_24667_, _24666_, _06396_);
  or (_24668_, _24667_, _06433_);
  or (_24669_, _24668_, _24664_);
  or (_24670_, _24600_, _06829_);
  and (_24672_, _24670_, _06444_);
  and (_24673_, _24672_, _24669_);
  and (_24674_, _15275_, _07823_);
  or (_24675_, _24674_, _24598_);
  and (_24676_, _24675_, _06440_);
  or (_24677_, _24676_, _01321_);
  or (_24678_, _24677_, _24673_);
  or (_24679_, _01317_, \oc8051_golden_model_1.TH0 [5]);
  and (_24680_, _24679_, _43100_);
  and (_43684_, _24680_, _24678_);
  and (_24682_, _11817_, \oc8051_golden_model_1.TH0 [6]);
  or (_24683_, _24682_, _08015_);
  and (_24684_, _15402_, _07823_);
  or (_24685_, _24684_, _24682_);
  and (_24686_, _24685_, _06306_);
  and (_24687_, _24686_, _24683_);
  and (_24688_, _15300_, _07823_);
  or (_24689_, _24688_, _24682_);
  or (_24690_, _24689_, _06161_);
  and (_24691_, _07823_, \oc8051_golden_model_1.ACC [6]);
  or (_24693_, _24691_, _24682_);
  and (_24694_, _24693_, _07056_);
  and (_24695_, _07057_, \oc8051_golden_model_1.TH0 [6]);
  or (_24696_, _24695_, _06160_);
  or (_24697_, _24696_, _24694_);
  and (_24698_, _24697_, _07075_);
  and (_24699_, _24698_, _24690_);
  and (_24700_, _08012_, _07823_);
  or (_24701_, _24700_, _24682_);
  and (_24702_, _24701_, _06217_);
  or (_24704_, _24702_, _24699_);
  and (_24705_, _24704_, _06229_);
  and (_24706_, _24693_, _06220_);
  or (_24707_, _24706_, _09842_);
  or (_24708_, _24707_, _24705_);
  or (_24709_, _24701_, _06132_);
  and (_24710_, _24709_, _24708_);
  or (_24711_, _24710_, _06116_);
  and (_24712_, _09207_, _07823_);
  or (_24713_, _24682_, _06117_);
  or (_24715_, _24713_, _24712_);
  and (_24716_, _24715_, _06114_);
  and (_24717_, _24716_, _24711_);
  and (_24718_, _15395_, _07823_);
  or (_24719_, _24718_, _24682_);
  and (_24720_, _24719_, _05787_);
  or (_24721_, _24720_, _11136_);
  or (_24722_, _24721_, _24717_);
  and (_24723_, _15413_, _07823_);
  or (_24724_, _24682_, _07127_);
  or (_24726_, _24724_, _24723_);
  or (_24727_, _24685_, _06111_);
  and (_24728_, _24727_, _07125_);
  and (_24729_, _24728_, _24726_);
  and (_24730_, _24729_, _24722_);
  and (_24731_, _10295_, _07823_);
  or (_24732_, _24731_, _24682_);
  and (_24733_, _24732_, _06402_);
  or (_24734_, _24733_, _24730_);
  and (_24735_, _24734_, _07132_);
  or (_24737_, _24735_, _24687_);
  and (_24738_, _24737_, _07130_);
  and (_24739_, _24693_, _06411_);
  and (_24740_, _24739_, _24683_);
  or (_24741_, _24740_, _06303_);
  or (_24742_, _24741_, _24738_);
  and (_24743_, _15410_, _07823_);
  or (_24744_, _24682_, _08819_);
  or (_24745_, _24744_, _24743_);
  and (_24746_, _24745_, _08824_);
  and (_24748_, _24746_, _24742_);
  nor (_24749_, _10294_, _11817_);
  or (_24750_, _24749_, _24682_);
  and (_24751_, _24750_, _06396_);
  or (_24752_, _24751_, _06433_);
  or (_24753_, _24752_, _24748_);
  or (_24754_, _24689_, _06829_);
  and (_24755_, _24754_, _06444_);
  and (_24756_, _24755_, _24753_);
  and (_24757_, _15478_, _07823_);
  or (_24759_, _24757_, _24682_);
  and (_24760_, _24759_, _06440_);
  or (_24761_, _24760_, _01321_);
  or (_24762_, _24761_, _24756_);
  or (_24763_, _01317_, \oc8051_golden_model_1.TH0 [6]);
  and (_24764_, _24763_, _43100_);
  and (_43685_, _24764_, _24762_);
  and (_24765_, _12744_, _12735_);
  nor (_24766_, _24765_, _05444_);
  and (_24767_, _12682_, \oc8051_golden_model_1.PC [0]);
  and (_24769_, _06758_, \oc8051_golden_model_1.PC [0]);
  nor (_24770_, _24769_, _12032_);
  nor (_24771_, _24770_, _12682_);
  nor (_24772_, _24771_, _24767_);
  and (_24773_, _24772_, _05748_);
  and (_24774_, _12711_, _12719_);
  nor (_24775_, _24774_, _05444_);
  and (_24776_, _11905_, _12693_);
  nor (_24777_, _24776_, _05444_);
  nor (_24778_, _10694_, _05444_);
  and (_24780_, _10694_, _05444_);
  nor (_24781_, _24780_, _24778_);
  nor (_24782_, _24781_, _12539_);
  and (_24783_, _11912_, _08819_);
  nor (_24784_, _24783_, _05444_);
  and (_24785_, _11914_, _07132_);
  nor (_24786_, _24785_, _05444_);
  and (_24787_, _11919_, _07127_);
  nor (_24788_, _24787_, _05444_);
  and (_24789_, _06110_, _05444_);
  not (_24791_, _05791_);
  nor (_24792_, _06758_, _24791_);
  nor (_24793_, _06758_, _05769_);
  and (_24794_, _06758_, _06581_);
  nor (_24795_, _12263_, _05444_);
  nor (_24796_, _12266_, _05444_);
  and (_24797_, _12266_, _05444_);
  nor (_24798_, _24797_, _24796_);
  and (_24799_, _12263_, _06582_);
  not (_24800_, _24799_);
  nor (_24802_, _24800_, _24798_);
  nor (_24803_, _24802_, _24795_);
  not (_24804_, _24803_);
  nor (_24805_, _24804_, _24794_);
  nor (_24806_, _24805_, _08445_);
  and (_24807_, _12258_, \oc8051_golden_model_1.PC [0]);
  and (_24808_, _06107_, _05444_);
  nor (_24809_, _24808_, _12200_);
  and (_24810_, _24809_, _12256_);
  or (_24811_, _24810_, _24807_);
  nor (_24813_, _24811_, _08443_);
  nor (_24814_, _24813_, _24806_);
  nor (_24815_, _24814_, _07064_);
  and (_24816_, _07064_, \oc8051_golden_model_1.PC [0]);
  nor (_24817_, _24816_, _06160_);
  not (_24818_, _24817_);
  nor (_24819_, _24818_, _24815_);
  not (_24820_, _24819_);
  not (_24821_, _12134_);
  not (_24822_, _24770_);
  and (_24824_, _24822_, _12139_);
  and (_24825_, _12141_, \oc8051_golden_model_1.PC [0]);
  or (_24826_, _24825_, _06161_);
  nor (_24827_, _24826_, _24824_);
  nor (_24828_, _24827_, _24821_);
  and (_24829_, _24828_, _24820_);
  nor (_24830_, _12134_, _05444_);
  nor (_24831_, _24830_, _07485_);
  not (_24832_, _24831_);
  nor (_24833_, _24832_, _24829_);
  nor (_24835_, _06758_, _05764_);
  and (_24836_, _12300_, _12292_);
  not (_24837_, _24836_);
  nor (_24838_, _24837_, _24835_);
  not (_24839_, _24838_);
  nor (_24840_, _24839_, _24833_);
  nor (_24841_, _24836_, _05444_);
  nor (_24842_, _24841_, _12304_);
  not (_24843_, _24842_);
  nor (_24844_, _24843_, _24840_);
  nor (_24846_, _24844_, _24793_);
  or (_24847_, _24846_, _12126_);
  and (_24848_, _12120_, \oc8051_golden_model_1.PC [0]);
  nor (_24849_, _24770_, _12120_);
  or (_24850_, _24849_, _12125_);
  or (_24851_, _24850_, _24848_);
  and (_24852_, _24851_, _12089_);
  and (_24853_, _24852_, _24847_);
  nor (_24854_, _24853_, _06236_);
  nor (_24855_, _11956_, \oc8051_golden_model_1.PC [0]);
  and (_24857_, _24770_, _11956_);
  or (_24858_, _24857_, _12089_);
  or (_24859_, _24858_, _24855_);
  and (_24860_, _24859_, _24854_);
  and (_24861_, _12329_, _05444_);
  nor (_24862_, _24822_, _12329_);
  nor (_24863_, _24862_, _24861_);
  nor (_24864_, _24863_, _06643_);
  nor (_24865_, _24864_, _24860_);
  nor (_24866_, _24865_, _06295_);
  and (_24868_, _12346_, _05444_);
  nor (_24869_, _24822_, _12346_);
  or (_24870_, _24869_, _24868_);
  and (_24871_, _24870_, _06295_);
  or (_24872_, _24871_, _24866_);
  and (_24873_, _24872_, _11925_);
  and (_24874_, _11924_, _05444_);
  or (_24875_, _24874_, _24873_);
  and (_24876_, _24875_, _05760_);
  nor (_24877_, _06758_, _05760_);
  nor (_24879_, _24877_, _12373_);
  not (_24880_, _24879_);
  nor (_24881_, _24880_, _24876_);
  not (_24882_, _05775_);
  nor (_24883_, _12369_, _05444_);
  nor (_24884_, _24883_, _24882_);
  not (_24885_, _24884_);
  nor (_24886_, _24885_, _24881_);
  nor (_24887_, _06758_, _05775_);
  and (_24888_, _12381_, _05805_);
  not (_24890_, _24888_);
  nor (_24891_, _24890_, _24887_);
  not (_24892_, _24891_);
  nor (_24893_, _24892_, _24886_);
  nor (_24894_, _24888_, _05444_);
  nor (_24895_, _24894_, _05791_);
  not (_24896_, _24895_);
  nor (_24897_, _24896_, _24893_);
  nor (_24898_, _06293_, _05787_);
  and (_24899_, _24898_, _11922_);
  not (_24901_, _24899_);
  or (_24902_, _24901_, _24897_);
  nor (_24903_, _24902_, _24792_);
  nor (_24904_, _24899_, _05444_);
  nor (_24905_, _24904_, _05829_);
  not (_24906_, _24905_);
  nor (_24907_, _24906_, _24903_);
  nor (_24908_, _06758_, _05830_);
  or (_24909_, _24908_, _12416_);
  nor (_24910_, _24909_, _24907_);
  nor (_24912_, _24809_, _12417_);
  nor (_24913_, _24912_, _24910_);
  and (_24914_, _24913_, _06111_);
  or (_24915_, _24914_, _24789_);
  and (_24916_, _24915_, _12432_);
  and (_24917_, _12431_, _05809_);
  or (_24918_, _24917_, _24916_);
  and (_24919_, _24918_, _05836_);
  nor (_24920_, _06758_, _05836_);
  or (_24921_, _24920_, _24919_);
  and (_24923_, _24921_, _12474_);
  not (_24924_, _24787_);
  nor (_24925_, _24809_, _11101_);
  and (_24926_, _11101_, _05444_);
  nor (_24927_, _24926_, _12474_);
  not (_24928_, _24927_);
  nor (_24929_, _24928_, _24925_);
  nor (_24930_, _24929_, _24924_);
  not (_24931_, _24930_);
  nor (_24932_, _24931_, _24923_);
  nor (_24934_, _24932_, _24788_);
  and (_24935_, _24934_, _05834_);
  nor (_24936_, _06758_, _05834_);
  or (_24937_, _24936_, _24935_);
  and (_24938_, _24937_, _12497_);
  not (_24939_, _24785_);
  nor (_24940_, _24809_, _12480_);
  nor (_24941_, _11101_, \oc8051_golden_model_1.PC [0]);
  nor (_24942_, _24941_, _12497_);
  not (_24943_, _24942_);
  nor (_24945_, _24943_, _24940_);
  nor (_24946_, _24945_, _24939_);
  not (_24947_, _24946_);
  nor (_24948_, _24947_, _24938_);
  nor (_24949_, _24948_, _24786_);
  and (_24950_, _24949_, _05848_);
  nor (_24951_, _06758_, _05848_);
  or (_24952_, _24951_, _24950_);
  and (_24953_, _24952_, _12518_);
  not (_24954_, _24783_);
  nor (_24956_, _24809_, \oc8051_golden_model_1.PSW [7]);
  and (_24957_, \oc8051_golden_model_1.PSW [7], _05444_);
  nor (_24958_, _24957_, _12518_);
  not (_24959_, _24958_);
  nor (_24960_, _24959_, _24956_);
  nor (_24961_, _24960_, _24954_);
  not (_24962_, _24961_);
  nor (_24963_, _24962_, _24953_);
  nor (_24964_, _24963_, _24784_);
  and (_24965_, _24964_, _05843_);
  nor (_24967_, _06758_, _05843_);
  or (_24968_, _24967_, _24965_);
  and (_24969_, _24968_, _12539_);
  and (_24970_, _11907_, _10926_);
  not (_24971_, _24970_);
  or (_24972_, _24971_, _24969_);
  nor (_24973_, _24972_, _24782_);
  nor (_24974_, _24970_, _05444_);
  nor (_24975_, _24974_, _06417_);
  not (_24976_, _24975_);
  nor (_24978_, _24976_, _24973_);
  and (_24979_, _09160_, _06417_);
  or (_24980_, _24979_, _24978_);
  and (_24981_, _24980_, _05846_);
  nor (_24982_, _06758_, _05846_);
  or (_24983_, _24982_, _24981_);
  and (_24984_, _24983_, _06421_);
  not (_24985_, _24776_);
  and (_24986_, _24822_, _12682_);
  nor (_24987_, _12682_, _05444_);
  or (_24989_, _24987_, _06421_);
  nor (_24990_, _24989_, _24986_);
  nor (_24991_, _24990_, _24985_);
  not (_24992_, _24991_);
  nor (_24993_, _24992_, _24984_);
  nor (_24994_, _24993_, _24777_);
  and (_24995_, _24994_, _06168_);
  and (_24996_, _09160_, _06167_);
  or (_24997_, _24996_, _24995_);
  and (_24998_, _24997_, _12703_);
  nor (_25000_, _06758_, _12703_);
  nor (_25001_, _25000_, _24998_);
  nor (_25002_, _25001_, _06165_);
  not (_25003_, _24774_);
  and (_25004_, _24772_, _06165_);
  nor (_25005_, _25004_, _25003_);
  not (_25006_, _25005_);
  nor (_25007_, _25006_, _25002_);
  or (_25008_, _25007_, _24775_);
  nand (_25009_, _25008_, _07160_);
  and (_25011_, _07577_, _06758_);
  nor (_25012_, _25011_, _05748_);
  nand (_25013_, _25012_, _25009_);
  nand (_25014_, _25013_, _24765_);
  nor (_25015_, _25014_, _24773_);
  or (_25016_, _25015_, _24766_);
  nor (_25017_, _06305_, _05821_);
  nand (_25018_, _25017_, _25016_);
  not (_25019_, _25017_);
  and (_25020_, _25019_, _06758_);
  nor (_25022_, _25020_, _12754_);
  and (_25023_, _25022_, _25018_);
  and (_25024_, _12754_, _05444_);
  or (_25025_, _25024_, _25023_);
  or (_25026_, _25025_, _01321_);
  or (_25027_, _01317_, \oc8051_golden_model_1.PC [0]);
  and (_25028_, _25027_, _43100_);
  and (_43687_, _25028_, _25026_);
  and (_25029_, _06440_, _05407_);
  and (_25030_, _12682_, _05879_);
  nor (_25032_, _12034_, _12032_);
  nor (_25033_, _25032_, _12035_);
  nor (_25034_, _25033_, _12682_);
  nor (_25035_, _25034_, _25030_);
  and (_25036_, _25035_, _05748_);
  and (_25037_, _06433_, _05407_);
  nor (_25038_, _08362_, _05879_);
  or (_25039_, _11905_, _05879_);
  or (_25040_, _11907_, _05879_);
  or (_25041_, _11914_, _05879_);
  or (_25043_, _11919_, _05879_);
  or (_25044_, _08787_, _05407_);
  or (_25045_, _12381_, _05879_);
  nor (_25046_, _12202_, _12200_);
  nor (_25047_, _25046_, _12203_);
  and (_25048_, _25047_, _12256_);
  and (_25049_, _12258_, _05407_);
  or (_25050_, _25049_, _25048_);
  or (_25051_, _25050_, _08443_);
  or (_25052_, _12263_, _05879_);
  nor (_25054_, _06945_, _06582_);
  not (_25055_, _12263_);
  and (_25056_, _06653_, _05444_);
  nor (_25057_, _12265_, _05444_);
  nor (_25058_, _25057_, _06545_);
  nor (_25059_, _25058_, _25056_);
  or (_25060_, _25059_, \oc8051_golden_model_1.PC [1]);
  nand (_25061_, _25059_, \oc8051_golden_model_1.PC [1]);
  and (_25062_, _25061_, _06582_);
  and (_25063_, _25062_, _25060_);
  or (_25065_, _25063_, _25055_);
  or (_25066_, _25065_, _25054_);
  and (_25067_, _25066_, _25052_);
  or (_25068_, _25067_, _08445_);
  and (_25069_, _25068_, _07065_);
  and (_25070_, _25069_, _25051_);
  and (_25071_, _07064_, _05879_);
  or (_25072_, _25071_, _06160_);
  or (_25073_, _25072_, _25070_);
  and (_25074_, _25033_, _12139_);
  and (_25076_, _12141_, _05878_);
  or (_25077_, _25076_, _06161_);
  or (_25078_, _25077_, _25074_);
  and (_25079_, _25078_, _25073_);
  or (_25080_, _25079_, _24821_);
  or (_25081_, _12134_, _05879_);
  and (_25082_, _25081_, _06157_);
  and (_25083_, _25082_, _25080_);
  and (_25084_, _06156_, _05407_);
  or (_25085_, _25084_, _07485_);
  or (_25087_, _25085_, _25083_);
  nand (_25088_, _06945_, _07485_);
  and (_25089_, _25088_, _07075_);
  and (_25090_, _25089_, _25087_);
  nand (_25091_, _06217_, _05407_);
  nand (_25092_, _25091_, _12292_);
  or (_25093_, _25092_, _25090_);
  or (_25094_, _12292_, _05879_);
  and (_25095_, _25094_, _06229_);
  and (_25096_, _25095_, _25093_);
  nand (_25098_, _06220_, _05407_);
  nand (_25099_, _25098_, _12300_);
  or (_25100_, _25099_, _25096_);
  or (_25101_, _12300_, _05879_);
  and (_25102_, _25101_, _06153_);
  and (_25103_, _25102_, _25100_);
  and (_25104_, _06152_, _05407_);
  or (_25105_, _25104_, _12304_);
  or (_25106_, _25105_, _25103_);
  nand (_25107_, _06945_, _12304_);
  and (_25109_, _25107_, _07191_);
  and (_25110_, _25109_, _25106_);
  nand (_25111_, _06151_, _05407_);
  nand (_25112_, _25111_, _12125_);
  or (_25113_, _25112_, _25110_);
  nor (_25114_, _06687_, _06236_);
  or (_25115_, _25033_, _12120_);
  nand (_25116_, _12120_, _05879_);
  and (_25117_, _25116_, _25115_);
  or (_25118_, _25117_, _12125_);
  and (_25120_, _25118_, _25114_);
  and (_25121_, _25120_, _25113_);
  and (_25122_, _12329_, _05878_);
  not (_25123_, _12329_);
  and (_25124_, _25033_, _25123_);
  or (_25125_, _25124_, _25122_);
  and (_25126_, _25125_, _06236_);
  and (_25127_, _11958_, _05878_);
  and (_25128_, _25033_, _11956_);
  or (_25129_, _25128_, _25127_);
  and (_25131_, _25129_, _06687_);
  or (_25132_, _25131_, _25126_);
  or (_25133_, _25132_, _25121_);
  and (_25134_, _25133_, _12317_);
  or (_25135_, _25033_, _12346_);
  nand (_25136_, _12346_, _05879_);
  and (_25137_, _25136_, _06295_);
  and (_25138_, _25137_, _25135_);
  or (_25139_, _25138_, _11924_);
  or (_25140_, _25139_, _25134_);
  nand (_25142_, _11924_, _05878_);
  and (_25143_, _25142_, _25140_);
  or (_25144_, _25143_, _06145_);
  nand (_25145_, _06145_, \oc8051_golden_model_1.PC [1]);
  and (_25146_, _25145_, _05760_);
  and (_25147_, _25146_, _25144_);
  nor (_25148_, _06945_, _05760_);
  nor (_25149_, _07292_, _06701_);
  and (_25150_, _25149_, _12359_);
  and (_25151_, _25150_, _12356_);
  not (_25152_, _25151_);
  or (_25153_, _25152_, _25148_);
  or (_25154_, _25153_, _25147_);
  or (_25155_, _25151_, _05407_);
  and (_25156_, _25155_, _12367_);
  and (_25157_, _25156_, _25154_);
  nand (_25158_, _12366_, _05879_);
  nand (_25159_, _25158_, _12368_);
  or (_25160_, _25159_, _25157_);
  or (_25161_, _12368_, _05879_);
  and (_25164_, _25161_, _13844_);
  and (_25165_, _25164_, _25160_);
  and (_25166_, _06255_, _05407_);
  or (_25167_, _25166_, _24882_);
  or (_25168_, _25167_, _25165_);
  nand (_25169_, _06945_, _24882_);
  and (_25170_, _25169_, _13843_);
  and (_25171_, _25170_, _25168_);
  or (_25172_, _12379_, _10545_);
  and (_25173_, _06254_, _05407_);
  nor (_25175_, _25173_, _25172_);
  nand (_25176_, _25175_, _10553_);
  or (_25177_, _25176_, _25171_);
  and (_25178_, _25177_, _25045_);
  or (_25179_, _25178_, _12386_);
  or (_25180_, _12385_, _05407_);
  and (_25181_, _25180_, _05805_);
  and (_25182_, _25181_, _25179_);
  nor (_25183_, _05878_, _05805_);
  or (_25184_, _25183_, _06139_);
  or (_25186_, _25184_, _25182_);
  nand (_25187_, _06139_, \oc8051_golden_model_1.PC [1]);
  and (_25188_, _25187_, _25186_);
  or (_25189_, _25188_, _05791_);
  nand (_25190_, _06945_, _05791_);
  and (_25191_, _25190_, _11296_);
  and (_25192_, _25191_, _25189_);
  nand (_25193_, _06293_, _05878_);
  nand (_25194_, _25193_, _06133_);
  or (_25195_, _25194_, _25192_);
  or (_25197_, _06133_, _05407_);
  and (_25198_, _25197_, _06114_);
  and (_25199_, _25198_, _25195_);
  nand (_25200_, _05878_, _05787_);
  nand (_25201_, _25200_, _11922_);
  or (_25202_, _25201_, _25199_);
  or (_25203_, _11922_, _05879_);
  and (_25204_, _25203_, _06762_);
  and (_25205_, _25204_, _25202_);
  and (_25206_, _06209_, _05407_);
  or (_25208_, _25206_, _05829_);
  or (_25209_, _25208_, _25205_);
  nand (_25210_, _06945_, _05829_);
  and (_25211_, _25210_, _12417_);
  and (_25212_, _25211_, _25209_);
  and (_25213_, _25047_, _12416_);
  or (_25214_, _25213_, _08788_);
  or (_25215_, _25214_, _25212_);
  and (_25216_, _25215_, _25044_);
  or (_25217_, _25216_, _06110_);
  nand (_25219_, _06110_, _05879_);
  and (_25220_, _25219_, _10752_);
  and (_25221_, _25220_, _25217_);
  and (_25222_, _10751_, _05407_);
  or (_25223_, _25222_, _12431_);
  or (_25224_, _25223_, _25221_);
  or (_25225_, _12432_, _05876_);
  and (_25226_, _25225_, _06768_);
  and (_25227_, _25226_, _25224_);
  and (_25228_, _06208_, _05407_);
  or (_25230_, _25228_, _06076_);
  or (_25231_, _25230_, _25227_);
  nand (_25232_, _06945_, _06076_);
  and (_25233_, _25232_, _12474_);
  and (_25234_, _25233_, _25231_);
  or (_25235_, _25047_, _11101_);
  nand (_25236_, _11101_, \oc8051_golden_model_1.PC [1]);
  and (_25237_, _25236_, _12473_);
  and (_25238_, _25237_, _25235_);
  or (_25239_, _25238_, _12478_);
  or (_25241_, _25239_, _25234_);
  and (_25242_, _25241_, _25043_);
  or (_25243_, _25242_, _11917_);
  or (_25244_, _11916_, _05407_);
  and (_25245_, _25244_, _07127_);
  and (_25246_, _25245_, _25243_);
  and (_25247_, _06297_, _05878_);
  or (_25248_, _25247_, _06402_);
  or (_25249_, _25248_, _25246_);
  nand (_25250_, _06402_, \oc8051_golden_model_1.PC [1]);
  and (_25252_, _25250_, _25249_);
  or (_25253_, _25252_, _12492_);
  nand (_25254_, _06945_, _12492_);
  and (_25255_, _25254_, _12497_);
  and (_25256_, _25255_, _25253_);
  or (_25257_, _25047_, _12480_);
  or (_25258_, _11101_, _05407_);
  and (_25259_, _25258_, _12496_);
  and (_25260_, _25259_, _25257_);
  or (_25261_, _25260_, _12505_);
  or (_25263_, _25261_, _25256_);
  and (_25264_, _25263_, _25041_);
  or (_25265_, _25264_, _10822_);
  or (_25266_, _10821_, _05407_);
  and (_25267_, _25266_, _07132_);
  and (_25268_, _25267_, _25265_);
  and (_25269_, _06306_, _05878_);
  or (_25270_, _25269_, _06411_);
  or (_25271_, _25270_, _25268_);
  nand (_25272_, _06411_, \oc8051_golden_model_1.PC [1]);
  and (_25274_, _25272_, _25271_);
  or (_25275_, _25274_, _07124_);
  nand (_25276_, _06945_, _07124_);
  and (_25277_, _25276_, _12518_);
  and (_25278_, _25277_, _25275_);
  or (_25279_, _25047_, \oc8051_golden_model_1.PSW [7]);
  nand (_25280_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_25281_, _25280_, _12517_);
  and (_25282_, _25281_, _25279_);
  or (_25283_, _25282_, _25278_);
  and (_25285_, _25283_, _11910_);
  nor (_25286_, _10466_, _06783_);
  and (_25287_, _11909_, _05879_);
  or (_25288_, _25287_, _25286_);
  or (_25289_, _25288_, _25285_);
  and (_25290_, _06281_, _05840_);
  and (_25291_, _25286_, _05878_);
  nor (_25292_, _25291_, _25290_);
  and (_25293_, _25292_, _25289_);
  nand (_25294_, _25290_, _05879_);
  nand (_25296_, _25294_, _10849_);
  or (_25297_, _25296_, _25293_);
  or (_25298_, _10849_, _05407_);
  and (_25299_, _25298_, _08819_);
  and (_25300_, _25299_, _25297_);
  nand (_25301_, _06303_, _05878_);
  nand (_25302_, _25301_, _12535_);
  or (_25303_, _25302_, _25300_);
  nand (_25304_, _06945_, _05842_);
  and (_25305_, _25304_, _12539_);
  or (_25307_, _05842_, _05407_);
  or (_25308_, _25307_, _08824_);
  and (_25309_, _25308_, _25305_);
  and (_25310_, _25309_, _25303_);
  or (_25311_, _25047_, _10693_);
  or (_25312_, \oc8051_golden_model_1.PSW [7], _05407_);
  and (_25313_, _25312_, _12538_);
  and (_25314_, _25313_, _25311_);
  or (_25315_, _25314_, _12547_);
  or (_25316_, _25315_, _25310_);
  and (_25318_, _25316_, _25040_);
  or (_25319_, _25318_, _10897_);
  or (_25320_, _10896_, _05407_);
  and (_25321_, _25320_, _10926_);
  and (_25322_, _25321_, _25319_);
  and (_25323_, _10925_, _05879_);
  or (_25324_, _25323_, _06417_);
  or (_25325_, _25324_, _25322_);
  or (_25326_, _09115_, _12558_);
  and (_25327_, _25326_, _25325_);
  or (_25329_, _25327_, _07142_);
  nand (_25330_, _06945_, _07142_);
  and (_25331_, _25330_, _06421_);
  and (_25332_, _25331_, _25329_);
  not (_25333_, _12682_);
  or (_25334_, _25033_, _25333_);
  or (_25335_, _12682_, _05878_);
  and (_25336_, _25335_, _06301_);
  and (_25337_, _25336_, _25334_);
  or (_25338_, _25337_, _12565_);
  or (_25340_, _25338_, _25332_);
  nand (_25341_, _25340_, _25039_);
  nand (_25342_, _25341_, _12690_);
  nor (_25343_, _12690_, _05407_);
  nor (_25344_, _25343_, _10262_);
  nand (_25345_, _25344_, _25342_);
  and (_25346_, _10262_, _05879_);
  nor (_25347_, _25346_, _06167_);
  and (_25348_, _25347_, _25345_);
  and (_25349_, _11935_, _06167_);
  or (_25351_, _25349_, _25348_);
  nand (_25352_, _25351_, _12703_);
  and (_25353_, _06945_, _05826_);
  nor (_25354_, _25353_, _06165_);
  nand (_25355_, _25354_, _25352_);
  not (_25356_, _08362_);
  and (_25357_, _25035_, _06165_);
  nor (_25358_, _25357_, _25356_);
  and (_25359_, _25358_, _25355_);
  or (_25360_, _25359_, _25038_);
  nand (_25362_, _25360_, _07154_);
  and (_25363_, _07153_, _05878_);
  nor (_25364_, _25363_, _06433_);
  and (_25365_, _25364_, _25362_);
  or (_25366_, _25365_, _25037_);
  nand (_25367_, _25366_, _12719_);
  nor (_25368_, _12719_, _05878_);
  nor (_25369_, _25368_, _07577_);
  nand (_25370_, _25369_, _25367_);
  and (_25371_, _07577_, _06945_);
  nor (_25373_, _25371_, _05748_);
  and (_25374_, _25373_, _25370_);
  or (_25375_, _25374_, _25036_);
  and (_25376_, _25375_, _09193_);
  nor (_25377_, _07168_, _05879_);
  nor (_25378_, _25377_, _12735_);
  or (_25379_, _25378_, _25376_);
  and (_25380_, _07168_, _05878_);
  nor (_25381_, _25380_, _06440_);
  and (_25382_, _25381_, _25379_);
  or (_25384_, _25382_, _25029_);
  nand (_25385_, _25384_, _12744_);
  nor (_25386_, _12744_, _05878_);
  nor (_25387_, _25386_, _25019_);
  nand (_25388_, _25387_, _25385_);
  and (_25389_, _25019_, _06945_);
  nor (_25390_, _25389_, _12754_);
  and (_25391_, _25390_, _25388_);
  and (_25392_, _12754_, _05879_);
  or (_25393_, _25392_, _25391_);
  or (_25395_, _25393_, _01321_);
  or (_25396_, _01317_, \oc8051_golden_model_1.PC [1]);
  and (_25397_, _25396_, _43100_);
  and (_43689_, _25397_, _25395_);
  and (_25398_, _06440_, _05921_);
  nor (_25399_, _11905_, _05907_);
  and (_25400_, _09070_, _06417_);
  nor (_25401_, _11907_, _05907_);
  nor (_25402_, _11912_, _05907_);
  nor (_25403_, _11914_, _05907_);
  nor (_25405_, _11919_, _05907_);
  nor (_25406_, _11922_, _05907_);
  nor (_25407_, _06131_, _05921_);
  not (_25408_, _05907_);
  and (_25409_, _11924_, _25408_);
  or (_25410_, _12028_, _11956_);
  and (_25411_, _12039_, _12036_);
  nor (_25412_, _25411_, _12040_);
  or (_25413_, _25412_, _11958_);
  nand (_25414_, _25413_, _25410_);
  nand (_25415_, _25414_, _06687_);
  and (_25416_, _06581_, _06521_);
  nor (_25417_, _12263_, _05907_);
  or (_25418_, _12265_, _25408_);
  nand (_25419_, _12266_, \oc8051_golden_model_1.PC [2]);
  and (_25420_, _25419_, _25418_);
  or (_25421_, _25420_, _07056_);
  and (_25422_, _06653_, _05907_);
  and (_25423_, _07056_, _05921_);
  nor (_25424_, _25423_, _25422_);
  and (_25427_, _25424_, _24799_);
  and (_25428_, _25427_, _25421_);
  or (_25429_, _25428_, _25417_);
  nor (_25430_, _25429_, _25416_);
  nor (_25431_, _25430_, _08445_);
  and (_25432_, _12207_, _12204_);
  nor (_25433_, _25432_, _12208_);
  nand (_25434_, _25433_, _12256_);
  or (_25435_, _12256_, _05923_);
  and (_25436_, _25435_, _08445_);
  and (_25438_, _25436_, _25434_);
  or (_25439_, _25438_, _25431_);
  nand (_25440_, _25439_, _07065_);
  and (_25441_, _07064_, _25408_);
  nor (_25442_, _25441_, _06160_);
  nand (_25443_, _25442_, _25440_);
  or (_25444_, _25412_, _12141_);
  or (_25445_, _12139_, _12028_);
  and (_25446_, _25445_, _06160_);
  nand (_25447_, _25446_, _25444_);
  and (_25449_, _25447_, _12134_);
  nand (_25450_, _25449_, _25443_);
  nor (_25451_, _12134_, _05907_);
  nor (_25452_, _25451_, _06156_);
  nand (_25453_, _25452_, _25450_);
  and (_25454_, _06156_, _05921_);
  nor (_25455_, _25454_, _07485_);
  nand (_25456_, _25455_, _25453_);
  and (_25457_, _06521_, _07485_);
  nor (_25458_, _25457_, _06217_);
  nand (_25460_, _25458_, _25456_);
  and (_25461_, _06217_, _05921_);
  nor (_25462_, _25461_, _12293_);
  nand (_25463_, _25462_, _25460_);
  nor (_25464_, _12292_, _05907_);
  nor (_25465_, _25464_, _06220_);
  nand (_25466_, _25465_, _25463_);
  and (_25467_, _06220_, _05921_);
  nor (_25468_, _25467_, _12302_);
  nand (_25469_, _25468_, _25466_);
  nor (_25471_, _12300_, _05907_);
  nor (_25472_, _25471_, _06152_);
  nand (_25473_, _25472_, _25469_);
  and (_25474_, _06152_, _05921_);
  nor (_25475_, _25474_, _12304_);
  nand (_25476_, _25475_, _25473_);
  and (_25477_, _06521_, _12304_);
  nor (_25478_, _25477_, _06151_);
  nand (_25479_, _25478_, _25476_);
  and (_25480_, _06151_, _05921_);
  nor (_25482_, _25480_, _12126_);
  and (_25483_, _25482_, _25479_);
  not (_25484_, _25412_);
  nor (_25485_, _25484_, _12120_);
  not (_25486_, _25485_);
  and (_25487_, _12120_, _12028_);
  nor (_25488_, _25487_, _12125_);
  and (_25489_, _25488_, _25486_);
  or (_25490_, _25489_, _25483_);
  nand (_25491_, _25490_, _12089_);
  nand (_25493_, _25491_, _25415_);
  nand (_25494_, _25493_, _06643_);
  and (_25495_, _12329_, _12028_);
  not (_25496_, _25495_);
  nor (_25497_, _25484_, _12329_);
  nor (_25498_, _25497_, _06643_);
  and (_25499_, _25498_, _25496_);
  nor (_25500_, _25499_, _06295_);
  nand (_25501_, _25500_, _25494_);
  nor (_25502_, _25412_, _12346_);
  and (_25504_, _12346_, _12029_);
  or (_25505_, _25504_, _12317_);
  or (_25506_, _25505_, _25502_);
  and (_25507_, _25506_, _11925_);
  and (_25508_, _25507_, _25501_);
  or (_25509_, _25508_, _25409_);
  nand (_25510_, _25509_, _06146_);
  and (_25511_, _06145_, _05923_);
  nor (_25512_, _25511_, _07388_);
  nand (_25513_, _25512_, _25510_);
  nor (_25515_, _06521_, _05760_);
  nor (_25516_, _25515_, _25152_);
  and (_25517_, _25516_, _25513_);
  nor (_25518_, _25151_, _05921_);
  or (_25519_, _25518_, _25517_);
  nand (_25520_, _25519_, _12369_);
  nor (_25521_, _12369_, _05907_);
  nor (_25522_, _25521_, _06255_);
  nand (_25523_, _25522_, _25520_);
  and (_25524_, _06255_, _05921_);
  nor (_25526_, _25524_, _24882_);
  nand (_25527_, _25526_, _25523_);
  and (_25528_, _06521_, _24882_);
  nor (_25529_, _25528_, _06254_);
  nand (_25530_, _25529_, _25527_);
  and (_25531_, _06254_, _05921_);
  nor (_25532_, _25531_, _12387_);
  and (_25533_, _25532_, _25530_);
  nor (_25534_, _12381_, _05907_);
  or (_25535_, _25534_, _25533_);
  nand (_25537_, _25535_, _12385_);
  nor (_25538_, _12385_, _05921_);
  nor (_25539_, _25538_, _05870_);
  nand (_25540_, _25539_, _25537_);
  nor (_25541_, _25408_, _05805_);
  nor (_25542_, _25541_, _06139_);
  and (_25543_, _25542_, _25540_);
  and (_25544_, _06139_, _05923_);
  or (_25545_, _25544_, _25543_);
  nand (_25546_, _25545_, _24791_);
  and (_25548_, _06521_, _05791_);
  nor (_25549_, _25548_, _06293_);
  nand (_25550_, _25549_, _25546_);
  and (_25551_, _12028_, _06293_);
  not (_25552_, _25551_);
  and (_25553_, _25552_, _06131_);
  and (_25554_, _25553_, _25550_);
  nor (_25555_, _25554_, _25407_);
  nor (_25556_, _07365_, _05797_);
  or (_25557_, _25556_, _25555_);
  and (_25559_, _25556_, _05923_);
  nor (_25560_, _25559_, _05787_);
  nand (_25561_, _25560_, _25557_);
  and (_25562_, _12028_, _05787_);
  nor (_25563_, _25562_, _12412_);
  and (_25564_, _25563_, _25561_);
  or (_25565_, _25564_, _25406_);
  and (_25566_, _25565_, _06762_);
  and (_25567_, _06209_, _05923_);
  or (_25568_, _25567_, _05829_);
  or (_25570_, _25568_, _25566_);
  nor (_25571_, _06521_, _05830_);
  nor (_25572_, _25571_, _12416_);
  and (_25573_, _25572_, _25570_);
  nor (_25574_, _25433_, _12417_);
  or (_25575_, _25574_, _25573_);
  nand (_25576_, _25575_, _07352_);
  and (_25577_, _07351_, _05923_);
  not (_25578_, _25577_);
  and (_25579_, _25578_, _08786_);
  nand (_25581_, _25579_, _25576_);
  nor (_25582_, _08786_, _05923_);
  nor (_25583_, _25582_, _06110_);
  nand (_25584_, _25583_, _25581_);
  and (_25585_, _12029_, _06110_);
  nor (_25586_, _25585_, _10751_);
  nand (_25587_, _25586_, _25584_);
  and (_25588_, _10751_, _05921_);
  nor (_25589_, _25588_, _12431_);
  nand (_25590_, _25589_, _25587_);
  and (_25592_, _12431_, _05936_);
  nor (_25593_, _25592_, _06208_);
  nand (_25594_, _25593_, _25590_);
  and (_25595_, _06208_, _05921_);
  nor (_25596_, _25595_, _06076_);
  nand (_25597_, _25596_, _25594_);
  and (_25598_, _06521_, _06076_);
  nor (_25599_, _25598_, _12473_);
  nand (_25600_, _25599_, _25597_);
  and (_25601_, _11101_, _05923_);
  nor (_25603_, _25433_, _11101_);
  or (_25604_, _25603_, _12474_);
  or (_25605_, _25604_, _25601_);
  and (_25606_, _25605_, _11919_);
  and (_25607_, _25606_, _25600_);
  or (_25608_, _25607_, _25405_);
  nand (_25609_, _25608_, _11916_);
  nor (_25610_, _11916_, _05921_);
  nor (_25611_, _25610_, _06297_);
  nand (_25612_, _25611_, _25609_);
  and (_25614_, _12028_, _06297_);
  nor (_25615_, _25614_, _06402_);
  and (_25616_, _25615_, _25612_);
  and (_25617_, _06402_, _05923_);
  or (_25618_, _25617_, _25616_);
  nand (_25619_, _25618_, _05834_);
  and (_25620_, _06521_, _12492_);
  nor (_25621_, _25620_, _12496_);
  nand (_25622_, _25621_, _25619_);
  nor (_25623_, _11101_, _05921_);
  nor (_25625_, _25433_, _12480_);
  or (_25626_, _25625_, _12497_);
  or (_25627_, _25626_, _25623_);
  and (_25628_, _25627_, _11914_);
  and (_25629_, _25628_, _25622_);
  or (_25630_, _25629_, _25403_);
  nand (_25631_, _25630_, _10821_);
  nor (_25632_, _10821_, _05921_);
  nor (_25633_, _25632_, _06306_);
  nand (_25634_, _25633_, _25631_);
  and (_25636_, _12028_, _06306_);
  nor (_25637_, _25636_, _06411_);
  and (_25638_, _25637_, _25634_);
  and (_25639_, _06411_, _05923_);
  or (_25640_, _25639_, _25638_);
  nand (_25641_, _25640_, _05848_);
  and (_25642_, _06521_, _07124_);
  nor (_25643_, _25642_, _12517_);
  nand (_25644_, _25643_, _25641_);
  nor (_25645_, _25433_, \oc8051_golden_model_1.PSW [7]);
  nor (_25647_, _05921_, _10693_);
  nor (_25648_, _25647_, _12518_);
  not (_25649_, _25648_);
  nor (_25650_, _25649_, _25645_);
  nor (_25651_, _25650_, _12522_);
  and (_25652_, _25651_, _25644_);
  or (_25653_, _25652_, _25402_);
  nand (_25654_, _25653_, _10849_);
  nor (_25655_, _10849_, _05921_);
  nor (_25656_, _25655_, _06303_);
  and (_25658_, _25656_, _25654_);
  and (_25659_, _12028_, _06303_);
  or (_25660_, _25659_, _06396_);
  nor (_25661_, _25660_, _25658_);
  and (_25662_, _06396_, _05923_);
  or (_25663_, _25662_, _25661_);
  nand (_25664_, _25663_, _05843_);
  and (_25665_, _06521_, _05842_);
  nor (_25666_, _25665_, _12538_);
  nand (_25667_, _25666_, _25664_);
  or (_25669_, _25433_, _10693_);
  or (_25670_, _05921_, \oc8051_golden_model_1.PSW [7]);
  and (_25671_, _25670_, _12538_);
  and (_25672_, _25671_, _25669_);
  nor (_25673_, _25672_, _12547_);
  and (_25674_, _25673_, _25667_);
  or (_25675_, _25674_, _25401_);
  nand (_25676_, _25675_, _10896_);
  nor (_25677_, _10896_, _05921_);
  nor (_25678_, _25677_, _10925_);
  nand (_25680_, _25678_, _25676_);
  and (_25681_, _10925_, _05907_);
  nor (_25682_, _25681_, _06417_);
  and (_25683_, _25682_, _25680_);
  or (_25684_, _25683_, _25400_);
  nand (_25685_, _25684_, _05846_);
  and (_25686_, _06521_, _07142_);
  nor (_25687_, _25686_, _06301_);
  nand (_25688_, _25687_, _25685_);
  nor (_25689_, _12028_, _12682_);
  and (_25691_, _25484_, _12682_);
  or (_25692_, _25691_, _06421_);
  nor (_25693_, _25692_, _25689_);
  nor (_25694_, _25693_, _12565_);
  and (_25695_, _25694_, _25688_);
  or (_25696_, _25695_, _25399_);
  nand (_25697_, _25696_, _12690_);
  nor (_25698_, _12690_, _05921_);
  nor (_25699_, _25698_, _10262_);
  nand (_25700_, _25699_, _25697_);
  and (_25702_, _10262_, _05907_);
  nor (_25703_, _25702_, _06167_);
  and (_25704_, _25703_, _25700_);
  and (_25705_, _09070_, _06167_);
  or (_25706_, _25705_, _25704_);
  nand (_25707_, _25706_, _12703_);
  and (_25708_, _06521_, _05826_);
  nor (_25709_, _25708_, _06165_);
  nand (_25710_, _25709_, _25707_);
  nor (_25711_, _25412_, _12682_);
  and (_25713_, _12029_, _12682_);
  nor (_25714_, _25713_, _25711_);
  and (_25715_, _25714_, _06165_);
  nor (_25716_, _25715_, _12712_);
  nand (_25717_, _25716_, _25710_);
  nor (_25718_, _12711_, _05907_);
  nor (_25719_, _25718_, _06433_);
  nand (_25720_, _25719_, _25717_);
  not (_25721_, _12719_);
  and (_25722_, _06433_, _05921_);
  nor (_25723_, _25722_, _25721_);
  and (_25724_, _25723_, _25720_);
  nor (_25725_, _12719_, _05907_);
  or (_25726_, _25725_, _25724_);
  nand (_25727_, _25726_, _07160_);
  and (_25728_, _07577_, _06521_);
  nor (_25729_, _25728_, _05748_);
  nand (_25730_, _25729_, _25727_);
  and (_25731_, _25714_, _05748_);
  nor (_25732_, _25731_, _12737_);
  nand (_25735_, _25732_, _25730_);
  nor (_25736_, _12735_, _05907_);
  nor (_25737_, _25736_, _06440_);
  and (_25738_, _25737_, _25735_);
  or (_25739_, _25738_, _25398_);
  nand (_25740_, _25739_, _12744_);
  nor (_25741_, _12744_, _25408_);
  nor (_25742_, _25741_, _25019_);
  nand (_25743_, _25742_, _25740_);
  and (_25744_, _25019_, _06521_);
  nor (_25746_, _25744_, _12754_);
  and (_25747_, _25746_, _25743_);
  and (_25748_, _12754_, _05907_);
  or (_25749_, _25748_, _25747_);
  or (_25750_, _25749_, _01321_);
  or (_25751_, _01317_, \oc8051_golden_model_1.PC [2]);
  and (_25752_, _25751_, _43100_);
  and (_43690_, _25752_, _25750_);
  and (_25753_, _06440_, _05974_);
  and (_25754_, _06433_, _05974_);
  or (_25756_, _11905_, _06324_);
  or (_25757_, _11907_, _06324_);
  or (_25758_, _11912_, _06324_);
  or (_25759_, _11914_, _06324_);
  or (_25760_, _11919_, _06324_);
  or (_25761_, _08787_, _05974_);
  or (_25762_, _25151_, _05974_);
  nand (_25763_, _11924_, _05951_);
  nor (_25764_, _06582_, _06389_);
  nand (_25765_, _07056_, _06322_);
  and (_25767_, _25765_, _12264_);
  and (_25768_, _12265_, \oc8051_golden_model_1.PC [3]);
  or (_25769_, _25768_, _07056_);
  and (_25770_, _25769_, _25767_);
  or (_25771_, _12266_, _05951_);
  nand (_25772_, _25771_, _12263_);
  or (_25773_, _25772_, _25770_);
  and (_25774_, _25773_, _06582_);
  or (_25775_, _25774_, _25764_);
  or (_25776_, _12263_, _06324_);
  and (_25778_, _25776_, _25775_);
  or (_25779_, _25778_, _08445_);
  or (_25780_, _12197_, _12196_);
  nand (_25781_, _25780_, _12209_);
  or (_25782_, _25780_, _12209_);
  and (_25783_, _25782_, _25781_);
  and (_25784_, _25783_, _12256_);
  and (_25785_, _12258_, _05974_);
  or (_25786_, _25785_, _08443_);
  or (_25787_, _25786_, _25784_);
  and (_25789_, _25787_, _25779_);
  or (_25790_, _25789_, _07064_);
  nand (_25791_, _07064_, _05951_);
  and (_25792_, _25791_, _06161_);
  and (_25793_, _25792_, _25790_);
  or (_25794_, _12139_, _12023_);
  or (_25795_, _12026_, _12025_);
  and (_25796_, _25795_, _12041_);
  nor (_25797_, _25795_, _12041_);
  nor (_25798_, _25797_, _25796_);
  or (_25800_, _25798_, _12141_);
  and (_25801_, _25800_, _06160_);
  and (_25802_, _25801_, _25794_);
  or (_25803_, _25802_, _24821_);
  or (_25804_, _25803_, _25793_);
  or (_25805_, _12134_, _06324_);
  and (_25806_, _25805_, _06157_);
  and (_25807_, _25806_, _25804_);
  and (_25808_, _06156_, _05974_);
  or (_25809_, _25808_, _07485_);
  or (_25811_, _25809_, _25807_);
  nand (_25812_, _06389_, _07485_);
  and (_25813_, _25812_, _07075_);
  and (_25814_, _25813_, _25811_);
  nand (_25815_, _06217_, _05974_);
  nand (_25816_, _25815_, _12292_);
  or (_25817_, _25816_, _25814_);
  or (_25818_, _12292_, _06324_);
  and (_25819_, _25818_, _06229_);
  and (_25820_, _25819_, _25817_);
  nand (_25822_, _06220_, _05974_);
  nand (_25823_, _25822_, _12300_);
  or (_25824_, _25823_, _25820_);
  or (_25825_, _12300_, _06324_);
  and (_25826_, _25825_, _06153_);
  and (_25827_, _25826_, _25824_);
  and (_25828_, _06152_, _05974_);
  or (_25829_, _25828_, _12304_);
  or (_25830_, _25829_, _25827_);
  nand (_25831_, _06389_, _12304_);
  and (_25833_, _25831_, _07191_);
  and (_25834_, _25833_, _25830_);
  nand (_25835_, _06151_, _05974_);
  nand (_25836_, _25835_, _12125_);
  or (_25837_, _25836_, _25834_);
  not (_25838_, _25798_);
  nor (_25839_, _25838_, _12120_);
  and (_25840_, _12120_, _12023_);
  or (_25841_, _25840_, _12125_);
  or (_25842_, _25841_, _25839_);
  and (_25844_, _25842_, _25114_);
  and (_25845_, _25844_, _25837_);
  and (_25846_, _12329_, _12023_);
  nor (_25847_, _25838_, _12329_);
  or (_25848_, _25847_, _25846_);
  and (_25849_, _25848_, _06236_);
  or (_25850_, _12023_, _11956_);
  or (_25851_, _25798_, _11958_);
  and (_25852_, _25851_, _06687_);
  and (_25853_, _25852_, _25850_);
  or (_25855_, _25853_, _25849_);
  or (_25856_, _25855_, _25845_);
  and (_25857_, _25856_, _12317_);
  nand (_25858_, _12346_, _12024_);
  or (_25859_, _25798_, _12346_);
  and (_25860_, _25859_, _06295_);
  and (_25861_, _25860_, _25858_);
  or (_25862_, _25861_, _11924_);
  or (_25863_, _25862_, _25857_);
  and (_25864_, _25863_, _25763_);
  or (_25866_, _25864_, _06145_);
  nand (_25867_, _06145_, _06322_);
  and (_25868_, _25867_, _05760_);
  and (_25869_, _25868_, _25866_);
  nor (_25870_, _06389_, _05760_);
  or (_25871_, _25870_, _25152_);
  or (_25872_, _25871_, _25869_);
  and (_25873_, _25872_, _25762_);
  or (_25874_, _25873_, _12373_);
  or (_25875_, _12369_, _06324_);
  and (_25876_, _25875_, _13844_);
  and (_25877_, _25876_, _25874_);
  and (_25878_, _06255_, _05974_);
  or (_25879_, _25878_, _24882_);
  or (_25880_, _25879_, _25877_);
  nand (_25881_, _06389_, _24882_);
  and (_25882_, _25881_, _13843_);
  and (_25883_, _25882_, _25880_);
  nand (_25884_, _06254_, _05974_);
  nand (_25885_, _25884_, _12381_);
  or (_25887_, _25885_, _25883_);
  or (_25888_, _12381_, _06324_);
  and (_25889_, _25888_, _25887_);
  or (_25890_, _25889_, _12386_);
  or (_25891_, _12385_, _05974_);
  and (_25892_, _25891_, _05805_);
  and (_25893_, _25892_, _25890_);
  nor (_25894_, _05805_, _05951_);
  or (_25895_, _25894_, _06139_);
  or (_25896_, _25895_, _25893_);
  nand (_25898_, _06139_, _06322_);
  and (_25899_, _25898_, _25896_);
  or (_25900_, _25899_, _05791_);
  nand (_25901_, _06389_, _05791_);
  and (_25902_, _25901_, _11296_);
  and (_25903_, _25902_, _25900_);
  nand (_25904_, _12023_, _06293_);
  nand (_25905_, _25904_, _06133_);
  or (_25906_, _25905_, _25903_);
  or (_25907_, _06133_, _05974_);
  and (_25908_, _25907_, _06114_);
  and (_25909_, _25908_, _25906_);
  nand (_25910_, _12023_, _05787_);
  nand (_25911_, _25910_, _11922_);
  or (_25912_, _25911_, _25909_);
  or (_25913_, _11922_, _06324_);
  and (_25914_, _25913_, _06762_);
  and (_25915_, _25914_, _25912_);
  and (_25916_, _06209_, _05974_);
  or (_25917_, _25916_, _05829_);
  or (_25918_, _25917_, _25915_);
  nand (_25919_, _06389_, _05829_);
  and (_25920_, _25919_, _12417_);
  and (_25921_, _25920_, _25918_);
  and (_25922_, _25783_, _12416_);
  or (_25923_, _25922_, _08788_);
  or (_25924_, _25923_, _25921_);
  and (_25925_, _25924_, _25761_);
  or (_25926_, _25925_, _06110_);
  nand (_25927_, _12024_, _06110_);
  and (_25928_, _25927_, _10752_);
  and (_25929_, _25928_, _25926_);
  and (_25930_, _10751_, _05974_);
  or (_25931_, _25930_, _12431_);
  or (_25932_, _25931_, _25929_);
  or (_25933_, _12432_, _05968_);
  and (_25934_, _25933_, _06768_);
  and (_25935_, _25934_, _25932_);
  and (_25936_, _06208_, _05974_);
  or (_25937_, _25936_, _06076_);
  or (_25938_, _25937_, _25935_);
  nand (_25939_, _06389_, _06076_);
  and (_25940_, _25939_, _12474_);
  and (_25941_, _25940_, _25938_);
  or (_25942_, _25783_, _11101_);
  nand (_25943_, _11101_, _06322_);
  and (_25944_, _25943_, _12473_);
  and (_25945_, _25944_, _25942_);
  or (_25946_, _25945_, _12478_);
  or (_25947_, _25946_, _25941_);
  and (_25948_, _25947_, _25760_);
  or (_25949_, _25948_, _11917_);
  or (_25950_, _11916_, _05974_);
  and (_25951_, _25950_, _07127_);
  and (_25952_, _25951_, _25949_);
  and (_25953_, _12023_, _06297_);
  or (_25954_, _25953_, _06402_);
  or (_25955_, _25954_, _25952_);
  nand (_25956_, _06402_, _06322_);
  and (_25957_, _25956_, _25955_);
  or (_25959_, _25957_, _12492_);
  nand (_25960_, _06389_, _12492_);
  and (_25961_, _25960_, _12497_);
  and (_25962_, _25961_, _25959_);
  or (_25963_, _25783_, _12480_);
  or (_25964_, _11101_, _05974_);
  and (_25965_, _25964_, _12496_);
  and (_25966_, _25965_, _25963_);
  or (_25967_, _25966_, _12505_);
  or (_25968_, _25967_, _25962_);
  and (_25970_, _25968_, _25759_);
  or (_25971_, _25970_, _10822_);
  or (_25972_, _10821_, _05974_);
  and (_25973_, _25972_, _07132_);
  and (_25974_, _25973_, _25971_);
  and (_25975_, _12023_, _06306_);
  or (_25976_, _25975_, _06411_);
  or (_25977_, _25976_, _25974_);
  nand (_25978_, _06411_, _06322_);
  and (_25979_, _25978_, _25977_);
  or (_25980_, _25979_, _07124_);
  nand (_25981_, _06389_, _07124_);
  and (_25982_, _25981_, _12518_);
  and (_25983_, _25982_, _25980_);
  or (_25984_, _25783_, \oc8051_golden_model_1.PSW [7]);
  or (_25985_, _05974_, _10693_);
  and (_25986_, _25985_, _12517_);
  and (_25987_, _25986_, _25984_);
  or (_25988_, _25987_, _12522_);
  or (_25989_, _25988_, _25983_);
  and (_25991_, _25989_, _25758_);
  or (_25992_, _25991_, _10850_);
  or (_25993_, _10849_, _05974_);
  and (_25994_, _25993_, _08819_);
  and (_25995_, _25994_, _25992_);
  and (_25996_, _12023_, _06303_);
  or (_25997_, _25996_, _06396_);
  or (_25998_, _25997_, _25995_);
  nand (_25999_, _06396_, _06322_);
  and (_26000_, _25999_, _25998_);
  or (_26002_, _26000_, _05842_);
  nand (_26003_, _06389_, _05842_);
  and (_26004_, _26003_, _12539_);
  and (_26005_, _26004_, _26002_);
  or (_26006_, _25783_, _10693_);
  or (_26007_, _05974_, \oc8051_golden_model_1.PSW [7]);
  and (_26008_, _26007_, _12538_);
  and (_26009_, _26008_, _26006_);
  or (_26010_, _26009_, _12547_);
  or (_26011_, _26010_, _26005_);
  and (_26013_, _26011_, _25757_);
  or (_26014_, _26013_, _10897_);
  or (_26015_, _10896_, _05974_);
  and (_26016_, _26015_, _10926_);
  and (_26017_, _26016_, _26014_);
  and (_26018_, _10925_, _06324_);
  or (_26019_, _26018_, _06417_);
  or (_26020_, _26019_, _26017_);
  or (_26021_, _09210_, _12558_);
  and (_26022_, _26021_, _26020_);
  or (_26024_, _26022_, _07142_);
  nand (_26025_, _06389_, _07142_);
  and (_26026_, _26025_, _06421_);
  and (_26027_, _26026_, _26024_);
  or (_26028_, _12023_, _12682_);
  nand (_26029_, _25838_, _12682_);
  and (_26030_, _26029_, _06301_);
  and (_26031_, _26030_, _26028_);
  or (_26032_, _26031_, _12565_);
  or (_26033_, _26032_, _26027_);
  and (_26034_, _26033_, _25756_);
  or (_26035_, _26034_, _12691_);
  or (_26036_, _12690_, _05974_);
  and (_26037_, _26036_, _12693_);
  and (_26038_, _26037_, _26035_);
  and (_26039_, _10262_, _06324_);
  or (_26040_, _26039_, _06167_);
  or (_26041_, _26040_, _26038_);
  or (_26042_, _09210_, _06168_);
  and (_26043_, _26042_, _26041_);
  or (_26044_, _26043_, _05826_);
  nand (_26045_, _06389_, _05826_);
  and (_26046_, _26045_, _06166_);
  and (_26047_, _26046_, _26044_);
  nor (_26048_, _25798_, _12682_);
  and (_26049_, _12024_, _12682_);
  nor (_26050_, _26049_, _26048_);
  and (_26051_, _26050_, _06165_);
  or (_26052_, _26051_, _12712_);
  or (_26053_, _26052_, _26047_);
  or (_26056_, _12711_, _06324_);
  and (_26057_, _26056_, _06829_);
  and (_26058_, _26057_, _26053_);
  or (_26059_, _26058_, _25754_);
  nand (_26060_, _26059_, _12719_);
  nor (_26061_, _12719_, _05951_);
  nor (_26062_, _26061_, _07577_);
  nand (_26063_, _26062_, _26060_);
  and (_26064_, _07577_, _06389_);
  nor (_26065_, _26064_, _05748_);
  nand (_26067_, _26065_, _26063_);
  and (_26068_, _26050_, _05748_);
  nor (_26069_, _26068_, _12737_);
  nand (_26070_, _26069_, _26067_);
  nor (_26071_, _12735_, _06324_);
  nor (_26072_, _26071_, _06440_);
  and (_26073_, _26072_, _26070_);
  or (_26074_, _26073_, _25753_);
  nand (_26075_, _26074_, _12744_);
  nor (_26076_, _12744_, _05951_);
  nor (_26078_, _26076_, _25019_);
  nand (_26079_, _26078_, _26075_);
  and (_26080_, _25019_, _06389_);
  nor (_26081_, _26080_, _12754_);
  and (_26082_, _26081_, _26079_);
  and (_26083_, _12754_, _06324_);
  or (_26084_, _26083_, _26082_);
  or (_26085_, _26084_, _01321_);
  or (_26086_, _01317_, \oc8051_golden_model_1.PC [3]);
  and (_26087_, _26086_, _43100_);
  and (_43691_, _26087_, _26085_);
  and (_26089_, _08670_, _07577_);
  nor (_26090_, _12194_, _11101_);
  and (_26091_, _12214_, _12211_);
  nor (_26092_, _26091_, _12215_);
  and (_26093_, _26092_, _11101_);
  or (_26094_, _26093_, _26090_);
  and (_26095_, _26094_, _12496_);
  and (_26096_, _12193_, _11101_);
  and (_26097_, _26092_, _12480_);
  or (_26098_, _26097_, _26096_);
  and (_26099_, _26098_, _12473_);
  nor (_26100_, _12193_, _08787_);
  nor (_26101_, _25151_, _12193_);
  and (_26102_, _05426_, \oc8051_golden_model_1.PC [4]);
  nor (_26103_, _05426_, \oc8051_golden_model_1.PC [4]);
  nor (_26104_, _26103_, _26102_);
  not (_26105_, _26104_);
  and (_26106_, _26105_, _11924_);
  nand (_26107_, _26105_, _12287_);
  and (_26109_, _12046_, _12043_);
  nor (_26110_, _26109_, _12047_);
  or (_26111_, _26110_, _12141_);
  or (_26112_, _12139_, _12018_);
  and (_26113_, _26112_, _26111_);
  or (_26114_, _26113_, _06161_);
  and (_26115_, _08670_, _06581_);
  and (_26116_, _12194_, _07056_);
  or (_26117_, _26116_, _06653_);
  nand (_26118_, _12265_, \oc8051_golden_model_1.PC [4]);
  and (_26120_, _26118_, _07057_);
  or (_26121_, _26120_, _26117_);
  or (_26122_, _26105_, _12266_);
  and (_26123_, _26122_, _06582_);
  and (_26124_, _26123_, _26121_);
  or (_26125_, _26124_, _25055_);
  or (_26126_, _26125_, _26115_);
  or (_26127_, _26105_, _12263_);
  and (_26128_, _26127_, _08443_);
  and (_26129_, _26128_, _26126_);
  or (_26131_, _12256_, _12194_);
  nand (_26132_, _26092_, _12256_);
  and (_26133_, _26132_, _08445_);
  and (_26134_, _26133_, _26131_);
  or (_26135_, _26134_, _26129_);
  nand (_26136_, _26135_, _12281_);
  and (_26137_, _26136_, _26114_);
  or (_26138_, _26137_, _24821_);
  nand (_26139_, _26138_, _26107_);
  nand (_26140_, _26139_, _06157_);
  and (_26142_, _12194_, _06156_);
  nor (_26143_, _26142_, _07485_);
  nand (_26144_, _26143_, _26140_);
  nor (_26145_, _08670_, _05764_);
  nor (_26146_, _26145_, _06217_);
  and (_26147_, _26146_, _26144_);
  and (_26148_, _12194_, _06217_);
  or (_26149_, _26148_, _26147_);
  and (_26150_, _26149_, _12292_);
  nor (_26151_, _26104_, _12292_);
  or (_26153_, _26151_, _26150_);
  nand (_26154_, _26153_, _06229_);
  and (_26155_, _12194_, _06220_);
  nor (_26156_, _26155_, _12302_);
  nand (_26157_, _26156_, _26154_);
  nor (_26158_, _26105_, _12300_);
  nor (_26159_, _26158_, _06152_);
  and (_26160_, _26159_, _26157_);
  and (_26161_, _12194_, _06152_);
  or (_26162_, _26161_, _26160_);
  nand (_26163_, _26162_, _05769_);
  and (_26164_, _08670_, _12304_);
  nor (_26165_, _26164_, _06151_);
  nand (_26166_, _26165_, _26163_);
  and (_26167_, _12193_, _06151_);
  nor (_26168_, _26167_, _12126_);
  nand (_26169_, _26168_, _26166_);
  and (_26170_, _12120_, _12018_);
  not (_26171_, _26110_);
  nor (_26172_, _26171_, _12120_);
  or (_26174_, _26172_, _12125_);
  nor (_26175_, _26174_, _26170_);
  not (_26176_, _26175_);
  and (_26177_, _26176_, _26169_);
  or (_26178_, _26177_, _06687_);
  and (_26179_, _26110_, _11956_);
  and (_26180_, _12018_, _11958_);
  or (_26181_, _26180_, _12089_);
  or (_26182_, _26181_, _26179_);
  nand (_26183_, _26182_, _26178_);
  nand (_26185_, _26183_, _06643_);
  nor (_26186_, _26171_, _12329_);
  not (_26187_, _26186_);
  and (_26188_, _12329_, _12018_);
  nor (_26189_, _26188_, _06643_);
  and (_26190_, _26189_, _26187_);
  nor (_26191_, _26190_, _06295_);
  nand (_26192_, _26191_, _26185_);
  nor (_26193_, _26110_, _12346_);
  and (_26194_, _12346_, _12019_);
  nor (_26196_, _26194_, _12317_);
  not (_26197_, _26196_);
  nor (_26198_, _26197_, _26193_);
  nor (_26199_, _26198_, _11924_);
  and (_26200_, _26199_, _26192_);
  or (_26201_, _26200_, _26106_);
  nand (_26202_, _26201_, _06146_);
  and (_26203_, _12194_, _06145_);
  nor (_26204_, _26203_, _07388_);
  nand (_26205_, _26204_, _26202_);
  nor (_26207_, _08670_, _05760_);
  nor (_26208_, _26207_, _25152_);
  and (_26209_, _26208_, _26205_);
  or (_26210_, _26209_, _26101_);
  nand (_26211_, _26210_, _12369_);
  nor (_26212_, _26104_, _12369_);
  nor (_26213_, _26212_, _06255_);
  nand (_26214_, _26213_, _26211_);
  and (_26215_, _12193_, _06255_);
  nor (_26216_, _26215_, _24882_);
  nand (_26218_, _26216_, _26214_);
  and (_26219_, _08670_, _24882_);
  nor (_26220_, _26219_, _06254_);
  and (_26221_, _26220_, _26218_);
  and (_26222_, _12193_, _06254_);
  or (_26223_, _26222_, _26221_);
  nand (_26224_, _26223_, _12381_);
  nor (_26225_, _26105_, _12381_);
  nor (_26226_, _26225_, _12386_);
  nand (_26227_, _26226_, _26224_);
  nor (_26228_, _12193_, _12385_);
  nor (_26229_, _26228_, _05870_);
  nand (_26230_, _26229_, _26227_);
  nor (_26231_, _26105_, _05805_);
  nor (_26232_, _26231_, _06139_);
  and (_26233_, _26232_, _26230_);
  and (_26234_, _12194_, _06139_);
  or (_26235_, _26234_, _26233_);
  nand (_26236_, _26235_, _24791_);
  and (_26237_, _08670_, _05791_);
  nor (_26239_, _26237_, _06293_);
  nand (_26240_, _26239_, _26236_);
  and (_26241_, _12018_, _06293_);
  nor (_26242_, _26241_, _13620_);
  nand (_26243_, _26242_, _26240_);
  nor (_26244_, _12193_, _06133_);
  nor (_26245_, _26244_, _05787_);
  nand (_26246_, _26245_, _26243_);
  and (_26247_, _12018_, _05787_);
  nor (_26248_, _26247_, _12412_);
  nand (_26250_, _26248_, _26246_);
  nor (_26251_, _26104_, _11922_);
  nor (_26252_, _26251_, _06209_);
  nand (_26253_, _26252_, _26250_);
  and (_26254_, _12193_, _06209_);
  nor (_26255_, _26254_, _05829_);
  nand (_26256_, _26255_, _26253_);
  and (_26257_, _08670_, _05829_);
  nor (_26258_, _26257_, _12416_);
  nand (_26259_, _26258_, _26256_);
  and (_26261_, _26092_, _12416_);
  nor (_26262_, _26261_, _08788_);
  and (_26263_, _26262_, _26259_);
  or (_26264_, _26263_, _26100_);
  nand (_26265_, _26264_, _06111_);
  and (_26266_, _12019_, _06110_);
  nor (_26267_, _26266_, _10751_);
  nand (_26268_, _26267_, _26265_);
  and (_26269_, _12193_, _10751_);
  nor (_26270_, _26269_, _12431_);
  nand (_26272_, _26270_, _26268_);
  and (_26273_, _12449_, _12446_);
  nor (_26274_, _26273_, _12450_);
  nor (_26275_, _26274_, _12432_);
  nor (_26276_, _26275_, _06208_);
  nand (_26277_, _26276_, _26272_);
  and (_26278_, _12193_, _06208_);
  nor (_26279_, _26278_, _06076_);
  nand (_26280_, _26279_, _26277_);
  and (_26281_, _08670_, _06076_);
  nor (_26283_, _26281_, _12473_);
  and (_26284_, _26283_, _26280_);
  or (_26285_, _26284_, _26099_);
  nand (_26286_, _26285_, _11919_);
  nor (_26287_, _26105_, _11919_);
  nor (_26288_, _26287_, _11917_);
  nand (_26289_, _26288_, _26286_);
  nor (_26290_, _12193_, _11916_);
  nor (_26291_, _26290_, _06297_);
  nand (_26292_, _26291_, _26289_);
  and (_26293_, _12018_, _06297_);
  nor (_26294_, _26293_, _06402_);
  and (_26295_, _26294_, _26292_);
  and (_26296_, _12194_, _06402_);
  or (_26297_, _26296_, _26295_);
  nand (_26298_, _26297_, _05834_);
  and (_26299_, _08670_, _12492_);
  nor (_26300_, _26299_, _12496_);
  and (_26301_, _26300_, _26298_);
  or (_26302_, _26301_, _26095_);
  nand (_26304_, _26302_, _11914_);
  nor (_26305_, _26105_, _11914_);
  nor (_26306_, _26305_, _10822_);
  nand (_26307_, _26306_, _26304_);
  nor (_26308_, _12193_, _10821_);
  nor (_26309_, _26308_, _06306_);
  nand (_26310_, _26309_, _26307_);
  and (_26311_, _12018_, _06306_);
  nor (_26312_, _26311_, _06411_);
  and (_26313_, _26312_, _26310_);
  and (_26315_, _12194_, _06411_);
  or (_26316_, _26315_, _26313_);
  nand (_26317_, _26316_, _05848_);
  and (_26318_, _08670_, _07124_);
  nor (_26319_, _26318_, _12517_);
  and (_26320_, _26319_, _26317_);
  and (_26321_, _12193_, \oc8051_golden_model_1.PSW [7]);
  and (_26322_, _26092_, _10693_);
  or (_26323_, _26322_, _26321_);
  and (_26324_, _26323_, _12517_);
  or (_26326_, _26324_, _26320_);
  nand (_26327_, _26326_, _11912_);
  nor (_26328_, _26105_, _11912_);
  nor (_26329_, _26328_, _10850_);
  nand (_26330_, _26329_, _26327_);
  nor (_26331_, _12193_, _10849_);
  nor (_26332_, _26331_, _06303_);
  nand (_26333_, _26332_, _26330_);
  and (_26334_, _12018_, _06303_);
  nor (_26335_, _26334_, _06396_);
  and (_26337_, _26335_, _26333_);
  and (_26338_, _12194_, _06396_);
  or (_26339_, _26338_, _26337_);
  nand (_26340_, _26339_, _05843_);
  and (_26341_, _08670_, _05842_);
  nor (_26342_, _26341_, _12538_);
  and (_26343_, _26342_, _26340_);
  and (_26344_, _12193_, _10693_);
  and (_26345_, _26092_, \oc8051_golden_model_1.PSW [7]);
  or (_26346_, _26345_, _26344_);
  and (_26348_, _26346_, _12538_);
  or (_26349_, _26348_, _26343_);
  nand (_26350_, _26349_, _11907_);
  nor (_26351_, _26105_, _11907_);
  nor (_26352_, _26351_, _10897_);
  nand (_26353_, _26352_, _26350_);
  nor (_26354_, _12193_, _10896_);
  nor (_26355_, _26354_, _10925_);
  nand (_26356_, _26355_, _26353_);
  and (_26357_, _26104_, _10925_);
  nor (_26359_, _26357_, _06417_);
  and (_26360_, _26359_, _26356_);
  and (_26361_, _08980_, _06417_);
  or (_26362_, _26361_, _26360_);
  nand (_26363_, _26362_, _05846_);
  and (_26364_, _08670_, _07142_);
  nor (_26365_, _26364_, _06301_);
  and (_26366_, _26365_, _26363_);
  nor (_26367_, _12019_, _12682_);
  and (_26368_, _26110_, _12682_);
  nor (_26370_, _26368_, _26367_);
  nor (_26371_, _26370_, _06421_);
  or (_26372_, _26371_, _26366_);
  nand (_26373_, _26372_, _11905_);
  nor (_26374_, _26105_, _11905_);
  nor (_26375_, _26374_, _12691_);
  nand (_26376_, _26375_, _26373_);
  nor (_26377_, _12690_, _12193_);
  nor (_26378_, _26377_, _10262_);
  nand (_26379_, _26378_, _26376_);
  and (_26380_, _26104_, _10262_);
  nor (_26381_, _26380_, _06167_);
  nand (_26382_, _26381_, _26379_);
  and (_26383_, _08980_, _06167_);
  nor (_26384_, _26383_, _05826_);
  nand (_26385_, _26384_, _26382_);
  nor (_26386_, _08670_, _12703_);
  nor (_26387_, _26386_, _06165_);
  nand (_26388_, _26387_, _26385_);
  and (_26389_, _12019_, _12682_);
  nor (_26391_, _26110_, _12682_);
  nor (_26392_, _26391_, _26389_);
  nor (_26393_, _26392_, _06166_);
  nor (_26394_, _26393_, _12712_);
  nand (_26395_, _26394_, _26388_);
  nor (_26396_, _26105_, _12711_);
  nor (_26397_, _26396_, _06433_);
  nand (_26398_, _26397_, _26395_);
  and (_26399_, _12194_, _06433_);
  nor (_26400_, _26399_, _25721_);
  nand (_26402_, _26400_, _26398_);
  nor (_26403_, _26105_, _12719_);
  nor (_26404_, _26403_, _07577_);
  and (_26405_, _26404_, _26402_);
  or (_26406_, _26405_, _26089_);
  nand (_26407_, _26406_, _05749_);
  nor (_26408_, _26392_, _05749_);
  nor (_26409_, _26408_, _12737_);
  nand (_26410_, _26409_, _26407_);
  nor (_26411_, _26105_, _12735_);
  nor (_26413_, _26411_, _06440_);
  nand (_26414_, _26413_, _26410_);
  not (_26415_, _12744_);
  and (_26416_, _12194_, _06440_);
  nor (_26417_, _26416_, _26415_);
  nand (_26418_, _26417_, _26414_);
  nor (_26419_, _26105_, _12744_);
  nor (_26420_, _26419_, _25019_);
  nand (_26421_, _26420_, _26418_);
  and (_26422_, _25019_, _08670_);
  nor (_26424_, _26422_, _12754_);
  and (_26425_, _26424_, _26421_);
  and (_26426_, _26104_, _12754_);
  or (_26427_, _26426_, _26425_);
  or (_26428_, _26427_, _01321_);
  or (_26429_, _01317_, \oc8051_golden_model_1.PC [4]);
  and (_26430_, _26429_, _43100_);
  and (_43692_, _26430_, _26428_);
  and (_26431_, _12188_, _06440_);
  and (_26432_, _12188_, _06433_);
  nor (_26434_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_26435_, _12188_, _05444_);
  nor (_26436_, _26435_, _26434_);
  nor (_26437_, _26436_, _11905_);
  and (_26438_, _08931_, _06417_);
  nor (_26439_, _26436_, _11907_);
  nor (_26440_, _26436_, _11912_);
  nor (_26441_, _26436_, _11914_);
  nor (_26442_, _26436_, _11919_);
  nor (_26443_, _12188_, _08787_);
  nor (_26444_, _25151_, _12188_);
  not (_26445_, _26436_);
  and (_26446_, _26445_, _11924_);
  nor (_26447_, _08701_, _06582_);
  and (_26448_, _12189_, _07056_);
  nor (_26449_, _26448_, _06653_);
  and (_26450_, _12265_, \oc8051_golden_model_1.PC [5]);
  or (_26451_, _26450_, _07056_);
  and (_26452_, _26451_, _26449_);
  or (_26453_, _26445_, _12266_);
  nand (_26455_, _26453_, _12263_);
  or (_26456_, _26455_, _26452_);
  and (_26457_, _26456_, _06582_);
  nor (_26458_, _26457_, _26447_);
  nor (_26459_, _26436_, _12263_);
  nor (_26460_, _26459_, _26458_);
  nor (_26461_, _26460_, _08445_);
  or (_26462_, _12256_, _12189_);
  or (_26463_, _12191_, _12190_);
  and (_26464_, _26463_, _12216_);
  nor (_26466_, _26463_, _12216_);
  or (_26467_, _26466_, _26464_);
  or (_26468_, _26467_, _12258_);
  and (_26469_, _26468_, _08445_);
  and (_26470_, _26469_, _26462_);
  or (_26471_, _26470_, _26461_);
  nand (_26472_, _26471_, _07065_);
  and (_26473_, _26445_, _07064_);
  nor (_26474_, _26473_, _06160_);
  and (_26475_, _26474_, _26472_);
  or (_26477_, _12139_, _12014_);
  or (_26478_, _12016_, _12015_);
  not (_26479_, _26478_);
  nor (_26480_, _26479_, _12048_);
  and (_26481_, _26479_, _12048_);
  nor (_26482_, _26481_, _26480_);
  or (_26483_, _26482_, _12141_);
  nand (_26484_, _26483_, _26477_);
  and (_26485_, _26484_, _06160_);
  or (_26486_, _26485_, _24821_);
  or (_26488_, _26486_, _26475_);
  nor (_26489_, _26436_, _12134_);
  nor (_26490_, _26489_, _06156_);
  nand (_26491_, _26490_, _26488_);
  and (_26492_, _12188_, _06156_);
  nor (_26493_, _26492_, _07485_);
  nand (_26494_, _26493_, _26491_);
  and (_26495_, _08701_, _07485_);
  nor (_26496_, _26495_, _06217_);
  nand (_26497_, _26496_, _26494_);
  and (_26499_, _12188_, _06217_);
  nor (_26500_, _26499_, _12293_);
  nand (_26501_, _26500_, _26497_);
  nor (_26502_, _26436_, _12292_);
  nor (_26503_, _26502_, _06220_);
  nand (_26504_, _26503_, _26501_);
  and (_26505_, _12188_, _06220_);
  nor (_26506_, _26505_, _12302_);
  nand (_26507_, _26506_, _26504_);
  nor (_26508_, _26436_, _12300_);
  nor (_26510_, _26508_, _06152_);
  nand (_26511_, _26510_, _26507_);
  and (_26512_, _12188_, _06152_);
  nor (_26513_, _26512_, _12304_);
  nand (_26514_, _26513_, _26511_);
  and (_26515_, _08701_, _12304_);
  nor (_26516_, _26515_, _06151_);
  nand (_26517_, _26516_, _26514_);
  and (_26518_, _12188_, _06151_);
  nor (_26519_, _26518_, _12126_);
  nand (_26520_, _26519_, _26517_);
  and (_26521_, _12120_, _12013_);
  nor (_26522_, _26482_, _12120_);
  or (_26523_, _26522_, _12125_);
  nor (_26524_, _26523_, _26521_);
  not (_26525_, _26524_);
  and (_26526_, _26525_, _26520_);
  or (_26527_, _26526_, _06687_);
  and (_26528_, _12013_, _11958_);
  not (_26529_, _26482_);
  and (_26532_, _26529_, _11956_);
  or (_26533_, _26532_, _12089_);
  or (_26534_, _26533_, _26528_);
  nand (_26535_, _26534_, _26527_);
  or (_26536_, _26535_, _06236_);
  nor (_26537_, _26482_, _12329_);
  and (_26538_, _12329_, _12013_);
  nor (_26539_, _26538_, _26537_);
  or (_26540_, _26539_, _06643_);
  and (_26541_, _26540_, _26536_);
  or (_26543_, _26541_, _06295_);
  and (_26544_, _12346_, _12013_);
  nor (_26545_, _26482_, _12346_);
  nor (_26546_, _26545_, _26544_);
  nor (_26547_, _26546_, _12317_);
  nor (_26548_, _26547_, _11924_);
  and (_26549_, _26548_, _26543_);
  or (_26550_, _26549_, _26446_);
  nand (_26551_, _26550_, _06146_);
  and (_26552_, _12189_, _06145_);
  nor (_26554_, _26552_, _07388_);
  nand (_26555_, _26554_, _26551_);
  nor (_26556_, _08701_, _05760_);
  nor (_26557_, _26556_, _25152_);
  and (_26558_, _26557_, _26555_);
  or (_26559_, _26558_, _26444_);
  nand (_26560_, _26559_, _12369_);
  nor (_26561_, _26436_, _12369_);
  nor (_26562_, _26561_, _06255_);
  nand (_26563_, _26562_, _26560_);
  and (_26565_, _12188_, _06255_);
  nor (_26566_, _26565_, _24882_);
  nand (_26567_, _26566_, _26563_);
  and (_26568_, _08701_, _24882_);
  nor (_26569_, _26568_, _06254_);
  nand (_26570_, _26569_, _26567_);
  and (_26571_, _12188_, _06254_);
  nor (_26572_, _26571_, _12387_);
  and (_26573_, _26572_, _26570_);
  nor (_26574_, _26436_, _12381_);
  or (_26576_, _26574_, _26573_);
  nand (_26577_, _26576_, _12385_);
  nor (_26578_, _12188_, _12385_);
  nor (_26579_, _26578_, _05870_);
  nand (_26580_, _26579_, _26577_);
  nor (_26581_, _26445_, _05805_);
  nor (_26582_, _26581_, _06139_);
  and (_26583_, _26582_, _26580_);
  and (_26584_, _12189_, _06139_);
  or (_26585_, _26584_, _26583_);
  nand (_26587_, _26585_, _24791_);
  and (_26588_, _08701_, _05791_);
  nor (_26589_, _26588_, _06293_);
  nand (_26590_, _26589_, _26587_);
  and (_26591_, _12013_, _06293_);
  nor (_26592_, _26591_, _13620_);
  nand (_26593_, _26592_, _26590_);
  nor (_26594_, _12188_, _06133_);
  nor (_26595_, _26594_, _05787_);
  nand (_26596_, _26595_, _26593_);
  and (_26598_, _12013_, _05787_);
  nor (_26599_, _26598_, _12412_);
  nand (_26600_, _26599_, _26596_);
  nor (_26601_, _26436_, _11922_);
  nor (_26602_, _26601_, _06209_);
  nand (_26603_, _26602_, _26600_);
  and (_26604_, _12188_, _06209_);
  nor (_26605_, _26604_, _05829_);
  nand (_26606_, _26605_, _26603_);
  and (_26607_, _08701_, _05829_);
  nor (_26609_, _26607_, _12416_);
  nand (_26610_, _26609_, _26606_);
  nor (_26611_, _26467_, _12417_);
  nor (_26612_, _26611_, _08788_);
  and (_26613_, _26612_, _26610_);
  or (_26614_, _26613_, _26443_);
  nand (_26615_, _26614_, _06111_);
  and (_26616_, _12014_, _06110_);
  nor (_26617_, _26616_, _10751_);
  nand (_26618_, _26617_, _26615_);
  and (_26620_, _12188_, _10751_);
  nor (_26621_, _26620_, _12431_);
  nand (_26622_, _26621_, _26618_);
  and (_26623_, _12451_, _12444_);
  nor (_26624_, _26623_, _12452_);
  nor (_26625_, _26624_, _12432_);
  nor (_26626_, _26625_, _06208_);
  nand (_26627_, _26626_, _26622_);
  and (_26628_, _12188_, _06208_);
  nor (_26629_, _26628_, _06076_);
  nand (_26631_, _26629_, _26627_);
  and (_26632_, _08701_, _06076_);
  nor (_26633_, _26632_, _12473_);
  nand (_26634_, _26633_, _26631_);
  and (_26635_, _12188_, _11101_);
  nor (_26636_, _26467_, _11101_);
  or (_26637_, _26636_, _26635_);
  and (_26638_, _26637_, _12473_);
  nor (_26639_, _26638_, _12478_);
  and (_26640_, _26639_, _26634_);
  or (_26642_, _26640_, _26442_);
  nand (_26643_, _26642_, _11916_);
  nor (_26644_, _12188_, _11916_);
  nor (_26645_, _26644_, _06297_);
  nand (_26646_, _26645_, _26643_);
  and (_26647_, _12013_, _06297_);
  nor (_26648_, _26647_, _06402_);
  and (_26649_, _26648_, _26646_);
  and (_26650_, _12189_, _06402_);
  or (_26651_, _26650_, _26649_);
  nand (_26653_, _26651_, _05834_);
  and (_26654_, _08701_, _12492_);
  nor (_26655_, _26654_, _12496_);
  nand (_26656_, _26655_, _26653_);
  and (_26657_, _26467_, _11101_);
  nor (_26658_, _12188_, _11101_);
  nor (_26659_, _26658_, _12497_);
  not (_26660_, _26659_);
  nor (_26661_, _26660_, _26657_);
  nor (_26662_, _26661_, _12505_);
  and (_26664_, _26662_, _26656_);
  or (_26665_, _26664_, _26441_);
  nand (_26666_, _26665_, _10821_);
  nor (_26667_, _12188_, _10821_);
  nor (_26668_, _26667_, _06306_);
  nand (_26669_, _26668_, _26666_);
  and (_26670_, _12013_, _06306_);
  nor (_26671_, _26670_, _06411_);
  and (_26672_, _26671_, _26669_);
  and (_26673_, _12189_, _06411_);
  or (_26675_, _26673_, _26672_);
  nand (_26676_, _26675_, _05848_);
  and (_26677_, _08701_, _07124_);
  nor (_26678_, _26677_, _12517_);
  nand (_26679_, _26678_, _26676_);
  and (_26680_, _12188_, \oc8051_golden_model_1.PSW [7]);
  nor (_26681_, _26467_, \oc8051_golden_model_1.PSW [7]);
  or (_26682_, _26681_, _26680_);
  and (_26683_, _26682_, _12517_);
  nor (_26684_, _26683_, _12522_);
  and (_26686_, _26684_, _26679_);
  or (_26687_, _26686_, _26440_);
  nand (_26688_, _26687_, _10849_);
  nor (_26689_, _12188_, _10849_);
  nor (_26690_, _26689_, _06303_);
  nand (_26691_, _26690_, _26688_);
  and (_26692_, _12013_, _06303_);
  nor (_26693_, _26692_, _06396_);
  and (_26694_, _26693_, _26691_);
  and (_26695_, _12189_, _06396_);
  or (_26697_, _26695_, _26694_);
  nand (_26698_, _26697_, _05843_);
  and (_26699_, _08701_, _05842_);
  nor (_26700_, _26699_, _12538_);
  nand (_26701_, _26700_, _26698_);
  nand (_26702_, _26467_, \oc8051_golden_model_1.PSW [7]);
  or (_26703_, _12188_, \oc8051_golden_model_1.PSW [7]);
  and (_26704_, _26703_, _12538_);
  and (_26705_, _26704_, _26702_);
  nor (_26706_, _26705_, _12547_);
  and (_26708_, _26706_, _26701_);
  or (_26709_, _26708_, _26439_);
  nand (_26710_, _26709_, _10896_);
  nor (_26711_, _12188_, _10896_);
  nor (_26712_, _26711_, _10925_);
  nand (_26713_, _26712_, _26710_);
  and (_26714_, _26436_, _10925_);
  nor (_26715_, _26714_, _06417_);
  and (_26716_, _26715_, _26713_);
  or (_26717_, _26716_, _26438_);
  nand (_26719_, _26717_, _05846_);
  and (_26720_, _08701_, _07142_);
  nor (_26721_, _26720_, _06301_);
  nand (_26722_, _26721_, _26719_);
  and (_26723_, _26482_, _12682_);
  nor (_26724_, _12013_, _12682_);
  or (_26725_, _26724_, _06421_);
  nor (_26726_, _26725_, _26723_);
  nor (_26727_, _26726_, _12565_);
  and (_26728_, _26727_, _26722_);
  or (_26730_, _26728_, _26437_);
  nand (_26731_, _26730_, _12690_);
  nor (_26732_, _12690_, _12188_);
  nor (_26733_, _26732_, _10262_);
  nand (_26734_, _26733_, _26731_);
  and (_26735_, _26436_, _10262_);
  nor (_26736_, _26735_, _06167_);
  and (_26737_, _26736_, _26734_);
  and (_26738_, _08931_, _06167_);
  or (_26739_, _26738_, _26737_);
  nand (_26741_, _26739_, _12703_);
  and (_26742_, _08701_, _05826_);
  nor (_26743_, _26742_, _06165_);
  nand (_26744_, _26743_, _26741_);
  nor (_26745_, _26529_, _12682_);
  and (_26746_, _12014_, _12682_);
  nor (_26747_, _26746_, _26745_);
  and (_26748_, _26747_, _06165_);
  nor (_26749_, _26748_, _12712_);
  nand (_26750_, _26749_, _26744_);
  nor (_26751_, _26436_, _12711_);
  nor (_26752_, _26751_, _06433_);
  and (_26753_, _26752_, _26750_);
  or (_26754_, _26753_, _26432_);
  nand (_26755_, _26754_, _12719_);
  nor (_26756_, _26445_, _12719_);
  nor (_26757_, _26756_, _07577_);
  nand (_26758_, _26757_, _26755_);
  and (_26759_, _08701_, _07577_);
  nor (_26760_, _26759_, _05748_);
  nand (_26763_, _26760_, _26758_);
  and (_26764_, _26747_, _05748_);
  nor (_26765_, _26764_, _12737_);
  nand (_26766_, _26765_, _26763_);
  nor (_26767_, _26436_, _12735_);
  nor (_26768_, _26767_, _06440_);
  and (_26769_, _26768_, _26766_);
  or (_26770_, _26769_, _26431_);
  nand (_26771_, _26770_, _12744_);
  nor (_26772_, _26445_, _12744_);
  nor (_26774_, _26772_, _25019_);
  nand (_26775_, _26774_, _26771_);
  and (_26776_, _25019_, _08701_);
  nor (_26777_, _26776_, _12754_);
  and (_26778_, _26777_, _26775_);
  and (_26779_, _26436_, _12754_);
  or (_26780_, _26779_, _26778_);
  or (_26781_, _26780_, _01321_);
  or (_26782_, _01317_, \oc8051_golden_model_1.PC [5]);
  and (_26783_, _26782_, _43100_);
  and (_43693_, _26783_, _26781_);
  and (_26785_, _08432_, _05426_);
  nor (_26786_, _26785_, \oc8051_golden_model_1.PC [6]);
  nor (_26787_, _26786_, _11894_);
  and (_26788_, _26787_, _12754_);
  and (_26789_, _08638_, _07577_);
  not (_26790_, _26787_);
  and (_26791_, _26790_, _10262_);
  and (_26792_, _12181_, _06209_);
  or (_26793_, _26792_, _05829_);
  nor (_26795_, _25151_, _12180_);
  and (_26796_, _12050_, _12010_);
  nor (_26797_, _26796_, _12051_);
  or (_26798_, _26797_, _12141_);
  or (_26799_, _12139_, _12005_);
  and (_26800_, _26799_, _06160_);
  nand (_26801_, _26800_, _26798_);
  or (_26802_, _12256_, _12181_);
  and (_26803_, _12218_, _12185_);
  nor (_26804_, _26803_, _12219_);
  nand (_26806_, _26804_, _12256_);
  and (_26807_, _26806_, _08445_);
  nand (_26808_, _26807_, _26802_);
  and (_26809_, _08638_, _06581_);
  and (_26810_, _12181_, _07056_);
  or (_26811_, _26810_, _06653_);
  nand (_26812_, _12265_, \oc8051_golden_model_1.PC [6]);
  and (_26813_, _26812_, _07057_);
  or (_26814_, _26813_, _26811_);
  or (_26815_, _26790_, _12266_);
  and (_26817_, _26815_, _06582_);
  and (_26818_, _26817_, _26814_);
  or (_26819_, _26818_, _25055_);
  or (_26820_, _26819_, _26809_);
  or (_26821_, _26790_, _12263_);
  and (_26822_, _26821_, _08443_);
  nand (_26823_, _26822_, _26820_);
  and (_26824_, _26823_, _12281_);
  nand (_26825_, _26824_, _26808_);
  nand (_26826_, _26825_, _26801_);
  and (_26828_, _26826_, _12134_);
  and (_26829_, _26787_, _12287_);
  or (_26830_, _26829_, _06156_);
  or (_26831_, _26830_, _26828_);
  and (_26832_, _12181_, _06156_);
  nor (_26833_, _26832_, _07485_);
  nand (_26834_, _26833_, _26831_);
  nor (_26835_, _08638_, _05764_);
  nor (_26836_, _26835_, _06217_);
  nand (_26837_, _26836_, _26834_);
  and (_26839_, _12181_, _06217_);
  nor (_26840_, _26839_, _12293_);
  nand (_26841_, _26840_, _26837_);
  nor (_26842_, _26790_, _12292_);
  nor (_26843_, _26842_, _06220_);
  nand (_26844_, _26843_, _26841_);
  and (_26845_, _12181_, _06220_);
  nor (_26846_, _26845_, _12302_);
  nand (_26847_, _26846_, _26844_);
  nor (_26848_, _26790_, _12300_);
  nor (_26850_, _26848_, _06152_);
  and (_26851_, _26850_, _26847_);
  and (_26852_, _12181_, _06152_);
  or (_26853_, _26852_, _26851_);
  nand (_26854_, _26853_, _05769_);
  and (_26855_, _08638_, _12304_);
  nor (_26856_, _26855_, _06151_);
  nand (_26857_, _26856_, _26854_);
  and (_26858_, _12180_, _06151_);
  nor (_26859_, _26858_, _12126_);
  nand (_26861_, _26859_, _26857_);
  not (_26862_, _25114_);
  and (_26863_, _12120_, _12005_);
  not (_26864_, _26797_);
  nor (_26865_, _26864_, _12120_);
  or (_26866_, _26865_, _26863_);
  nor (_26867_, _26866_, _12125_);
  nor (_26868_, _26867_, _26862_);
  nand (_26869_, _26868_, _26861_);
  nor (_26870_, _26864_, _12329_);
  and (_26872_, _12329_, _12005_);
  nor (_26873_, _26872_, _26870_);
  nor (_26874_, _26873_, _06643_);
  or (_26875_, _12005_, _11956_);
  or (_26876_, _26797_, _11958_);
  and (_26877_, _26876_, _06687_);
  and (_26878_, _26877_, _26875_);
  nor (_26879_, _26878_, _26874_);
  nand (_26880_, _26879_, _26869_);
  nand (_26881_, _26880_, _12317_);
  nand (_26883_, _12346_, _12005_);
  nand (_26884_, _26797_, _12347_);
  and (_26885_, _26884_, _26883_);
  or (_26886_, _26885_, _12317_);
  and (_26887_, _26886_, _26881_);
  or (_26888_, _26887_, _11924_);
  nand (_26889_, _26787_, _11924_);
  and (_26890_, _26889_, _26888_);
  nand (_26891_, _26890_, _06146_);
  and (_26892_, _12181_, _06145_);
  nor (_26894_, _26892_, _07388_);
  nand (_26895_, _26894_, _26891_);
  nor (_26896_, _08638_, _05760_);
  nor (_26897_, _26896_, _25152_);
  and (_26898_, _26897_, _26895_);
  or (_26899_, _26898_, _26795_);
  nand (_26900_, _26899_, _12369_);
  nor (_26901_, _26787_, _12369_);
  nor (_26902_, _26901_, _06255_);
  nand (_26903_, _26902_, _26900_);
  and (_26905_, _12180_, _06255_);
  nor (_26906_, _26905_, _24882_);
  nand (_26907_, _26906_, _26903_);
  and (_26908_, _08638_, _24882_);
  nor (_26909_, _26908_, _06254_);
  nand (_26910_, _26909_, _26907_);
  and (_26911_, _12180_, _06254_);
  nor (_26912_, _26911_, _12387_);
  nand (_26913_, _26912_, _26910_);
  nor (_26914_, _26787_, _12381_);
  nor (_26916_, _26914_, _12386_);
  nand (_26917_, _26916_, _26913_);
  nor (_26918_, _12181_, _12385_);
  nor (_26919_, _26918_, _05870_);
  and (_26920_, _26919_, _26917_);
  nor (_26921_, _26787_, _05805_);
  or (_26922_, _26921_, _26920_);
  nand (_26923_, _26922_, _06140_);
  and (_26924_, _12181_, _06139_);
  nor (_26925_, _26924_, _05791_);
  nand (_26927_, _26925_, _26923_);
  nor (_26928_, _08638_, _24791_);
  nor (_26929_, _26928_, _06293_);
  and (_26930_, _26929_, _26927_);
  and (_26931_, _12006_, _06293_);
  or (_26932_, _26931_, _26930_);
  and (_26933_, _26932_, _06133_);
  nor (_26934_, _12180_, _06133_);
  or (_26935_, _26934_, _26933_);
  nand (_26936_, _26935_, _06114_);
  and (_26938_, _12006_, _05787_);
  nor (_26939_, _26938_, _12412_);
  nand (_26940_, _26939_, _26936_);
  nor (_26941_, _26790_, _11922_);
  nor (_26942_, _26941_, _06209_);
  and (_26943_, _26942_, _26940_);
  or (_26944_, _26943_, _26793_);
  nor (_26945_, _08638_, _05830_);
  nor (_26946_, _26945_, _12416_);
  and (_26947_, _26946_, _26944_);
  nor (_26949_, _26804_, _12417_);
  nor (_26950_, _26949_, _26947_);
  nand (_26951_, _26950_, _08787_);
  nor (_26952_, _12181_, _08787_);
  nor (_26953_, _26952_, _06110_);
  nand (_26954_, _26953_, _26951_);
  and (_26955_, _12006_, _06110_);
  nor (_26956_, _26955_, _10751_);
  nand (_26957_, _26956_, _26954_);
  and (_26958_, _12180_, _10751_);
  nor (_26960_, _26958_, _12431_);
  nand (_26961_, _26960_, _26957_);
  and (_26962_, _12453_, _12440_);
  nor (_26963_, _26962_, _12454_);
  nor (_26964_, _26963_, _12432_);
  nor (_26965_, _26964_, _06208_);
  nand (_26966_, _26965_, _26961_);
  and (_26967_, _12180_, _06208_);
  nor (_26968_, _26967_, _06076_);
  nand (_26969_, _26968_, _26966_);
  and (_26971_, _08638_, _06076_);
  nor (_26972_, _26971_, _12473_);
  nand (_26973_, _26972_, _26969_);
  and (_26974_, _12180_, _11101_);
  and (_26975_, _26804_, _12480_);
  or (_26976_, _26975_, _26974_);
  and (_26977_, _26976_, _12473_);
  nor (_26978_, _26977_, _12478_);
  nand (_26979_, _26978_, _26973_);
  nor (_26980_, _26787_, _11919_);
  nor (_26982_, _26980_, _11917_);
  nand (_26983_, _26982_, _26979_);
  nor (_26984_, _12181_, _11916_);
  nor (_26985_, _26984_, _06297_);
  and (_26986_, _26985_, _26983_);
  and (_26987_, _12006_, _06297_);
  or (_26988_, _26987_, _26986_);
  nand (_26989_, _26988_, _07125_);
  and (_26990_, _12181_, _06402_);
  nor (_26991_, _26990_, _12492_);
  and (_26993_, _26991_, _26989_);
  nor (_26994_, _08638_, _05834_);
  or (_26995_, _26994_, _26993_);
  nand (_26996_, _26995_, _12497_);
  nor (_26997_, _12181_, _11101_);
  and (_26998_, _26804_, _11101_);
  or (_26999_, _26998_, _26997_);
  and (_27000_, _26999_, _12496_);
  nor (_27001_, _27000_, _12505_);
  nand (_27002_, _27001_, _26996_);
  nor (_27004_, _26787_, _11914_);
  nor (_27005_, _27004_, _10822_);
  nand (_27006_, _27005_, _27002_);
  nor (_27007_, _12181_, _10821_);
  nor (_27008_, _27007_, _06306_);
  and (_27009_, _27008_, _27006_);
  and (_27010_, _12006_, _06306_);
  or (_27011_, _27010_, _27009_);
  nand (_27012_, _27011_, _07130_);
  and (_27013_, _12181_, _06411_);
  nor (_27015_, _27013_, _07124_);
  and (_27016_, _27015_, _27012_);
  nor (_27017_, _08638_, _05848_);
  or (_27018_, _27017_, _27016_);
  nand (_27019_, _27018_, _12518_);
  and (_27020_, _12180_, \oc8051_golden_model_1.PSW [7]);
  and (_27021_, _26804_, _10693_);
  or (_27022_, _27021_, _27020_);
  and (_27023_, _27022_, _12517_);
  nor (_27024_, _27023_, _12522_);
  nand (_27026_, _27024_, _27019_);
  nor (_27027_, _26787_, _11912_);
  nor (_27028_, _27027_, _10850_);
  nand (_27029_, _27028_, _27026_);
  nor (_27030_, _12181_, _10849_);
  nor (_27031_, _27030_, _06303_);
  and (_27032_, _27031_, _27029_);
  and (_27033_, _12006_, _06303_);
  or (_27034_, _27033_, _27032_);
  nand (_27035_, _27034_, _08824_);
  and (_27037_, _12181_, _06396_);
  nor (_27038_, _27037_, _05842_);
  and (_27039_, _27038_, _27035_);
  nor (_27040_, _08638_, _05843_);
  or (_27041_, _27040_, _27039_);
  nand (_27042_, _27041_, _12539_);
  or (_27043_, _26804_, _10693_);
  or (_27044_, _12180_, \oc8051_golden_model_1.PSW [7]);
  and (_27045_, _27044_, _12538_);
  and (_27046_, _27045_, _27043_);
  nor (_27048_, _27046_, _12547_);
  nand (_27049_, _27048_, _27042_);
  nor (_27050_, _26787_, _11907_);
  nor (_27051_, _27050_, _10897_);
  nand (_27052_, _27051_, _27049_);
  nor (_27053_, _12181_, _10896_);
  nor (_27054_, _27053_, _10925_);
  nand (_27055_, _27054_, _27052_);
  and (_27056_, _26790_, _10925_);
  nor (_27057_, _27056_, _06417_);
  nand (_27059_, _27057_, _27055_);
  and (_27060_, _09207_, _06417_);
  nor (_27061_, _27060_, _07142_);
  nand (_27062_, _27061_, _27059_);
  and (_27063_, _08638_, _07142_);
  nor (_27064_, _27063_, _06301_);
  nand (_27065_, _27064_, _27062_);
  and (_27066_, _26864_, _12682_);
  nor (_27067_, _12005_, _12682_);
  or (_27068_, _27067_, _06421_);
  nor (_27070_, _27068_, _27066_);
  nor (_27071_, _27070_, _12565_);
  nand (_27072_, _27071_, _27065_);
  nor (_27073_, _26787_, _11905_);
  nor (_27074_, _27073_, _12691_);
  nand (_27075_, _27074_, _27072_);
  nor (_27076_, _12690_, _12181_);
  nor (_27077_, _27076_, _10262_);
  and (_27078_, _27077_, _27075_);
  or (_27079_, _27078_, _26791_);
  nand (_27081_, _27079_, _06168_);
  and (_27082_, _08883_, _06167_);
  nor (_27083_, _27082_, _05826_);
  nand (_27084_, _27083_, _27081_);
  nor (_27085_, _08638_, _12703_);
  nor (_27086_, _27085_, _06165_);
  and (_27087_, _27086_, _27084_);
  and (_27088_, _12006_, _12682_);
  nor (_27089_, _26797_, _12682_);
  nor (_27090_, _27089_, _27088_);
  nor (_27092_, _27090_, _06166_);
  or (_27093_, _27092_, _27087_);
  and (_27094_, _27093_, _12711_);
  nor (_27095_, _26787_, _12711_);
  or (_27096_, _27095_, _27094_);
  nand (_27097_, _27096_, _06829_);
  and (_27098_, _12181_, _06433_);
  nor (_27099_, _27098_, _25721_);
  nand (_27100_, _27099_, _27097_);
  nor (_27101_, _26790_, _12719_);
  nor (_27103_, _27101_, _07577_);
  and (_27104_, _27103_, _27100_);
  or (_27105_, _27104_, _26789_);
  nand (_27106_, _27105_, _05749_);
  nor (_27107_, _27090_, _05749_);
  nor (_27108_, _27107_, _12737_);
  nand (_27109_, _27108_, _27106_);
  nor (_27110_, _26790_, _12735_);
  nor (_27111_, _27110_, _06440_);
  nand (_27112_, _27111_, _27109_);
  and (_27114_, _12181_, _06440_);
  nor (_27115_, _27114_, _26415_);
  nand (_27116_, _27115_, _27112_);
  nor (_27117_, _26790_, _12744_);
  nor (_27118_, _27117_, _25019_);
  nand (_27119_, _27118_, _27116_);
  and (_27120_, _25019_, _08638_);
  nor (_27121_, _27120_, _12754_);
  and (_27122_, _27121_, _27119_);
  or (_27123_, _27122_, _26788_);
  or (_27125_, _27123_, _01321_);
  or (_27126_, _01317_, \oc8051_golden_model_1.PC [6]);
  and (_27127_, _27126_, _43100_);
  and (_43694_, _27127_, _27125_);
  and (_27128_, _08437_, _06440_);
  nor (_27129_, _11894_, \oc8051_golden_model_1.PC [7]);
  nor (_27130_, _27129_, _11895_);
  nor (_27131_, _27130_, _11905_);
  nor (_27132_, _27130_, _11907_);
  nor (_27133_, _27130_, _11912_);
  nor (_27135_, _27130_, _11914_);
  nor (_27136_, _27130_, _11919_);
  nor (_27137_, _08787_, _08437_);
  nor (_27138_, _25151_, _08437_);
  not (_27139_, _27130_);
  nand (_27140_, _27139_, _11924_);
  and (_27141_, _12141_, _09180_);
  or (_27142_, _12001_, _12002_);
  and (_27143_, _27142_, _12052_);
  nor (_27144_, _27142_, _12052_);
  nor (_27146_, _27144_, _27143_);
  and (_27147_, _27146_, _12139_);
  or (_27148_, _27147_, _27141_);
  and (_27149_, _27148_, _06160_);
  or (_27150_, _12176_, _12177_);
  and (_27151_, _27150_, _12220_);
  nor (_27152_, _27150_, _12220_);
  nor (_27153_, _27152_, _27151_);
  and (_27154_, _27153_, _12256_);
  and (_27155_, _12258_, _08437_);
  or (_27157_, _27155_, _27154_);
  and (_27158_, _27157_, _08445_);
  nor (_27159_, _08395_, _06582_);
  nand (_27160_, _08573_, _07056_);
  and (_27161_, _27160_, _12264_);
  and (_27162_, _12265_, \oc8051_golden_model_1.PC [7]);
  or (_27163_, _27162_, _07056_);
  and (_27164_, _27163_, _27161_);
  or (_27165_, _27139_, _12266_);
  nand (_27166_, _27165_, _12263_);
  or (_27168_, _27166_, _27164_);
  and (_27169_, _27168_, _06582_);
  or (_27170_, _27169_, _27159_);
  or (_27171_, _27130_, _12263_);
  and (_27172_, _27171_, _08443_);
  and (_27173_, _27172_, _27170_);
  or (_27174_, _27173_, _07064_);
  or (_27175_, _27174_, _27158_);
  nand (_27176_, _27139_, _07064_);
  and (_27177_, _27176_, _06161_);
  and (_27179_, _27177_, _27175_);
  or (_27180_, _27179_, _27149_);
  or (_27181_, _27180_, _24821_);
  or (_27182_, _27130_, _12134_);
  and (_27183_, _27182_, _06157_);
  and (_27184_, _27183_, _27181_);
  and (_27185_, _08437_, _06156_);
  or (_27186_, _27185_, _07485_);
  or (_27187_, _27186_, _27184_);
  nand (_27188_, _08395_, _07485_);
  and (_27190_, _27188_, _07075_);
  and (_27191_, _27190_, _27187_);
  nand (_27192_, _08437_, _06217_);
  nand (_27193_, _27192_, _12292_);
  or (_27194_, _27193_, _27191_);
  or (_27195_, _27130_, _12292_);
  and (_27196_, _27195_, _06229_);
  and (_27197_, _27196_, _27194_);
  nand (_27198_, _08437_, _06220_);
  nand (_27199_, _27198_, _12300_);
  or (_27201_, _27199_, _27197_);
  or (_27202_, _27130_, _12300_);
  and (_27203_, _27202_, _06153_);
  and (_27204_, _27203_, _27201_);
  and (_27205_, _08437_, _06152_);
  or (_27206_, _27205_, _12304_);
  or (_27207_, _27206_, _27204_);
  nand (_27208_, _08395_, _12304_);
  and (_27209_, _27208_, _07191_);
  and (_27210_, _27209_, _27207_);
  nand (_27212_, _08437_, _06151_);
  nand (_27213_, _27212_, _12125_);
  or (_27214_, _27213_, _27210_);
  not (_27215_, _27146_);
  nor (_27216_, _27215_, _12120_);
  and (_27217_, _12120_, _09180_);
  or (_27218_, _27217_, _12125_);
  or (_27219_, _27218_, _27216_);
  and (_27220_, _27219_, _12089_);
  and (_27221_, _27220_, _27214_);
  and (_27223_, _27146_, _11956_);
  and (_27224_, _11958_, _09180_);
  or (_27225_, _27224_, _27223_);
  and (_27226_, _27225_, _06687_);
  or (_27227_, _27226_, _06236_);
  or (_27228_, _27227_, _27221_);
  and (_27229_, _12329_, _09180_);
  nor (_27230_, _27215_, _12329_);
  or (_27231_, _27230_, _06643_);
  or (_27232_, _27231_, _27229_);
  and (_27234_, _27232_, _12317_);
  and (_27235_, _27234_, _27228_);
  or (_27236_, _27146_, _12346_);
  nand (_27237_, _12346_, _09181_);
  and (_27238_, _27237_, _06295_);
  and (_27239_, _27238_, _27236_);
  or (_27240_, _27239_, _11924_);
  or (_27241_, _27240_, _27235_);
  nand (_27242_, _27241_, _27140_);
  nand (_27243_, _27242_, _06146_);
  and (_27245_, _08573_, _06145_);
  nor (_27246_, _27245_, _07388_);
  nand (_27247_, _27246_, _27243_);
  nor (_27248_, _08395_, _05760_);
  nor (_27249_, _27248_, _25152_);
  and (_27250_, _27249_, _27247_);
  or (_27251_, _27250_, _27138_);
  nand (_27252_, _27251_, _12369_);
  nor (_27253_, _27130_, _12369_);
  nor (_27254_, _27253_, _06255_);
  nand (_27256_, _27254_, _27252_);
  and (_27257_, _08437_, _06255_);
  nor (_27258_, _27257_, _24882_);
  nand (_27259_, _27258_, _27256_);
  and (_27260_, _08395_, _24882_);
  nor (_27261_, _27260_, _06254_);
  nand (_27262_, _27261_, _27259_);
  and (_27263_, _08437_, _06254_);
  nor (_27264_, _27263_, _12387_);
  and (_27265_, _27264_, _27262_);
  nor (_27267_, _27130_, _12381_);
  or (_27268_, _27267_, _27265_);
  nand (_27269_, _27268_, _12385_);
  nor (_27270_, _12385_, _08437_);
  nor (_27271_, _27270_, _05870_);
  nand (_27272_, _27271_, _27269_);
  nor (_27273_, _27139_, _05805_);
  nor (_27274_, _27273_, _06139_);
  and (_27275_, _27274_, _27272_);
  and (_27276_, _08573_, _06139_);
  or (_27278_, _27276_, _27275_);
  nand (_27279_, _27278_, _24791_);
  and (_27280_, _08395_, _05791_);
  nor (_27281_, _27280_, _06293_);
  nand (_27282_, _27281_, _27279_);
  and (_27283_, _09180_, _06293_);
  nor (_27284_, _27283_, _13620_);
  nand (_27285_, _27284_, _27282_);
  nor (_27286_, _08437_, _06133_);
  nor (_27287_, _27286_, _05787_);
  nand (_27289_, _27287_, _27285_);
  and (_27290_, _09180_, _05787_);
  nor (_27291_, _27290_, _12412_);
  nand (_27292_, _27291_, _27289_);
  nor (_27293_, _27130_, _11922_);
  nor (_27294_, _27293_, _06209_);
  nand (_27295_, _27294_, _27292_);
  and (_27296_, _08437_, _06209_);
  nor (_27297_, _27296_, _05829_);
  nand (_27298_, _27297_, _27295_);
  and (_27300_, _08395_, _05829_);
  nor (_27301_, _27300_, _12416_);
  nand (_27302_, _27301_, _27298_);
  and (_27303_, _27153_, _12416_);
  nor (_27304_, _27303_, _08788_);
  and (_27305_, _27304_, _27302_);
  or (_27306_, _27305_, _27137_);
  nand (_27307_, _27306_, _06111_);
  and (_27308_, _09181_, _06110_);
  nor (_27309_, _27308_, _10751_);
  and (_27311_, _27309_, _27307_);
  and (_27312_, _10751_, _08437_);
  or (_27313_, _27312_, _27311_);
  nand (_27314_, _27313_, _12432_);
  or (_27315_, _12436_, _12435_);
  nor (_27316_, _27315_, _12455_);
  not (_27317_, _27316_);
  and (_27318_, _27315_, _12455_);
  nor (_27319_, _27318_, _12432_);
  and (_27320_, _27319_, _27317_);
  nor (_27322_, _27320_, _06208_);
  and (_27323_, _27322_, _27314_);
  and (_27324_, _08573_, _06208_);
  or (_27325_, _27324_, _27323_);
  nand (_27326_, _27325_, _05836_);
  and (_27327_, _08395_, _06076_);
  nor (_27328_, _27327_, _12473_);
  nand (_27329_, _27328_, _27326_);
  and (_27330_, _11101_, _08437_);
  and (_27331_, _27153_, _12480_);
  or (_27332_, _27331_, _27330_);
  and (_27333_, _27332_, _12473_);
  nor (_27334_, _27333_, _12478_);
  and (_27335_, _27334_, _27329_);
  or (_27336_, _27335_, _27136_);
  nand (_27337_, _27336_, _11916_);
  nor (_27338_, _11916_, _08437_);
  nor (_27339_, _27338_, _06297_);
  nand (_27340_, _27339_, _27337_);
  and (_27341_, _09180_, _06297_);
  nor (_27344_, _27341_, _06402_);
  and (_27345_, _27344_, _27340_);
  and (_27346_, _08573_, _06402_);
  or (_27347_, _27346_, _27345_);
  nand (_27348_, _27347_, _05834_);
  and (_27349_, _08395_, _12492_);
  nor (_27350_, _27349_, _12496_);
  nand (_27351_, _27350_, _27348_);
  nor (_27352_, _27153_, _12480_);
  nor (_27353_, _11101_, _08437_);
  nor (_27355_, _27353_, _12497_);
  not (_27356_, _27355_);
  nor (_27357_, _27356_, _27352_);
  nor (_27358_, _27357_, _12505_);
  and (_27359_, _27358_, _27351_);
  or (_27360_, _27359_, _27135_);
  nand (_27361_, _27360_, _10821_);
  nor (_27362_, _10821_, _08437_);
  nor (_27363_, _27362_, _06306_);
  nand (_27364_, _27363_, _27361_);
  and (_27366_, _09180_, _06306_);
  nor (_27367_, _27366_, _06411_);
  and (_27368_, _27367_, _27364_);
  and (_27369_, _08573_, _06411_);
  or (_27370_, _27369_, _27368_);
  nand (_27371_, _27370_, _05848_);
  and (_27372_, _08395_, _07124_);
  nor (_27373_, _27372_, _12517_);
  nand (_27374_, _27373_, _27371_);
  and (_27375_, _08437_, \oc8051_golden_model_1.PSW [7]);
  and (_27377_, _27153_, _10693_);
  or (_27378_, _27377_, _27375_);
  and (_27379_, _27378_, _12517_);
  nor (_27380_, _27379_, _12522_);
  and (_27381_, _27380_, _27374_);
  or (_27382_, _27381_, _27133_);
  nand (_27383_, _27382_, _10849_);
  nor (_27384_, _10849_, _08437_);
  nor (_27385_, _27384_, _06303_);
  nand (_27386_, _27385_, _27383_);
  and (_27388_, _09180_, _06303_);
  nor (_27389_, _27388_, _06396_);
  and (_27390_, _27389_, _27386_);
  and (_27391_, _08573_, _06396_);
  or (_27392_, _27391_, _27390_);
  nand (_27393_, _27392_, _05843_);
  and (_27394_, _08395_, _05842_);
  nor (_27395_, _27394_, _12538_);
  nand (_27396_, _27395_, _27393_);
  and (_27397_, _08437_, _10693_);
  and (_27399_, _27153_, \oc8051_golden_model_1.PSW [7]);
  or (_27400_, _27399_, _27397_);
  and (_27401_, _27400_, _12538_);
  nor (_27402_, _27401_, _12547_);
  and (_27403_, _27402_, _27396_);
  or (_27404_, _27403_, _27132_);
  nand (_27405_, _27404_, _10896_);
  nor (_27406_, _10896_, _08437_);
  nor (_27407_, _27406_, _10925_);
  nand (_27408_, _27407_, _27405_);
  and (_27410_, _27130_, _10925_);
  nor (_27411_, _27410_, _06417_);
  and (_27412_, _27411_, _27408_);
  and (_27413_, _08838_, _06417_);
  or (_27414_, _27413_, _27412_);
  nand (_27415_, _27414_, _05846_);
  and (_27416_, _08395_, _07142_);
  nor (_27417_, _27416_, _06301_);
  nand (_27418_, _27417_, _27415_);
  and (_27419_, _27215_, _12682_);
  nor (_27421_, _09180_, _12682_);
  or (_27422_, _27421_, _06421_);
  nor (_27423_, _27422_, _27419_);
  nor (_27424_, _27423_, _12565_);
  and (_27425_, _27424_, _27418_);
  or (_27426_, _27425_, _27131_);
  nand (_27427_, _27426_, _12690_);
  nor (_27428_, _12690_, _08437_);
  nor (_27429_, _27428_, _10262_);
  nand (_27430_, _27429_, _27427_);
  and (_27432_, _27130_, _10262_);
  nor (_27433_, _27432_, _06167_);
  and (_27434_, _27433_, _27430_);
  and (_27435_, _08838_, _06167_);
  or (_27436_, _27435_, _27434_);
  nand (_27437_, _27436_, _12703_);
  and (_27438_, _08395_, _05826_);
  nor (_27439_, _27438_, _06165_);
  nand (_27440_, _27439_, _27437_);
  nor (_27441_, _27146_, _12682_);
  and (_27443_, _09181_, _12682_);
  nor (_27444_, _27443_, _27441_);
  and (_27445_, _27444_, _06165_);
  nor (_27446_, _27445_, _12712_);
  nand (_27447_, _27446_, _27440_);
  nor (_27448_, _27130_, _12711_);
  nor (_27449_, _27448_, _06433_);
  nand (_27450_, _27449_, _27447_);
  and (_27451_, _08437_, _06433_);
  nor (_27452_, _27451_, _25721_);
  and (_27454_, _27452_, _27450_);
  nor (_27455_, _27130_, _12719_);
  or (_27456_, _27455_, _27454_);
  nand (_27457_, _27456_, _07160_);
  and (_27458_, _08395_, _07577_);
  nor (_27459_, _27458_, _05748_);
  nand (_27460_, _27459_, _27457_);
  and (_27461_, _27444_, _05748_);
  nor (_27462_, _27461_, _12737_);
  nand (_27463_, _27462_, _27460_);
  nor (_27465_, _27130_, _12735_);
  nor (_27466_, _27465_, _06440_);
  and (_27467_, _27466_, _27463_);
  or (_27468_, _27467_, _27128_);
  nand (_27469_, _27468_, _12744_);
  nor (_27470_, _27139_, _12744_);
  nor (_27471_, _27470_, _25019_);
  nand (_27472_, _27471_, _27469_);
  and (_27473_, _25019_, _08395_);
  nor (_27474_, _27473_, _12754_);
  and (_27476_, _27474_, _27472_);
  and (_27477_, _27130_, _12754_);
  or (_27478_, _27477_, _27476_);
  or (_27479_, _27478_, _01321_);
  or (_27480_, _01317_, \oc8051_golden_model_1.PC [7]);
  and (_27481_, _27480_, _43100_);
  and (_43695_, _27481_, _27479_);
  nor (_27482_, _12747_, _06107_);
  nor (_27483_, _12723_, _06107_);
  nor (_27484_, _12538_, _05842_);
  nor (_27486_, _12416_, _05829_);
  and (_27487_, _12224_, _06209_);
  and (_27488_, _12224_, _06152_);
  nor (_27489_, _06217_, _07485_);
  and (_27490_, _12224_, _06156_);
  and (_27491_, _11895_, \oc8051_golden_model_1.PC [8]);
  nor (_27492_, _11895_, \oc8051_golden_model_1.PC [8]);
  nor (_27493_, _27492_, _27491_);
  nor (_27494_, _27493_, _12266_);
  not (_27495_, _12224_);
  and (_27497_, _27495_, _07056_);
  nor (_27498_, _07056_, \oc8051_golden_model_1.PC [8]);
  and (_27499_, _27498_, _12265_);
  or (_27500_, _27499_, _27497_);
  and (_27501_, _27500_, _12264_);
  nor (_27502_, _27501_, _27494_);
  nor (_27503_, _27502_, _24800_);
  nor (_27504_, _27493_, _12263_);
  nor (_27505_, _27504_, _27503_);
  nor (_27506_, _27505_, _08445_);
  or (_27508_, _12256_, _27495_);
  nor (_27509_, _12227_, _12222_);
  nor (_27510_, _27509_, _12228_);
  nand (_27511_, _27510_, _12256_);
  and (_27512_, _27511_, _08445_);
  and (_27513_, _27512_, _27508_);
  or (_27514_, _27513_, _27506_);
  nand (_27515_, _27514_, _07065_);
  not (_27516_, _27493_);
  and (_27517_, _27516_, _07064_);
  nor (_27519_, _27517_, _06160_);
  nand (_27520_, _27519_, _27515_);
  or (_27521_, _12139_, _12056_);
  nor (_27522_, _12060_, _12054_);
  nor (_27523_, _27522_, _12061_);
  or (_27524_, _27523_, _12141_);
  and (_27525_, _27524_, _06160_);
  nand (_27526_, _27525_, _27521_);
  and (_27527_, _27526_, _12134_);
  nand (_27528_, _27527_, _27520_);
  nor (_27530_, _27493_, _12134_);
  nor (_27531_, _27530_, _06156_);
  and (_27532_, _27531_, _27528_);
  or (_27533_, _27532_, _27490_);
  nand (_27534_, _27533_, _27489_);
  and (_27535_, _12224_, _06217_);
  nor (_27536_, _27535_, _12293_);
  nand (_27537_, _27536_, _27534_);
  nor (_27538_, _27493_, _12292_);
  nor (_27539_, _27538_, _06220_);
  nand (_27541_, _27539_, _27537_);
  and (_27542_, _12224_, _06220_);
  nor (_27543_, _27542_, _12302_);
  nand (_27544_, _27543_, _27541_);
  nor (_27545_, _27493_, _12300_);
  nor (_27546_, _27545_, _06152_);
  and (_27547_, _27546_, _27544_);
  or (_27548_, _27547_, _27488_);
  nand (_27549_, _27548_, _12305_);
  and (_27550_, _12224_, _06151_);
  nor (_27552_, _27550_, _12126_);
  nand (_27553_, _27552_, _27549_);
  and (_27554_, _12120_, _12056_);
  not (_27555_, _27523_);
  nor (_27556_, _27555_, _12120_);
  or (_27557_, _27556_, _27554_);
  nor (_27558_, _27557_, _12125_);
  nor (_27559_, _27558_, _26862_);
  nand (_27560_, _27559_, _27553_);
  nor (_27561_, _27555_, _12329_);
  and (_27563_, _12329_, _12056_);
  nor (_27564_, _27563_, _27561_);
  nor (_27565_, _27564_, _06643_);
  or (_27566_, _12056_, _11956_);
  nand (_27567_, _27555_, _11956_);
  and (_27568_, _27567_, _06687_);
  and (_27569_, _27568_, _27566_);
  nor (_27570_, _27569_, _27565_);
  nand (_27571_, _27570_, _27560_);
  nand (_27572_, _27571_, _12317_);
  nor (_27574_, _27523_, _12346_);
  and (_27575_, _12346_, _12057_);
  nor (_27576_, _27575_, _12317_);
  not (_27577_, _27576_);
  nor (_27578_, _27577_, _27574_);
  nor (_27579_, _27578_, _11924_);
  nand (_27580_, _27579_, _27572_);
  and (_27581_, _27516_, _11924_);
  nor (_27582_, _27581_, _06145_);
  nand (_27583_, _27582_, _27580_);
  and (_27585_, _12224_, _06145_);
  nor (_27586_, _27585_, _07388_);
  nand (_27587_, _27586_, _27583_);
  nand (_27588_, _27587_, _25151_);
  nor (_27589_, _25151_, _27495_);
  nor (_27590_, _27589_, _12373_);
  nand (_27591_, _27590_, _27588_);
  nor (_27592_, _27493_, _12369_);
  nor (_27593_, _27592_, _06255_);
  nand (_27594_, _27593_, _27591_);
  and (_27596_, _12224_, _06255_);
  nor (_27597_, _27596_, _24882_);
  nand (_27598_, _27597_, _27594_);
  nand (_27599_, _27598_, _13843_);
  and (_27600_, _12224_, _06254_);
  nor (_27601_, _27600_, _12387_);
  nand (_27602_, _27601_, _27599_);
  nor (_27603_, _27493_, _12381_);
  nor (_27604_, _27603_, _12386_);
  and (_27605_, _27604_, _27602_);
  nor (_27607_, _27495_, _12385_);
  or (_27608_, _27607_, _05870_);
  nor (_27609_, _27608_, _27605_);
  nor (_27610_, _27493_, _05805_);
  or (_27611_, _27610_, _27609_);
  nand (_27612_, _27611_, _06140_);
  and (_27613_, _27495_, _06139_);
  nor (_27614_, _06293_, _05791_);
  not (_27615_, _27614_);
  nor (_27616_, _27615_, _27613_);
  nand (_27618_, _27616_, _27612_);
  and (_27619_, _12056_, _06293_);
  nor (_27620_, _27619_, _13620_);
  nand (_27621_, _27620_, _27618_);
  nor (_27622_, _12224_, _06133_);
  nor (_27623_, _27622_, _05787_);
  nand (_27624_, _27623_, _27621_);
  and (_27625_, _12056_, _05787_);
  nor (_27626_, _27625_, _12412_);
  nand (_27627_, _27626_, _27624_);
  nor (_27629_, _27493_, _11922_);
  nor (_27630_, _27629_, _06209_);
  and (_27631_, _27630_, _27627_);
  or (_27632_, _27631_, _27487_);
  nand (_27633_, _27632_, _27486_);
  and (_27634_, _27510_, _12416_);
  nor (_27635_, _27634_, _08788_);
  and (_27636_, _27635_, _27633_);
  nor (_27637_, _12224_, _08787_);
  or (_27638_, _27637_, _27636_);
  nand (_27640_, _27638_, _06111_);
  and (_27641_, _12057_, _06110_);
  nor (_27642_, _27641_, _10751_);
  nand (_27643_, _27642_, _27640_);
  and (_27644_, _12224_, _10751_);
  nor (_27645_, _27644_, _12431_);
  nand (_27646_, _27645_, _27643_);
  and (_27647_, _12457_, _12434_);
  nor (_27648_, _27647_, _12458_);
  nor (_27649_, _27648_, _12432_);
  nor (_27651_, _27649_, _06208_);
  nand (_27652_, _27651_, _27646_);
  and (_27653_, _12224_, _06208_);
  nor (_27654_, _27653_, _06076_);
  nand (_27655_, _27654_, _27652_);
  nand (_27656_, _27655_, _12474_);
  and (_27657_, _12224_, _11101_);
  and (_27658_, _27510_, _12480_);
  or (_27659_, _27658_, _27657_);
  and (_27660_, _27659_, _12473_);
  nor (_27662_, _27660_, _12478_);
  nand (_27663_, _27662_, _27656_);
  nor (_27664_, _27493_, _11919_);
  nor (_27665_, _27664_, _11917_);
  nand (_27666_, _27665_, _27663_);
  nor (_27667_, _27495_, _11916_);
  nor (_27668_, _27667_, _06297_);
  nand (_27669_, _27668_, _27666_);
  and (_27670_, _12057_, _06297_);
  nor (_27671_, _27670_, _06402_);
  nand (_27673_, _27671_, _27669_);
  and (_27674_, _12224_, _06402_);
  nor (_27675_, _27674_, _12492_);
  nand (_27676_, _27675_, _27673_);
  nand (_27677_, _27676_, _12497_);
  nor (_27678_, _27510_, _12480_);
  nor (_27679_, _12224_, _11101_);
  nor (_27680_, _27679_, _12497_);
  not (_27681_, _27680_);
  nor (_27682_, _27681_, _27678_);
  nor (_27684_, _27682_, _12505_);
  nand (_27685_, _27684_, _27677_);
  nor (_27686_, _27493_, _11914_);
  nor (_27687_, _27686_, _10822_);
  nand (_27688_, _27687_, _27685_);
  nor (_27689_, _27495_, _10821_);
  nor (_27690_, _27689_, _06306_);
  and (_27691_, _27690_, _27688_);
  and (_27692_, _12057_, _06306_);
  or (_27693_, _27692_, _27691_);
  nand (_27695_, _27693_, _07130_);
  nor (_27696_, _12517_, _07124_);
  and (_27697_, _27495_, _06411_);
  not (_27698_, _27697_);
  and (_27699_, _27698_, _27696_);
  nand (_27700_, _27699_, _27695_);
  and (_27701_, _12224_, \oc8051_golden_model_1.PSW [7]);
  and (_27702_, _27510_, _10693_);
  or (_27703_, _27702_, _27701_);
  and (_27704_, _27703_, _12517_);
  nor (_27706_, _27704_, _12522_);
  nand (_27707_, _27706_, _27700_);
  nor (_27708_, _27493_, _11912_);
  nor (_27709_, _27708_, _10850_);
  and (_27710_, _27709_, _27707_);
  nor (_27711_, _27495_, _10849_);
  or (_27712_, _27711_, _06303_);
  or (_27713_, _27712_, _27710_);
  and (_27714_, _12057_, _06303_);
  nor (_27715_, _27714_, _06396_);
  and (_27717_, _27715_, _27713_);
  and (_27718_, _12224_, _06396_);
  or (_27719_, _27718_, _27717_);
  nand (_27720_, _27719_, _27484_);
  and (_27721_, _12224_, _10693_);
  and (_27722_, _27510_, \oc8051_golden_model_1.PSW [7]);
  or (_27723_, _27722_, _27721_);
  and (_27724_, _27723_, _12538_);
  nor (_27725_, _27724_, _12547_);
  nand (_27726_, _27725_, _27720_);
  nor (_27728_, _27493_, _11907_);
  nor (_27729_, _27728_, _10897_);
  nand (_27730_, _27729_, _27726_);
  nor (_27731_, _27495_, _10896_);
  nor (_27732_, _27731_, _10925_);
  nand (_27733_, _27732_, _27730_);
  and (_27734_, _27516_, _10925_);
  nor (_27735_, _27734_, _06417_);
  nand (_27736_, _27735_, _27733_);
  and (_27737_, _07049_, _06417_);
  nor (_27739_, _27737_, _07142_);
  nand (_27740_, _27739_, _27736_);
  nand (_27741_, _27740_, _06421_);
  and (_27742_, _27555_, _12682_);
  nor (_27743_, _12056_, _12682_);
  or (_27744_, _27743_, _06421_);
  nor (_27745_, _27744_, _27742_);
  nor (_27746_, _27745_, _12565_);
  nand (_27747_, _27746_, _27741_);
  nor (_27748_, _27493_, _11905_);
  nor (_27750_, _27748_, _12691_);
  nand (_27751_, _27750_, _27747_);
  nor (_27752_, _12690_, _27495_);
  nor (_27753_, _27752_, _10262_);
  nand (_27754_, _27753_, _27751_);
  and (_27755_, _27516_, _10262_);
  nor (_27756_, _27755_, _06167_);
  nand (_27757_, _27756_, _27754_);
  and (_27758_, _07049_, _06167_);
  nor (_27759_, _27758_, _05826_);
  nand (_27761_, _27759_, _27757_);
  nand (_27762_, _27761_, _06166_);
  nor (_27763_, _27523_, _12682_);
  and (_27764_, _12057_, _12682_);
  nor (_27765_, _27764_, _27763_);
  and (_27766_, _27765_, _06165_);
  nor (_27767_, _27766_, _12712_);
  nand (_27768_, _27767_, _27762_);
  nor (_27769_, _27493_, _12711_);
  nor (_27770_, _27769_, _06433_);
  nand (_27772_, _27770_, _27768_);
  and (_27773_, _12224_, _06433_);
  nor (_27774_, _27773_, _25721_);
  nand (_27775_, _27774_, _27772_);
  nor (_27776_, _27493_, _12719_);
  nor (_27777_, _27776_, _06310_);
  and (_27778_, _27777_, _27775_);
  or (_27779_, _27778_, _27483_);
  nor (_27780_, _05823_, _05748_);
  nand (_27781_, _27780_, _27779_);
  and (_27783_, _27765_, _05748_);
  nor (_27784_, _27783_, _12737_);
  nand (_27785_, _27784_, _27781_);
  nor (_27786_, _27493_, _12735_);
  nor (_27787_, _27786_, _06440_);
  nand (_27788_, _27787_, _27785_);
  and (_27789_, _12224_, _06440_);
  nor (_27790_, _27789_, _26415_);
  nand (_27791_, _27790_, _27788_);
  nor (_27792_, _27493_, _12744_);
  nor (_27794_, _27792_, _06305_);
  and (_27795_, _27794_, _27791_);
  or (_27796_, _27795_, _27482_);
  nor (_27797_, _12754_, _05821_);
  and (_27798_, _27797_, _27796_);
  and (_27799_, _27493_, _12754_);
  or (_27800_, _27799_, _27798_);
  or (_27801_, _27800_, _01321_);
  or (_27802_, _01317_, \oc8051_golden_model_1.PC [8]);
  and (_27803_, _27802_, _43100_);
  and (_43696_, _27803_, _27801_);
  nor (_27805_, _06912_, _12747_);
  nor (_27806_, _06912_, _12723_);
  nor (_27807_, _27491_, \oc8051_golden_model_1.PC [9]);
  nor (_27808_, _27807_, _11896_);
  nor (_27809_, _27808_, _11905_);
  nor (_27810_, _27808_, _11907_);
  and (_27811_, _11996_, _06303_);
  nor (_27812_, _27808_, _11912_);
  and (_27813_, _11996_, _06306_);
  nor (_27815_, _27808_, _11914_);
  and (_27816_, _11996_, _06297_);
  nor (_27817_, _27808_, _11919_);
  nor (_27818_, _12172_, _08787_);
  and (_27819_, _12172_, _06209_);
  and (_27820_, _12172_, _06254_);
  nor (_27821_, _06254_, _24882_);
  and (_27822_, _12172_, _06255_);
  or (_27823_, _12139_, _11996_);
  nor (_27824_, _12061_, _12058_);
  and (_27826_, _27824_, _12000_);
  nor (_27827_, _27824_, _12000_);
  nor (_27828_, _27827_, _27826_);
  not (_27829_, _27828_);
  or (_27830_, _27829_, _12141_);
  and (_27831_, _27830_, _27823_);
  or (_27832_, _27831_, _06161_);
  nor (_27833_, _12228_, _12225_);
  and (_27834_, _27833_, _12175_);
  nor (_27835_, _27833_, _12175_);
  nor (_27837_, _27835_, _27834_);
  or (_27838_, _27837_, _12258_);
  not (_27839_, _12172_);
  or (_27840_, _12256_, _27839_);
  and (_27841_, _27840_, _08445_);
  nand (_27842_, _27841_, _27838_);
  and (_27843_, _12265_, _12263_);
  or (_27844_, _27843_, _27808_);
  and (_27845_, _27839_, _07056_);
  nor (_27846_, _27845_, _06653_);
  nor (_27848_, _07056_, \oc8051_golden_model_1.PC [9]);
  nand (_27849_, _27848_, _12265_);
  nand (_27850_, _27849_, _27846_);
  nand (_27851_, _27850_, _24799_);
  and (_27852_, _27851_, _27844_);
  and (_27853_, _27808_, _06653_);
  nor (_27854_, _27853_, _08445_);
  not (_27855_, _27854_);
  nor (_27856_, _27855_, _27852_);
  nor (_27857_, _27856_, _07064_);
  and (_27859_, _27857_, _27842_);
  and (_27860_, _27808_, _07064_);
  or (_27861_, _27860_, _06160_);
  or (_27862_, _27861_, _27859_);
  nand (_27863_, _27862_, _27832_);
  nand (_27864_, _27863_, _12134_);
  nor (_27865_, _27808_, _12134_);
  nor (_27866_, _27865_, _06156_);
  nand (_27867_, _27866_, _27864_);
  and (_27868_, _12172_, _06156_);
  nor (_27870_, _27868_, _07485_);
  nand (_27871_, _27870_, _27867_);
  nand (_27872_, _27871_, _07075_);
  and (_27873_, _12172_, _06217_);
  nor (_27874_, _27873_, _12293_);
  nand (_27875_, _27874_, _27872_);
  nor (_27876_, _27808_, _12292_);
  nor (_27877_, _27876_, _06220_);
  nand (_27878_, _27877_, _27875_);
  and (_27879_, _12172_, _06220_);
  nor (_27881_, _27879_, _12302_);
  nand (_27882_, _27881_, _27878_);
  nor (_27883_, _27808_, _12300_);
  nor (_27884_, _27883_, _06152_);
  nand (_27885_, _27884_, _27882_);
  and (_27886_, _12172_, _06152_);
  nor (_27887_, _27886_, _12304_);
  nand (_27888_, _27887_, _27885_);
  nand (_27889_, _27888_, _07191_);
  and (_27890_, _12172_, _06151_);
  nor (_27892_, _27890_, _12126_);
  nand (_27893_, _27892_, _27889_);
  and (_27894_, _12120_, _11996_);
  nor (_27895_, _27828_, _12120_);
  or (_27896_, _27895_, _27894_);
  nor (_27897_, _27896_, _12125_);
  nor (_27898_, _27897_, _06687_);
  and (_27899_, _27898_, _27893_);
  and (_27900_, _27829_, _11956_);
  and (_27901_, _11996_, _11958_);
  or (_27903_, _27901_, _27900_);
  and (_27904_, _27903_, _06687_);
  or (_27905_, _27904_, _06236_);
  or (_27906_, _27905_, _27899_);
  nor (_27907_, _27828_, _12329_);
  not (_27908_, _27907_);
  and (_27909_, _12329_, _11996_);
  nor (_27910_, _27909_, _06643_);
  and (_27911_, _27910_, _27908_);
  nor (_27912_, _27911_, _06295_);
  nand (_27914_, _27912_, _27906_);
  nand (_27915_, _12346_, _11996_);
  or (_27916_, _27828_, _12346_);
  and (_27917_, _27916_, _27915_);
  or (_27918_, _27917_, _12317_);
  and (_27919_, _27918_, _27914_);
  or (_27920_, _27919_, _11924_);
  nand (_27921_, _27808_, _11924_);
  and (_27922_, _27921_, _27920_);
  nand (_27923_, _27922_, _06146_);
  and (_27925_, _27839_, _06145_);
  nor (_27926_, _27925_, _07388_);
  and (_27927_, _27926_, _25151_);
  nand (_27928_, _27927_, _27923_);
  nor (_27929_, _25151_, _27839_);
  nor (_27930_, _27929_, _12373_);
  nand (_27931_, _27930_, _27928_);
  nor (_27932_, _27808_, _12369_);
  nor (_27933_, _27932_, _06255_);
  and (_27934_, _27933_, _27931_);
  or (_27936_, _27934_, _27822_);
  and (_27937_, _27936_, _27821_);
  or (_27938_, _27937_, _27820_);
  nand (_27939_, _27938_, _12381_);
  and (_27940_, _27808_, _12387_);
  nor (_27941_, _27940_, _12386_);
  nand (_27942_, _27941_, _27939_);
  nor (_27943_, _12172_, _12385_);
  nor (_27944_, _27943_, _05870_);
  nand (_27945_, _27944_, _27942_);
  and (_27947_, _27808_, _05870_);
  nor (_27948_, _27947_, _06139_);
  nand (_27949_, _27948_, _27945_);
  and (_27950_, _27839_, _06139_);
  nor (_27951_, _27950_, _27615_);
  nand (_27952_, _27951_, _27949_);
  and (_27953_, _11996_, _06293_);
  nor (_27954_, _27953_, _13620_);
  nand (_27955_, _27954_, _27952_);
  nor (_27956_, _12172_, _06133_);
  nor (_27958_, _27956_, _05787_);
  nand (_27959_, _27958_, _27955_);
  and (_27960_, _11996_, _05787_);
  nor (_27961_, _27960_, _12412_);
  nand (_27962_, _27961_, _27959_);
  nor (_27963_, _27808_, _11922_);
  nor (_27964_, _27963_, _06209_);
  and (_27965_, _27964_, _27962_);
  or (_27966_, _27965_, _27819_);
  nand (_27967_, _27966_, _27486_);
  nor (_27968_, _27837_, _12417_);
  nor (_27969_, _27968_, _08788_);
  and (_27970_, _27969_, _27967_);
  or (_27971_, _27970_, _27818_);
  nand (_27972_, _27971_, _06111_);
  and (_27973_, _11997_, _06110_);
  nor (_27974_, _27973_, _10751_);
  nand (_27975_, _27974_, _27972_);
  and (_27976_, _12172_, _10751_);
  nor (_27977_, _27976_, _12431_);
  nand (_27980_, _27977_, _27975_);
  nor (_27981_, _12458_, \oc8051_golden_model_1.DPH [1]);
  nor (_27982_, _27981_, _12459_);
  nor (_27983_, _27982_, _12432_);
  nor (_27984_, _27983_, _06208_);
  nand (_27985_, _27984_, _27980_);
  and (_27986_, _12172_, _06208_);
  nor (_27987_, _27986_, _06076_);
  nand (_27988_, _27987_, _27985_);
  nand (_27989_, _27988_, _12474_);
  and (_27991_, _12172_, _11101_);
  nor (_27992_, _27837_, _11101_);
  or (_27993_, _27992_, _27991_);
  and (_27994_, _27993_, _12473_);
  nor (_27995_, _27994_, _12478_);
  and (_27996_, _27995_, _27989_);
  or (_27997_, _27996_, _27817_);
  nand (_27998_, _27997_, _11916_);
  nor (_27999_, _12172_, _11916_);
  nor (_28000_, _27999_, _06297_);
  and (_28002_, _28000_, _27998_);
  or (_28003_, _28002_, _27816_);
  nand (_28004_, _28003_, _07125_);
  and (_28005_, _12172_, _06402_);
  nor (_28006_, _28005_, _12492_);
  nand (_28007_, _28006_, _28004_);
  nand (_28008_, _28007_, _12497_);
  and (_28009_, _12172_, _12480_);
  nor (_28010_, _27837_, _12480_);
  or (_28011_, _28010_, _28009_);
  and (_28013_, _28011_, _12496_);
  nor (_28014_, _28013_, _12505_);
  and (_28015_, _28014_, _28008_);
  or (_28016_, _28015_, _27815_);
  nand (_28017_, _28016_, _10821_);
  nor (_28018_, _12172_, _10821_);
  nor (_28019_, _28018_, _06306_);
  and (_28020_, _28019_, _28017_);
  or (_28021_, _28020_, _27813_);
  nand (_28022_, _28021_, _07130_);
  and (_28024_, _12172_, _06411_);
  nor (_28025_, _28024_, _07124_);
  nand (_28026_, _28025_, _28022_);
  nand (_28027_, _28026_, _12518_);
  and (_28028_, _12172_, \oc8051_golden_model_1.PSW [7]);
  nor (_28029_, _27837_, \oc8051_golden_model_1.PSW [7]);
  or (_28030_, _28029_, _28028_);
  and (_28031_, _28030_, _12517_);
  nor (_28032_, _28031_, _12522_);
  and (_28033_, _28032_, _28027_);
  or (_28035_, _28033_, _27812_);
  nand (_28036_, _28035_, _10849_);
  nor (_28037_, _12172_, _10849_);
  nor (_28038_, _28037_, _06303_);
  and (_28039_, _28038_, _28036_);
  or (_28040_, _28039_, _27811_);
  nand (_28041_, _28040_, _08824_);
  and (_28042_, _12172_, _06396_);
  nor (_28043_, _28042_, _05842_);
  nand (_28044_, _28043_, _28041_);
  nand (_28046_, _28044_, _12539_);
  nand (_28047_, _27837_, \oc8051_golden_model_1.PSW [7]);
  or (_28048_, _12172_, \oc8051_golden_model_1.PSW [7]);
  and (_28049_, _28048_, _12538_);
  and (_28050_, _28049_, _28047_);
  nor (_28051_, _28050_, _12547_);
  and (_28052_, _28051_, _28046_);
  or (_28053_, _28052_, _27810_);
  nand (_28054_, _28053_, _10896_);
  nor (_28055_, _12172_, _10896_);
  nor (_28057_, _28055_, _10925_);
  nand (_28058_, _28057_, _28054_);
  and (_28059_, _27808_, _10925_);
  nor (_28060_, _28059_, _06417_);
  nand (_28061_, _28060_, _28058_);
  nor (_28062_, _06301_, _07142_);
  not (_28063_, _28062_);
  and (_28064_, _07252_, _06417_);
  nor (_28065_, _28064_, _28063_);
  nand (_28066_, _28065_, _28061_);
  nor (_28068_, _11996_, _12682_);
  and (_28069_, _27828_, _12682_);
  or (_28070_, _28069_, _06421_);
  nor (_28071_, _28070_, _28068_);
  nor (_28072_, _28071_, _12565_);
  and (_28073_, _28072_, _28066_);
  or (_28074_, _28073_, _27809_);
  nand (_28075_, _28074_, _12690_);
  nor (_28076_, _12690_, _12172_);
  nor (_28077_, _28076_, _10262_);
  nand (_28079_, _28077_, _28075_);
  and (_28080_, _27808_, _10262_);
  nor (_28081_, _28080_, _06167_);
  nand (_28082_, _28081_, _28079_);
  nor (_28083_, _06165_, _05826_);
  not (_28084_, _28083_);
  and (_28085_, _07252_, _06167_);
  nor (_28086_, _28085_, _28084_);
  nand (_28087_, _28086_, _28082_);
  nor (_28088_, _27829_, _12682_);
  and (_28090_, _11997_, _12682_);
  nor (_28091_, _28090_, _28088_);
  and (_28092_, _28091_, _06165_);
  nor (_28093_, _28092_, _12712_);
  nand (_28094_, _28093_, _28087_);
  nor (_28095_, _27808_, _12711_);
  nor (_28096_, _28095_, _06433_);
  nand (_28097_, _28096_, _28094_);
  and (_28098_, _12172_, _06433_);
  nor (_28099_, _28098_, _25721_);
  nand (_28101_, _28099_, _28097_);
  nor (_28102_, _27808_, _12719_);
  nor (_28103_, _28102_, _06310_);
  and (_28104_, _28103_, _28101_);
  or (_28105_, _28104_, _27806_);
  nand (_28106_, _28105_, _27780_);
  and (_28107_, _28091_, _05748_);
  nor (_28108_, _28107_, _12737_);
  nand (_28109_, _28108_, _28106_);
  nor (_28110_, _27808_, _12735_);
  nor (_28112_, _28110_, _06440_);
  nand (_28113_, _28112_, _28109_);
  and (_28114_, _12172_, _06440_);
  nor (_28115_, _28114_, _26415_);
  nand (_28116_, _28115_, _28113_);
  nor (_28117_, _27808_, _12744_);
  nor (_28118_, _28117_, _06305_);
  and (_28119_, _28118_, _28116_);
  or (_28120_, _28119_, _27805_);
  and (_28121_, _28120_, _27797_);
  and (_28123_, _27808_, _12754_);
  or (_28124_, _28123_, _28121_);
  or (_28125_, _28124_, _01321_);
  or (_28126_, _01317_, \oc8051_golden_model_1.PC [9]);
  and (_28127_, _28126_, _43100_);
  and (_43697_, _28127_, _28125_);
  nor (_28128_, _11896_, \oc8051_golden_model_1.PC [10]);
  nor (_28129_, _28128_, _11897_);
  not (_28130_, _28129_);
  nand (_28131_, _28130_, _10925_);
  nand (_28133_, _11989_, _06303_);
  nand (_28134_, _11989_, _06306_);
  nand (_28135_, _11989_, _06297_);
  nor (_28136_, _12473_, _06076_);
  not (_28137_, _06286_);
  or (_28138_, _28129_, _12292_);
  and (_28139_, _12159_, _07056_);
  and (_28140_, _07057_, \oc8051_golden_model_1.PC [10]);
  and (_28141_, _28140_, _12265_);
  or (_28142_, _28141_, _28139_);
  and (_28144_, _28142_, _12264_);
  or (_28145_, _28144_, _06581_);
  and (_28146_, _28145_, _12263_);
  nor (_28147_, _28130_, _12267_);
  or (_28148_, _28147_, _08445_);
  or (_28149_, _28148_, _28146_);
  and (_28150_, _12258_, _12159_);
  nor (_28151_, _12232_, _12229_);
  not (_28152_, _28151_);
  and (_28153_, _28152_, _12168_);
  nor (_28155_, _28152_, _12168_);
  nor (_28156_, _28155_, _28153_);
  and (_28157_, _28156_, _12256_);
  or (_28158_, _28157_, _28150_);
  or (_28159_, _28158_, _08443_);
  and (_28160_, _28159_, _28149_);
  or (_28161_, _28160_, _07064_);
  nand (_28162_, _28130_, _07064_);
  and (_28163_, _28162_, _06161_);
  and (_28164_, _28163_, _28161_);
  not (_28166_, _11992_);
  nor (_28167_, _12065_, _12062_);
  nor (_28168_, _28167_, _28166_);
  and (_28169_, _28167_, _28166_);
  nor (_28170_, _28169_, _28168_);
  or (_28171_, _28170_, _12141_);
  or (_28172_, _12139_, _11988_);
  and (_28173_, _28172_, _06160_);
  and (_28174_, _28173_, _28171_);
  or (_28175_, _28174_, _24821_);
  or (_28177_, _28175_, _28164_);
  or (_28178_, _28129_, _12134_);
  and (_28179_, _28178_, _06157_);
  and (_28180_, _28179_, _28177_);
  or (_28181_, _28180_, _07485_);
  and (_28182_, _28181_, _07075_);
  not (_28183_, _12159_);
  or (_28184_, _28183_, _06221_);
  nand (_28185_, _28184_, _12292_);
  or (_28186_, _28185_, _28182_);
  and (_28188_, _28186_, _28138_);
  or (_28189_, _28188_, _06220_);
  nand (_28190_, _28183_, _06220_);
  and (_28191_, _28190_, _12300_);
  and (_28192_, _28191_, _28189_);
  nor (_28193_, _28130_, _12300_);
  or (_28194_, _28193_, _28192_);
  and (_28195_, _28194_, _06153_);
  and (_28196_, _12159_, _06152_);
  or (_28197_, _28196_, _12304_);
  or (_28199_, _28197_, _28195_);
  and (_28200_, _28199_, _07191_);
  nand (_28201_, _12159_, _06151_);
  nand (_28202_, _28201_, _12125_);
  or (_28203_, _28202_, _28200_);
  or (_28204_, _28170_, _12120_);
  nand (_28205_, _12120_, _11989_);
  and (_28206_, _28205_, _28204_);
  or (_28207_, _28206_, _12125_);
  and (_28208_, _28207_, _28203_);
  or (_28210_, _28208_, _28137_);
  and (_28211_, _11988_, _11958_);
  and (_28212_, _28170_, _11956_);
  or (_28213_, _28212_, _28211_);
  or (_28214_, _28213_, _12089_);
  and (_28215_, _28214_, _28210_);
  or (_28216_, _28215_, _06236_);
  and (_28217_, _12329_, _11988_);
  and (_28218_, _28170_, _25123_);
  or (_28219_, _28218_, _06643_);
  or (_28221_, _28219_, _28217_);
  and (_28222_, _28221_, _12317_);
  and (_28223_, _28222_, _28216_);
  or (_28224_, _28170_, _12346_);
  nand (_28225_, _12346_, _11989_);
  and (_28226_, _28225_, _06295_);
  and (_28227_, _28226_, _28224_);
  or (_28228_, _28227_, _11924_);
  or (_28229_, _28228_, _28223_);
  nand (_28230_, _28130_, _11924_);
  and (_28232_, _25151_, _06146_);
  and (_28233_, _28232_, _28230_);
  and (_28234_, _28233_, _28229_);
  nor (_28235_, _28232_, _28183_);
  nand (_28236_, _12369_, _05760_);
  or (_28237_, _28236_, _28235_);
  or (_28238_, _28237_, _28234_);
  or (_28239_, _28129_, _12369_);
  and (_28240_, _28239_, _13844_);
  and (_28241_, _28240_, _28238_);
  or (_28243_, _28241_, _24882_);
  and (_28244_, _28243_, _13843_);
  or (_28245_, _28183_, _06256_);
  nand (_28246_, _28245_, _12381_);
  or (_28247_, _28246_, _28244_);
  or (_28248_, _28129_, _12381_);
  and (_28249_, _28248_, _12385_);
  and (_28250_, _28249_, _28247_);
  nor (_28251_, _28183_, _12385_);
  or (_28252_, _28251_, _05870_);
  or (_28254_, _28252_, _28250_);
  or (_28255_, _28129_, _05805_);
  and (_28256_, _28255_, _06140_);
  and (_28257_, _28256_, _28254_);
  nand (_28258_, _12159_, _06139_);
  nand (_28259_, _28258_, _27614_);
  or (_28260_, _28259_, _28257_);
  nand (_28261_, _11989_, _06293_);
  and (_28262_, _28261_, _06133_);
  and (_28263_, _28262_, _28260_);
  nor (_28265_, _28183_, _06133_);
  or (_28266_, _28265_, _05787_);
  or (_28267_, _28266_, _28263_);
  nand (_28268_, _11989_, _05787_);
  and (_28269_, _28268_, _11922_);
  and (_28270_, _28269_, _28267_);
  nor (_28271_, _28130_, _11922_);
  or (_28272_, _28271_, _28270_);
  and (_28273_, _28272_, _06762_);
  nand (_28274_, _12159_, _06209_);
  nand (_28275_, _28274_, _27486_);
  or (_28276_, _28275_, _28273_);
  or (_28277_, _28156_, _12417_);
  and (_28278_, _28277_, _08787_);
  and (_28279_, _28278_, _28276_);
  nor (_28280_, _28183_, _08787_);
  or (_28281_, _28280_, _06110_);
  or (_28282_, _28281_, _28279_);
  nand (_28283_, _11989_, _06110_);
  and (_28284_, _28283_, _10752_);
  and (_28287_, _28284_, _28282_);
  and (_28288_, _12159_, _10751_);
  or (_28289_, _28288_, _12431_);
  or (_28290_, _28289_, _28287_);
  nor (_28291_, _12459_, \oc8051_golden_model_1.DPH [2]);
  nor (_28292_, _28291_, _12460_);
  or (_28293_, _28292_, _12432_);
  and (_28294_, _28293_, _06768_);
  and (_28295_, _28294_, _28290_);
  and (_28296_, _12159_, _06208_);
  or (_28298_, _28296_, _28295_);
  and (_28299_, _28298_, _28136_);
  or (_28300_, _28156_, _11101_);
  or (_28301_, _12159_, _12480_);
  and (_28302_, _28301_, _12473_);
  and (_28303_, _28302_, _28300_);
  or (_28304_, _28303_, _12478_);
  or (_28305_, _28304_, _28299_);
  or (_28306_, _28129_, _11919_);
  and (_28307_, _28306_, _11916_);
  and (_28309_, _28307_, _28305_);
  nor (_28310_, _28183_, _11916_);
  or (_28311_, _28310_, _06297_);
  or (_28312_, _28311_, _28309_);
  and (_28313_, _28312_, _28135_);
  or (_28314_, _28313_, _06402_);
  nand (_28315_, _28183_, _06402_);
  nor (_28316_, _12496_, _12492_);
  and (_28317_, _28316_, _28315_);
  and (_28318_, _28317_, _28314_);
  or (_28320_, _28156_, _12480_);
  or (_28321_, _12159_, _11101_);
  and (_28322_, _28321_, _12496_);
  and (_28323_, _28322_, _28320_);
  or (_28324_, _28323_, _12505_);
  or (_28325_, _28324_, _28318_);
  or (_28326_, _28129_, _11914_);
  and (_28327_, _28326_, _10821_);
  and (_28328_, _28327_, _28325_);
  nor (_28329_, _28183_, _10821_);
  or (_28331_, _28329_, _06306_);
  or (_28332_, _28331_, _28328_);
  and (_28333_, _28332_, _28134_);
  or (_28334_, _28333_, _06411_);
  nand (_28335_, _28183_, _06411_);
  and (_28336_, _28335_, _27696_);
  and (_28337_, _28336_, _28334_);
  or (_28338_, _28156_, \oc8051_golden_model_1.PSW [7]);
  or (_28339_, _12159_, _10693_);
  and (_28340_, _28339_, _12517_);
  and (_28342_, _28340_, _28338_);
  or (_28343_, _28342_, _12522_);
  or (_28344_, _28343_, _28337_);
  or (_28345_, _28129_, _11912_);
  and (_28346_, _28345_, _10849_);
  and (_28347_, _28346_, _28344_);
  nor (_28348_, _28183_, _10849_);
  or (_28349_, _28348_, _06303_);
  or (_28350_, _28349_, _28347_);
  and (_28351_, _28350_, _28133_);
  or (_28353_, _28351_, _06396_);
  nand (_28354_, _28183_, _06396_);
  and (_28355_, _28354_, _27484_);
  and (_28356_, _28355_, _28353_);
  or (_28357_, _28156_, _10693_);
  or (_28358_, _12159_, \oc8051_golden_model_1.PSW [7]);
  and (_28359_, _28358_, _12538_);
  and (_28360_, _28359_, _28357_);
  or (_28361_, _28360_, _12547_);
  or (_28362_, _28361_, _28356_);
  or (_28364_, _28129_, _11907_);
  and (_28365_, _28364_, _10896_);
  and (_28366_, _28365_, _28362_);
  nor (_28367_, _28183_, _10896_);
  or (_28368_, _28367_, _10925_);
  or (_28369_, _28368_, _28366_);
  and (_28370_, _28369_, _28131_);
  or (_28371_, _28370_, _06417_);
  or (_28372_, _07708_, _12558_);
  and (_28373_, _28372_, _28062_);
  and (_28375_, _28373_, _28371_);
  or (_28376_, _28170_, _25333_);
  or (_28377_, _11988_, _12682_);
  and (_28378_, _28377_, _06301_);
  and (_28379_, _28378_, _28376_);
  or (_28380_, _28379_, _12565_);
  or (_28381_, _28380_, _28375_);
  or (_28382_, _28129_, _11905_);
  and (_28383_, _28382_, _12690_);
  and (_28384_, _28383_, _28381_);
  nor (_28386_, _12690_, _28183_);
  or (_28387_, _28386_, _10262_);
  or (_28388_, _28387_, _28384_);
  nand (_28389_, _28130_, _10262_);
  and (_28390_, _28389_, _28388_);
  or (_28391_, _28390_, _06167_);
  or (_28392_, _07708_, _06168_);
  and (_28393_, _28392_, _28083_);
  and (_28394_, _28393_, _28391_);
  nor (_28395_, _28170_, _12682_);
  and (_28397_, _11989_, _12682_);
  nor (_28398_, _28397_, _28395_);
  and (_28399_, _28398_, _06165_);
  or (_28400_, _28399_, _12712_);
  or (_28401_, _28400_, _28394_);
  or (_28402_, _28129_, _12711_);
  and (_28403_, _28402_, _28401_);
  nor (_28404_, _28403_, _06433_);
  and (_28405_, _28183_, _06433_);
  nor (_28406_, _28405_, _25721_);
  not (_28408_, _28406_);
  nor (_28409_, _28408_, _28404_);
  nor (_28410_, _28130_, _12719_);
  nor (_28411_, _28410_, _06310_);
  not (_28412_, _28411_);
  nor (_28413_, _28412_, _28409_);
  not (_28414_, _27780_);
  and (_28415_, _06625_, _06310_);
  nor (_28416_, _28415_, _28414_);
  not (_28417_, _28416_);
  nor (_28419_, _28417_, _28413_);
  and (_28420_, _28398_, _05748_);
  nor (_28421_, _28420_, _12737_);
  not (_28422_, _28421_);
  nor (_28423_, _28422_, _28419_);
  nor (_28424_, _28129_, _12735_);
  or (_28425_, _28424_, _28423_);
  nand (_28426_, _28425_, _06444_);
  and (_28427_, _28183_, _06440_);
  nor (_28428_, _28427_, _26415_);
  and (_28430_, _28428_, _28426_);
  nor (_28431_, _28130_, _12744_);
  or (_28432_, _28431_, _06305_);
  or (_28433_, _28432_, _28430_);
  not (_28434_, _27797_);
  and (_28435_, _06625_, _06305_);
  nor (_28436_, _28435_, _28434_);
  and (_28437_, _28436_, _28433_);
  and (_28438_, _28129_, _12754_);
  or (_28439_, _28438_, _28437_);
  or (_28441_, _28439_, _01321_);
  or (_28442_, _01317_, \oc8051_golden_model_1.PC [10]);
  and (_28443_, _28442_, _43100_);
  and (_43698_, _28443_, _28441_);
  nor (_28444_, _11897_, \oc8051_golden_model_1.PC [11]);
  nor (_28445_, _28444_, _11898_);
  or (_28446_, _28445_, _11905_);
  nor (_28447_, _28153_, _12160_);
  nor (_28448_, _28447_, _12166_);
  and (_28449_, _28447_, _12166_);
  or (_28451_, _28449_, _28448_);
  or (_28452_, _28451_, _10693_);
  or (_28453_, _12163_, \oc8051_golden_model_1.PSW [7]);
  and (_28454_, _28453_, _12538_);
  and (_28455_, _28454_, _28452_);
  or (_28456_, _28451_, \oc8051_golden_model_1.PSW [7]);
  or (_28457_, _12163_, _10693_);
  and (_28458_, _28457_, _12517_);
  and (_28459_, _28458_, _28456_);
  or (_28460_, _28445_, _11914_);
  or (_28462_, _28445_, _11919_);
  or (_28463_, _12163_, _08787_);
  and (_28464_, _11981_, _05787_);
  or (_28465_, _11981_, _11956_);
  nor (_28466_, _28168_, _11990_);
  and (_28467_, _28466_, _11985_);
  nor (_28468_, _28466_, _11985_);
  nor (_28469_, _28468_, _28467_);
  not (_28470_, _28469_);
  or (_28471_, _28470_, _11958_);
  and (_28473_, _28471_, _06687_);
  and (_28474_, _28473_, _28465_);
  nand (_28475_, _12120_, _11982_);
  or (_28476_, _28470_, _12120_);
  and (_28477_, _28476_, _12126_);
  and (_28478_, _28477_, _28475_);
  and (_28479_, _12163_, _06220_);
  or (_28480_, _12131_, _12163_);
  or (_28481_, _12139_, _11981_);
  or (_28482_, _28470_, _12141_);
  and (_28484_, _28482_, _06160_);
  and (_28485_, _28484_, _28481_);
  and (_28486_, _12258_, _12163_);
  and (_28487_, _28451_, _12256_);
  or (_28488_, _28487_, _08443_);
  or (_28489_, _28488_, _28486_);
  or (_28490_, _28445_, _12267_);
  or (_28491_, _12163_, _06582_);
  or (_28492_, _12163_, _07057_);
  nor (_28493_, _07056_, \oc8051_golden_model_1.PC [11]);
  nand (_28495_, _28493_, _12265_);
  and (_28496_, _28495_, _28492_);
  nor (_28497_, _28496_, _06653_);
  nand (_28498_, _28497_, _24799_);
  and (_28499_, _28498_, _28491_);
  and (_28500_, _28499_, _28490_);
  or (_28501_, _28500_, _08445_);
  and (_28502_, _28501_, _12281_);
  and (_28503_, _28502_, _28489_);
  or (_28504_, _28503_, _28485_);
  and (_28506_, _28504_, _12134_);
  and (_28507_, _28445_, _12287_);
  or (_28508_, _28507_, _12286_);
  or (_28509_, _28508_, _28506_);
  and (_28510_, _28509_, _28480_);
  or (_28511_, _28510_, _12293_);
  or (_28512_, _28445_, _12292_);
  and (_28513_, _28512_, _06229_);
  and (_28514_, _28513_, _28511_);
  or (_28515_, _28514_, _28479_);
  and (_28517_, _28515_, _12300_);
  and (_28518_, _28445_, _12302_);
  or (_28519_, _28518_, _12307_);
  or (_28520_, _28519_, _28517_);
  or (_28521_, _12306_, _12163_);
  and (_28522_, _28521_, _12125_);
  and (_28523_, _28522_, _28520_);
  or (_28524_, _28523_, _28478_);
  and (_28525_, _28524_, _12089_);
  or (_28526_, _28525_, _06236_);
  or (_28528_, _28526_, _28474_);
  and (_28529_, _12329_, _11981_);
  nor (_28530_, _28469_, _12329_);
  or (_28531_, _28530_, _06643_);
  or (_28532_, _28531_, _28529_);
  and (_28533_, _28532_, _12317_);
  and (_28534_, _28533_, _28528_);
  nand (_28535_, _28469_, _12347_);
  nand (_28536_, _12346_, _11982_);
  and (_28537_, _28536_, _06295_);
  and (_28539_, _28537_, _28535_);
  or (_28540_, _28539_, _28534_);
  and (_28541_, _28540_, _11925_);
  nand (_28542_, _28445_, _11924_);
  nand (_28543_, _28542_, _12363_);
  or (_28544_, _28543_, _28541_);
  or (_28545_, _12363_, _12163_);
  and (_28546_, _28545_, _12369_);
  and (_28547_, _28546_, _28544_);
  and (_28548_, _28445_, _12373_);
  or (_28550_, _28548_, _12376_);
  or (_28551_, _28550_, _28547_);
  or (_28552_, _12375_, _12163_);
  and (_28553_, _28552_, _12381_);
  and (_28554_, _28553_, _28551_);
  and (_28555_, _28445_, _12387_);
  or (_28556_, _28555_, _12386_);
  or (_28557_, _28556_, _28554_);
  or (_28558_, _12163_, _12385_);
  and (_28559_, _28558_, _05805_);
  and (_28561_, _28559_, _28557_);
  nand (_28562_, _28445_, _05870_);
  nand (_28563_, _28562_, _12395_);
  or (_28564_, _28563_, _28561_);
  or (_28565_, _12395_, _12163_);
  and (_28566_, _28565_, _11296_);
  and (_28567_, _28566_, _28564_);
  nand (_28568_, _11981_, _06293_);
  nand (_28569_, _28568_, _06133_);
  or (_28570_, _28569_, _28567_);
  or (_28572_, _12163_, _06133_);
  and (_28573_, _28572_, _06114_);
  and (_28574_, _28573_, _28570_);
  or (_28575_, _28574_, _28464_);
  and (_28576_, _28575_, _11922_);
  and (_28577_, _28445_, _12412_);
  or (_28578_, _28577_, _12411_);
  or (_28579_, _28578_, _28576_);
  or (_28580_, _12410_, _12163_);
  and (_28581_, _28580_, _12417_);
  and (_28583_, _28581_, _28579_);
  and (_28584_, _28451_, _12416_);
  or (_28585_, _28584_, _08788_);
  or (_28586_, _28585_, _28583_);
  and (_28587_, _28586_, _28463_);
  or (_28588_, _28587_, _06110_);
  nand (_28589_, _11982_, _06110_);
  and (_28590_, _28589_, _10752_);
  and (_28591_, _28590_, _28588_);
  and (_28592_, _12163_, _10751_);
  or (_28594_, _28592_, _28591_);
  and (_28595_, _28594_, _12432_);
  or (_28596_, _12460_, \oc8051_golden_model_1.DPH [3]);
  nor (_28597_, _12461_, _12432_);
  and (_28598_, _28597_, _28596_);
  or (_28599_, _28598_, _12470_);
  or (_28600_, _28599_, _28595_);
  or (_28601_, _12469_, _12163_);
  and (_28602_, _28601_, _12474_);
  and (_28603_, _28602_, _28600_);
  or (_28605_, _28451_, _11101_);
  or (_28606_, _12163_, _12480_);
  and (_28607_, _28606_, _12473_);
  and (_28608_, _28607_, _28605_);
  or (_28609_, _28608_, _12478_);
  or (_28610_, _28609_, _28603_);
  and (_28611_, _28610_, _28462_);
  or (_28612_, _28611_, _11917_);
  or (_28613_, _12163_, _11916_);
  and (_28614_, _28613_, _07127_);
  and (_28616_, _28614_, _28612_);
  nand (_28617_, _11981_, _06297_);
  nand (_28618_, _28617_, _12493_);
  or (_28619_, _28618_, _28616_);
  or (_28620_, _12493_, _12163_);
  and (_28621_, _28620_, _12497_);
  and (_28622_, _28621_, _28619_);
  or (_28623_, _28451_, _12480_);
  or (_28624_, _12163_, _11101_);
  and (_28625_, _28624_, _12496_);
  and (_28626_, _28625_, _28623_);
  or (_28627_, _28626_, _12505_);
  or (_28628_, _28627_, _28622_);
  and (_28629_, _28628_, _28460_);
  or (_28630_, _28629_, _10822_);
  or (_28631_, _12163_, _10821_);
  and (_28632_, _28631_, _07132_);
  and (_28633_, _28632_, _28630_);
  nand (_28634_, _11981_, _06306_);
  nand (_28635_, _28634_, _12514_);
  or (_28638_, _28635_, _28633_);
  or (_28639_, _12514_, _12163_);
  and (_28640_, _28639_, _12518_);
  and (_28641_, _28640_, _28638_);
  or (_28642_, _28641_, _28459_);
  and (_28643_, _28642_, _11912_);
  and (_28644_, _28445_, _12522_);
  or (_28645_, _28644_, _10850_);
  or (_28646_, _28645_, _28643_);
  or (_28647_, _12163_, _10849_);
  and (_28649_, _28647_, _08819_);
  and (_28650_, _28649_, _28646_);
  nand (_28651_, _11981_, _06303_);
  nand (_28652_, _28651_, _12535_);
  or (_28653_, _28652_, _28650_);
  or (_28654_, _12535_, _12163_);
  and (_28655_, _28654_, _12539_);
  and (_28656_, _28655_, _28653_);
  or (_28657_, _28656_, _28455_);
  and (_28658_, _28657_, _11907_);
  and (_28660_, _28445_, _12547_);
  or (_28661_, _28660_, _10897_);
  or (_28662_, _28661_, _28658_);
  or (_28663_, _12163_, _10896_);
  and (_28664_, _28663_, _10926_);
  and (_28665_, _28664_, _28662_);
  and (_28666_, _28445_, _10925_);
  or (_28667_, _28666_, _06417_);
  or (_28668_, _28667_, _28665_);
  or (_28669_, _07544_, _12558_);
  and (_28671_, _28669_, _28668_);
  or (_28672_, _28671_, _07142_);
  nor (_28673_, _12163_, _05846_);
  nor (_28674_, _28673_, _06301_);
  and (_28675_, _28674_, _28672_);
  nand (_28676_, _28469_, _12682_);
  or (_28677_, _11981_, _12682_);
  and (_28678_, _28677_, _06301_);
  and (_28679_, _28678_, _28676_);
  or (_28680_, _28679_, _12565_);
  or (_28682_, _28680_, _28675_);
  and (_28683_, _28682_, _28446_);
  or (_28684_, _28683_, _12691_);
  or (_28685_, _12690_, _12163_);
  and (_28686_, _28685_, _12693_);
  and (_28687_, _28686_, _28684_);
  and (_28688_, _28445_, _10262_);
  or (_28689_, _28688_, _06167_);
  or (_28690_, _28689_, _28687_);
  or (_28691_, _07544_, _06168_);
  and (_28693_, _28691_, _28690_);
  or (_28694_, _28693_, _05826_);
  or (_28695_, _12163_, _12703_);
  and (_28696_, _28695_, _06166_);
  and (_28697_, _28696_, _28694_);
  or (_28698_, _28470_, _12682_);
  nand (_28699_, _11982_, _12682_);
  and (_28700_, _28699_, _28698_);
  and (_28701_, _28700_, _06165_);
  or (_28702_, _28701_, _12712_);
  or (_28704_, _28702_, _28697_);
  or (_28705_, _28445_, _12711_);
  and (_28706_, _28705_, _06829_);
  and (_28707_, _28706_, _28704_);
  nand (_28708_, _12163_, _06433_);
  nand (_28709_, _28708_, _12719_);
  or (_28710_, _28709_, _28707_);
  or (_28711_, _28445_, _12719_);
  and (_28712_, _28711_, _12723_);
  and (_28713_, _28712_, _28710_);
  nor (_28715_, _12723_, _06070_);
  or (_28716_, _28715_, _05823_);
  or (_28717_, _28716_, _28713_);
  or (_28718_, _12163_, _12730_);
  and (_28719_, _28718_, _05749_);
  and (_28720_, _28719_, _28717_);
  and (_28721_, _28700_, _05748_);
  or (_28722_, _28721_, _12737_);
  or (_28723_, _28722_, _28720_);
  or (_28724_, _28445_, _12735_);
  and (_28726_, _28724_, _06444_);
  and (_28727_, _28726_, _28723_);
  nand (_28728_, _12163_, _06440_);
  nand (_28729_, _28728_, _12744_);
  or (_28730_, _28729_, _28727_);
  or (_28731_, _28445_, _12744_);
  and (_28732_, _28731_, _12747_);
  and (_28733_, _28732_, _28730_);
  nor (_28734_, _12747_, _06070_);
  or (_28735_, _28734_, _05821_);
  or (_28737_, _28735_, _28733_);
  or (_28738_, _12163_, _05822_);
  and (_28739_, _28738_, _12755_);
  and (_28740_, _28739_, _28737_);
  and (_28741_, _28445_, _12754_);
  or (_28742_, _28741_, _28740_);
  or (_28743_, _28742_, _01321_);
  or (_28744_, _01317_, \oc8051_golden_model_1.PC [11]);
  and (_28745_, _28744_, _43100_);
  and (_43700_, _28745_, _28743_);
  and (_28747_, _11895_, _09242_);
  and (_28748_, _28747_, \oc8051_golden_model_1.PC [11]);
  and (_28749_, _28748_, \oc8051_golden_model_1.PC [12]);
  nor (_28750_, _28748_, \oc8051_golden_model_1.PC [12]);
  nor (_28751_, _28750_, _28749_);
  not (_28752_, _28751_);
  and (_28753_, _28752_, _12754_);
  and (_28754_, _06876_, _06305_);
  or (_28755_, _28754_, _05821_);
  and (_28756_, _12156_, _10693_);
  and (_28758_, _12239_, _12236_);
  nor (_28759_, _28758_, _12240_);
  and (_28760_, _28759_, \oc8051_golden_model_1.PSW [7]);
  or (_28761_, _28760_, _28756_);
  and (_28762_, _28761_, _12538_);
  and (_28763_, _12156_, \oc8051_golden_model_1.PSW [7]);
  and (_28764_, _28759_, _10693_);
  or (_28765_, _28764_, _28763_);
  and (_28766_, _28765_, _12517_);
  and (_28767_, _12156_, _11101_);
  and (_28769_, _28759_, _12480_);
  or (_28770_, _28769_, _28767_);
  and (_28771_, _28770_, _12473_);
  nor (_28772_, _12156_, _08787_);
  and (_28773_, _11977_, _05787_);
  and (_28774_, _28751_, _11924_);
  and (_28775_, _12072_, _12069_);
  nor (_28776_, _28775_, _12073_);
  not (_28777_, _28776_);
  and (_28778_, _28777_, _11956_);
  nor (_28780_, _11977_, _11956_);
  or (_28781_, _28780_, _12089_);
  or (_28782_, _28781_, _28778_);
  and (_28783_, _12329_, _11977_);
  nor (_28784_, _28777_, _12329_);
  nor (_28785_, _28784_, _28783_);
  nor (_28786_, _28785_, _06643_);
  not (_28787_, _28786_);
  nand (_28788_, _12120_, _11978_);
  or (_28789_, _28776_, _12120_);
  and (_28791_, _28789_, _12126_);
  and (_28792_, _28791_, _28788_);
  or (_28793_, _12139_, _11977_);
  or (_28794_, _28776_, _12141_);
  and (_28795_, _28794_, _06160_);
  nand (_28796_, _28795_, _28793_);
  nand (_28797_, _28759_, _12256_);
  not (_28798_, _12156_);
  or (_28799_, _12256_, _28798_);
  and (_28800_, _28799_, _28797_);
  nand (_28802_, _28800_, _08445_);
  and (_28803_, _12263_, _28798_);
  nor (_28804_, _28751_, _12263_);
  nor (_28805_, _28804_, _28803_);
  nor (_28806_, _28805_, _24799_);
  nor (_28807_, _28752_, _12267_);
  not (_28808_, _28807_);
  and (_28809_, _28798_, _07056_);
  nor (_28810_, _28809_, _06653_);
  not (_28811_, _28810_);
  and (_28813_, _12265_, \oc8051_golden_model_1.PC [12]);
  nor (_28814_, _28813_, _07056_);
  nor (_28815_, _28814_, _28811_);
  nor (_28816_, _28815_, _06581_);
  and (_28817_, _28816_, _28808_);
  nor (_28818_, _28817_, _28806_);
  nor (_28819_, _28818_, _08445_);
  not (_28820_, _28819_);
  and (_28821_, _28820_, _12281_);
  nand (_28822_, _28821_, _28802_);
  nand (_28824_, _28822_, _28796_);
  and (_28825_, _28824_, _12134_);
  and (_28826_, _28751_, _12287_);
  or (_28827_, _28826_, _12286_);
  or (_28828_, _28827_, _28825_);
  nor (_28829_, _12131_, _12156_);
  nor (_28830_, _28829_, _12293_);
  nand (_28831_, _28830_, _28828_);
  nor (_28832_, _28752_, _12292_);
  nor (_28833_, _28832_, _06220_);
  nand (_28835_, _28833_, _28831_);
  and (_28836_, _28798_, _06220_);
  nor (_28837_, _28836_, _12302_);
  nand (_28838_, _28837_, _28835_);
  nor (_28839_, _28752_, _12300_);
  nor (_28840_, _28839_, _12307_);
  nand (_28841_, _28840_, _28838_);
  nor (_28842_, _12306_, _12156_);
  not (_28843_, _28842_);
  and (_28844_, _28843_, _12125_);
  and (_28846_, _28844_, _28841_);
  nor (_28847_, _28846_, _28792_);
  or (_28848_, _28847_, _26862_);
  and (_28849_, _28848_, _28787_);
  nand (_28850_, _28849_, _28782_);
  nand (_28851_, _28850_, _12317_);
  nand (_28852_, _12346_, _11977_);
  nand (_28853_, _28776_, _12347_);
  and (_28854_, _28853_, _28852_);
  or (_28855_, _28854_, _12317_);
  nand (_28857_, _28855_, _28851_);
  nand (_28858_, _28857_, _11925_);
  nand (_28859_, _28858_, _12363_);
  or (_28860_, _28859_, _28774_);
  nor (_28861_, _12363_, _12156_);
  nor (_28862_, _28861_, _12373_);
  nand (_28863_, _28862_, _28860_);
  nor (_28864_, _28752_, _12369_);
  nor (_28865_, _28864_, _12376_);
  nand (_28866_, _28865_, _28863_);
  nor (_28868_, _12375_, _12156_);
  nor (_28869_, _28868_, _12387_);
  nand (_28870_, _28869_, _28866_);
  nor (_28871_, _28752_, _12381_);
  nor (_28872_, _28871_, _12386_);
  nand (_28873_, _28872_, _28870_);
  nor (_28874_, _12156_, _12385_);
  nor (_28875_, _28874_, _05870_);
  nand (_28876_, _28875_, _28873_);
  nor (_28877_, _28752_, _05805_);
  nor (_28879_, _28877_, _12396_);
  nand (_28880_, _28879_, _28876_);
  nor (_28881_, _12395_, _12156_);
  nor (_28882_, _28881_, _06293_);
  nand (_28883_, _28882_, _28880_);
  and (_28884_, _11977_, _06293_);
  nor (_28885_, _28884_, _13620_);
  nand (_28886_, _28885_, _28883_);
  nor (_28887_, _12156_, _06133_);
  nor (_28888_, _28887_, _05787_);
  and (_28890_, _28888_, _28886_);
  or (_28891_, _28890_, _28773_);
  nand (_28892_, _28891_, _11922_);
  nor (_28893_, _28752_, _11922_);
  nor (_28894_, _28893_, _12411_);
  nand (_28895_, _28894_, _28892_);
  nor (_28896_, _12410_, _12156_);
  nor (_28897_, _28896_, _12416_);
  nand (_28898_, _28897_, _28895_);
  and (_28899_, _28759_, _12416_);
  nor (_28901_, _28899_, _08788_);
  and (_28902_, _28901_, _28898_);
  or (_28903_, _28902_, _28772_);
  nand (_28904_, _28903_, _06111_);
  and (_28905_, _11978_, _06110_);
  nor (_28906_, _28905_, _10751_);
  and (_28907_, _28906_, _28904_);
  and (_28908_, _12156_, _10751_);
  or (_28909_, _28908_, _28907_);
  nand (_28910_, _28909_, _12432_);
  nor (_28912_, _12461_, \oc8051_golden_model_1.DPH [4]);
  nor (_28913_, _28912_, _12462_);
  and (_28914_, _28913_, _12431_);
  nor (_28915_, _28914_, _12470_);
  nand (_28916_, _28915_, _28910_);
  nor (_28917_, _12469_, _12156_);
  nor (_28918_, _28917_, _12473_);
  and (_28919_, _28918_, _28916_);
  or (_28920_, _28919_, _28771_);
  nand (_28921_, _28920_, _11919_);
  nor (_28923_, _28752_, _11919_);
  nor (_28924_, _28923_, _11917_);
  nand (_28925_, _28924_, _28921_);
  nor (_28926_, _12156_, _11916_);
  nor (_28927_, _28926_, _06297_);
  nand (_28928_, _28927_, _28925_);
  and (_28929_, _11977_, _06297_);
  not (_28930_, _28929_);
  and (_28931_, _28930_, _12493_);
  nand (_28932_, _28931_, _28928_);
  nor (_28934_, _12493_, _12156_);
  nor (_28935_, _28934_, _12496_);
  and (_28936_, _28935_, _28932_);
  and (_28937_, _12156_, _12480_);
  and (_28938_, _28759_, _11101_);
  or (_28939_, _28938_, _28937_);
  and (_28940_, _28939_, _12496_);
  or (_28941_, _28940_, _28936_);
  nand (_28942_, _28941_, _11914_);
  nor (_28943_, _28752_, _11914_);
  nor (_28945_, _28943_, _10822_);
  nand (_28946_, _28945_, _28942_);
  nor (_28947_, _12156_, _10821_);
  nor (_28948_, _28947_, _06306_);
  nand (_28949_, _28948_, _28946_);
  and (_28950_, _11977_, _06306_);
  not (_28951_, _28950_);
  and (_28952_, _28951_, _12514_);
  nand (_28953_, _28952_, _28949_);
  nor (_28954_, _12514_, _12156_);
  nor (_28956_, _28954_, _12517_);
  and (_28957_, _28956_, _28953_);
  or (_28958_, _28957_, _28766_);
  nand (_28959_, _28958_, _11912_);
  nor (_28960_, _28752_, _11912_);
  nor (_28961_, _28960_, _10850_);
  nand (_28962_, _28961_, _28959_);
  nor (_28963_, _12156_, _10849_);
  nor (_28964_, _28963_, _06303_);
  nand (_28965_, _28964_, _28962_);
  not (_28967_, _12535_);
  and (_28968_, _11977_, _06303_);
  nor (_28969_, _28968_, _28967_);
  nand (_28970_, _28969_, _28965_);
  nor (_28971_, _12535_, _12156_);
  nor (_28972_, _28971_, _12538_);
  and (_28973_, _28972_, _28970_);
  or (_28974_, _28973_, _28762_);
  nand (_28975_, _28974_, _11907_);
  nor (_28976_, _28752_, _11907_);
  nor (_28978_, _28976_, _10897_);
  nand (_28979_, _28978_, _28975_);
  nor (_28980_, _12156_, _10896_);
  nor (_28981_, _28980_, _10925_);
  nand (_28982_, _28981_, _28979_);
  and (_28983_, _28751_, _10925_);
  nor (_28984_, _28983_, _06417_);
  and (_28985_, _28984_, _28982_);
  and (_28986_, _08349_, _06417_);
  or (_28987_, _28986_, _28985_);
  nand (_28989_, _28987_, _05846_);
  nor (_28990_, _12156_, _05846_);
  nor (_28991_, _28990_, _06301_);
  and (_28992_, _28991_, _28989_);
  nor (_28993_, _11978_, _12682_);
  and (_28994_, _28776_, _12682_);
  nor (_28995_, _28994_, _28993_);
  nor (_28996_, _28995_, _06421_);
  or (_28997_, _28996_, _28992_);
  nand (_28998_, _28997_, _11905_);
  nor (_28999_, _28752_, _11905_);
  nor (_29000_, _28999_, _12691_);
  nand (_29001_, _29000_, _28998_);
  nor (_29002_, _12690_, _12156_);
  nor (_29003_, _29002_, _10262_);
  nand (_29004_, _29003_, _29001_);
  and (_29005_, _28751_, _10262_);
  nor (_29006_, _29005_, _06167_);
  nand (_29007_, _29006_, _29004_);
  and (_29008_, _08349_, _06167_);
  nor (_29011_, _29008_, _05826_);
  and (_29012_, _29011_, _29007_);
  and (_29013_, _12156_, _05826_);
  or (_29014_, _29013_, _06165_);
  or (_29015_, _29014_, _29012_);
  and (_29016_, _11978_, _12682_);
  nor (_29017_, _28776_, _12682_);
  nor (_29018_, _29017_, _29016_);
  nor (_29019_, _29018_, _06166_);
  nor (_29020_, _29019_, _12712_);
  nand (_29022_, _29020_, _29015_);
  nor (_29023_, _28752_, _12711_);
  nor (_29024_, _29023_, _06433_);
  nand (_29025_, _29024_, _29022_);
  and (_29026_, _28798_, _06433_);
  nor (_29027_, _29026_, _25721_);
  nand (_29028_, _29027_, _29025_);
  nor (_29029_, _28752_, _12719_);
  nor (_29030_, _29029_, _06310_);
  nand (_29031_, _29030_, _29028_);
  and (_29033_, _06876_, _06310_);
  nor (_29034_, _29033_, _05823_);
  and (_29035_, _29034_, _29031_);
  and (_29036_, _12156_, _05823_);
  or (_29037_, _29036_, _05748_);
  or (_29038_, _29037_, _29035_);
  nor (_29039_, _29018_, _05749_);
  nor (_29040_, _29039_, _12737_);
  nand (_29041_, _29040_, _29038_);
  nor (_29042_, _28752_, _12735_);
  nor (_29044_, _29042_, _06440_);
  nand (_29045_, _29044_, _29041_);
  and (_29046_, _28798_, _06440_);
  nor (_29047_, _29046_, _26415_);
  nand (_29048_, _29047_, _29045_);
  nor (_29049_, _28752_, _12744_);
  nor (_29050_, _29049_, _06305_);
  and (_29051_, _29050_, _29048_);
  or (_29052_, _29051_, _28755_);
  and (_29053_, _12156_, _05821_);
  nor (_29055_, _29053_, _12754_);
  and (_29056_, _29055_, _29052_);
  nor (_29057_, _29056_, _28753_);
  or (_29058_, _29057_, _01321_);
  or (_29059_, _01317_, \oc8051_golden_model_1.PC [12]);
  and (_29060_, _29059_, _43100_);
  and (_43701_, _29060_, _29058_);
  and (_29061_, _12152_, _05823_);
  and (_29062_, _28749_, \oc8051_golden_model_1.PC [13]);
  nor (_29063_, _28749_, \oc8051_golden_model_1.PC [13]);
  nor (_29065_, _29063_, _29062_);
  or (_29066_, _29065_, _12719_);
  or (_29067_, _29065_, _11905_);
  or (_29068_, _29065_, _11912_);
  or (_29069_, _29065_, _11919_);
  and (_29070_, _11972_, _05787_);
  or (_29071_, _11975_, _11974_);
  not (_29072_, _29071_);
  nor (_29073_, _29072_, _12074_);
  and (_29074_, _29072_, _12074_);
  nor (_29076_, _29074_, _29073_);
  not (_29077_, _29076_);
  or (_29078_, _29077_, _11958_);
  or (_29079_, _11972_, _11956_);
  and (_29080_, _29079_, _06687_);
  and (_29081_, _29080_, _29078_);
  and (_29082_, _12152_, _06220_);
  and (_29083_, _29065_, _12287_);
  or (_29084_, _29077_, _12141_);
  or (_29085_, _12139_, _11972_);
  and (_29087_, _29085_, _06160_);
  and (_29088_, _29087_, _29084_);
  or (_29089_, _29065_, _12267_);
  not (_29090_, _12152_);
  nand (_29091_, _29090_, _06581_);
  nand (_29092_, _29090_, _07056_);
  nor (_29093_, _07056_, \oc8051_golden_model_1.PC [13]);
  nand (_29094_, _29093_, _12265_);
  nand (_29095_, _29094_, _29092_);
  and (_29096_, _29095_, _12264_);
  nand (_29098_, _29096_, _24799_);
  and (_29099_, _29098_, _08443_);
  and (_29100_, _29099_, _29091_);
  and (_29101_, _29100_, _29089_);
  or (_29102_, _12256_, _12152_);
  or (_29103_, _12154_, _12153_);
  not (_29104_, _29103_);
  nor (_29105_, _29104_, _12241_);
  and (_29106_, _29104_, _12241_);
  or (_29107_, _29106_, _29105_);
  or (_29109_, _29107_, _12258_);
  and (_29110_, _29109_, _08445_);
  and (_29111_, _29110_, _29102_);
  or (_29112_, _29111_, _29101_);
  and (_29113_, _29112_, _12281_);
  or (_29114_, _29113_, _29088_);
  and (_29115_, _29114_, _12134_);
  or (_29116_, _29115_, _29083_);
  and (_29117_, _29116_, _12131_);
  or (_29118_, _12131_, _29090_);
  nand (_29120_, _29118_, _12292_);
  or (_29121_, _29120_, _29117_);
  or (_29122_, _29065_, _12292_);
  and (_29123_, _29122_, _06229_);
  and (_29124_, _29123_, _29121_);
  or (_29125_, _29124_, _29082_);
  and (_29126_, _29125_, _12300_);
  not (_29127_, _29065_);
  or (_29128_, _29127_, _12300_);
  nand (_29129_, _29128_, _12306_);
  or (_29131_, _29129_, _29126_);
  or (_29132_, _12306_, _12152_);
  and (_29133_, _29132_, _29131_);
  or (_29134_, _29133_, _12126_);
  and (_29135_, _12120_, _11972_);
  nor (_29136_, _29076_, _12120_);
  or (_29137_, _29136_, _29135_);
  or (_29138_, _29137_, _12125_);
  and (_29139_, _29138_, _12089_);
  and (_29140_, _29139_, _29134_);
  or (_29142_, _29140_, _06236_);
  or (_29143_, _29142_, _29081_);
  and (_29144_, _12329_, _11972_);
  nor (_29145_, _29076_, _12329_);
  or (_29146_, _29145_, _06643_);
  or (_29147_, _29146_, _29144_);
  and (_29148_, _29147_, _12317_);
  and (_29149_, _29148_, _29143_);
  nand (_29150_, _29076_, _12347_);
  nand (_29151_, _12346_, _11973_);
  and (_29153_, _29151_, _06295_);
  and (_29154_, _29153_, _29150_);
  or (_29155_, _29154_, _29149_);
  and (_29156_, _29155_, _11925_);
  nand (_29157_, _29065_, _11924_);
  nand (_29158_, _29157_, _12363_);
  or (_29159_, _29158_, _29156_);
  or (_29160_, _12363_, _12152_);
  and (_29161_, _29160_, _12369_);
  and (_29162_, _29161_, _29159_);
  nor (_29164_, _29127_, _12369_);
  or (_29165_, _29164_, _12376_);
  or (_29166_, _29165_, _29162_);
  or (_29167_, _12375_, _12152_);
  and (_29168_, _29167_, _12381_);
  and (_29169_, _29168_, _29166_);
  nor (_29170_, _29127_, _12381_);
  or (_29171_, _29170_, _12386_);
  or (_29172_, _29171_, _29169_);
  or (_29173_, _12152_, _12385_);
  and (_29175_, _29173_, _05805_);
  and (_29176_, _29175_, _29172_);
  or (_29177_, _29127_, _05805_);
  nand (_29178_, _29177_, _12395_);
  or (_29179_, _29178_, _29176_);
  or (_29180_, _12395_, _12152_);
  and (_29181_, _29180_, _11296_);
  and (_29182_, _29181_, _29179_);
  nand (_29183_, _11972_, _06293_);
  nand (_29184_, _29183_, _06133_);
  or (_29186_, _29184_, _29182_);
  or (_29187_, _12152_, _06133_);
  and (_29188_, _29187_, _06114_);
  and (_29189_, _29188_, _29186_);
  or (_29190_, _29189_, _29070_);
  and (_29191_, _29190_, _11922_);
  nor (_29192_, _29127_, _11922_);
  or (_29193_, _29192_, _12411_);
  or (_29194_, _29193_, _29191_);
  or (_29195_, _12410_, _12152_);
  and (_29197_, _29195_, _12417_);
  and (_29198_, _29197_, _29194_);
  and (_29199_, _29107_, _12416_);
  or (_29200_, _29199_, _08788_);
  or (_29201_, _29200_, _29198_);
  or (_29202_, _12152_, _08787_);
  and (_29203_, _29202_, _06111_);
  and (_29204_, _29203_, _29201_);
  and (_29205_, _11972_, _06110_);
  or (_29206_, _29205_, _10751_);
  or (_29208_, _29206_, _29204_);
  nand (_29209_, _29090_, _10751_);
  and (_29210_, _29209_, _12432_);
  and (_29211_, _29210_, _29208_);
  or (_29212_, _12462_, \oc8051_golden_model_1.DPH [5]);
  nor (_29213_, _12463_, _12432_);
  and (_29214_, _29213_, _29212_);
  or (_29215_, _29214_, _12470_);
  or (_29216_, _29215_, _29211_);
  or (_29217_, _12469_, _12152_);
  and (_29219_, _29217_, _12474_);
  and (_29220_, _29219_, _29216_);
  or (_29221_, _29107_, _11101_);
  or (_29222_, _12152_, _12480_);
  and (_29223_, _29222_, _12473_);
  and (_29224_, _29223_, _29221_);
  or (_29225_, _29224_, _12478_);
  or (_29226_, _29225_, _29220_);
  and (_29227_, _29226_, _29069_);
  or (_29228_, _29227_, _11917_);
  or (_29230_, _12152_, _11916_);
  and (_29231_, _29230_, _07127_);
  and (_29232_, _29231_, _29228_);
  nand (_29233_, _11972_, _06297_);
  nand (_29234_, _29233_, _12493_);
  or (_29235_, _29234_, _29232_);
  or (_29236_, _12493_, _12152_);
  and (_29237_, _29236_, _12497_);
  and (_29238_, _29237_, _29235_);
  or (_29239_, _29107_, _12480_);
  or (_29241_, _12152_, _11101_);
  and (_29242_, _29241_, _12496_);
  and (_29243_, _29242_, _29239_);
  or (_29244_, _29243_, _29238_);
  and (_29245_, _29244_, _11914_);
  nor (_29246_, _29127_, _11914_);
  or (_29247_, _29246_, _10822_);
  or (_29248_, _29247_, _29245_);
  or (_29249_, _12152_, _10821_);
  and (_29250_, _29249_, _07132_);
  and (_29252_, _29250_, _29248_);
  nand (_29253_, _11972_, _06306_);
  nand (_29254_, _29253_, _12514_);
  or (_29255_, _29254_, _29252_);
  or (_29256_, _12514_, _12152_);
  and (_29257_, _29256_, _12518_);
  and (_29258_, _29257_, _29255_);
  or (_29259_, _29107_, \oc8051_golden_model_1.PSW [7]);
  or (_29260_, _12152_, _10693_);
  and (_29261_, _29260_, _12517_);
  and (_29263_, _29261_, _29259_);
  or (_29264_, _29263_, _12522_);
  or (_29265_, _29264_, _29258_);
  and (_29266_, _29265_, _29068_);
  or (_29267_, _29266_, _10850_);
  or (_29268_, _12152_, _10849_);
  and (_29269_, _29268_, _08819_);
  and (_29270_, _29269_, _29267_);
  nand (_29271_, _11972_, _06303_);
  nand (_29272_, _29271_, _12535_);
  or (_29274_, _29272_, _29270_);
  or (_29275_, _12535_, _12152_);
  and (_29276_, _29275_, _12539_);
  and (_29277_, _29276_, _29274_);
  or (_29278_, _29107_, _10693_);
  or (_29279_, _12152_, \oc8051_golden_model_1.PSW [7]);
  and (_29280_, _29279_, _12538_);
  and (_29281_, _29280_, _29278_);
  or (_29282_, _29281_, _29277_);
  and (_29283_, _29282_, _11907_);
  nor (_29285_, _29127_, _11907_);
  or (_29286_, _29285_, _10897_);
  or (_29287_, _29286_, _29283_);
  or (_29288_, _12152_, _10896_);
  and (_29289_, _29288_, _10926_);
  and (_29290_, _29289_, _29287_);
  and (_29291_, _29065_, _10925_);
  or (_29292_, _29291_, _06417_);
  or (_29293_, _29292_, _29290_);
  or (_29294_, _08101_, _12558_);
  and (_29296_, _29294_, _29293_);
  or (_29297_, _29296_, _07142_);
  nor (_29298_, _12152_, _05846_);
  nor (_29299_, _29298_, _06301_);
  and (_29300_, _29299_, _29297_);
  or (_29301_, _11972_, _12682_);
  nand (_29302_, _29076_, _12682_);
  and (_29303_, _29302_, _06301_);
  and (_29304_, _29303_, _29301_);
  or (_29305_, _29304_, _12565_);
  or (_29307_, _29305_, _29300_);
  and (_29308_, _29307_, _29067_);
  or (_29309_, _29308_, _12691_);
  or (_29310_, _12690_, _12152_);
  and (_29311_, _29310_, _12693_);
  and (_29312_, _29311_, _29309_);
  and (_29313_, _29065_, _10262_);
  or (_29314_, _29313_, _06167_);
  or (_29315_, _29314_, _29312_);
  or (_29316_, _08101_, _06168_);
  and (_29318_, _29316_, _29315_);
  or (_29319_, _29318_, _05826_);
  nand (_29320_, _29090_, _05826_);
  and (_29321_, _29320_, _06166_);
  and (_29322_, _29321_, _29319_);
  or (_29323_, _29077_, _12682_);
  nand (_29324_, _11973_, _12682_);
  and (_29325_, _29324_, _29323_);
  and (_29326_, _29325_, _06165_);
  or (_29327_, _29326_, _12712_);
  or (_29329_, _29327_, _29322_);
  or (_29330_, _29065_, _12711_);
  and (_29331_, _29330_, _06829_);
  and (_29332_, _29331_, _29329_);
  nand (_29333_, _12152_, _06433_);
  nand (_29334_, _29333_, _12719_);
  or (_29335_, _29334_, _29332_);
  and (_29336_, _29335_, _29066_);
  or (_29337_, _29336_, _06310_);
  nand (_29338_, _06477_, _06310_);
  and (_29340_, _29338_, _12730_);
  and (_29341_, _29340_, _29337_);
  or (_29342_, _29341_, _29061_);
  and (_29343_, _29342_, _05749_);
  and (_29344_, _29325_, _05748_);
  or (_29345_, _29344_, _12737_);
  or (_29346_, _29345_, _29343_);
  or (_29347_, _29065_, _12735_);
  and (_29348_, _29347_, _06444_);
  and (_29349_, _29348_, _29346_);
  nand (_29351_, _12152_, _06440_);
  nand (_29352_, _29351_, _12744_);
  or (_29353_, _29352_, _29349_);
  or (_29354_, _29065_, _12744_);
  and (_29355_, _29354_, _12747_);
  and (_29356_, _29355_, _29353_);
  nor (_29357_, _06477_, _12747_);
  or (_29358_, _29357_, _05821_);
  or (_29359_, _29358_, _29356_);
  nand (_29360_, _29090_, _05821_);
  and (_29362_, _29360_, _12755_);
  and (_29363_, _29362_, _29359_);
  and (_29364_, _29065_, _12754_);
  or (_29365_, _29364_, _29363_);
  or (_29366_, _29365_, _01321_);
  or (_29367_, _01317_, \oc8051_golden_model_1.PC [13]);
  and (_29368_, _29367_, _43100_);
  and (_43702_, _29368_, _29366_);
  and (_29369_, _06305_, _06203_);
  or (_29370_, _29369_, _05821_);
  nor (_29372_, _29062_, \oc8051_golden_model_1.PC [14]);
  nor (_29373_, _29372_, _11901_);
  not (_29374_, _29373_);
  and (_29375_, _29374_, _10262_);
  not (_29376_, _12146_);
  or (_29377_, _12535_, _29376_);
  or (_29378_, _12514_, _29376_);
  or (_29379_, _12493_, _29376_);
  nor (_29380_, _12410_, _12146_);
  and (_29381_, _12076_, _11970_);
  or (_29383_, _29381_, _12077_);
  and (_29384_, _29383_, _11956_);
  nor (_29385_, _11965_, _11956_);
  or (_29386_, _29385_, _12089_);
  or (_29387_, _29386_, _29384_);
  or (_29388_, _29383_, _12329_);
  nand (_29389_, _12329_, _11965_);
  and (_29390_, _29389_, _29388_);
  or (_29391_, _29390_, _06643_);
  and (_29392_, _29376_, _06220_);
  and (_29394_, _29374_, _12287_);
  and (_29395_, _29383_, _12139_);
  and (_29396_, _12141_, _11966_);
  or (_29397_, _29396_, _29395_);
  and (_29398_, _29397_, _06160_);
  nor (_29399_, _29373_, _12263_);
  and (_29400_, _12263_, _29376_);
  or (_29401_, _29400_, _29399_);
  and (_29402_, _29401_, _24800_);
  or (_29403_, _29374_, _12267_);
  and (_29405_, _29376_, _07056_);
  or (_29406_, _29405_, _06653_);
  nand (_29407_, _12265_, \oc8051_golden_model_1.PC [14]);
  and (_29408_, _29407_, _07057_);
  or (_29409_, _29408_, _29406_);
  and (_29410_, _29409_, _06582_);
  and (_29411_, _29410_, _29403_);
  or (_29412_, _29411_, _29402_);
  and (_29413_, _29412_, _08443_);
  or (_29414_, _12256_, _29376_);
  and (_29416_, _12243_, _12150_);
  nor (_29417_, _29416_, _12244_);
  nand (_29418_, _29417_, _12256_);
  and (_29419_, _29418_, _08445_);
  and (_29420_, _29419_, _29414_);
  or (_29421_, _29420_, _29413_);
  and (_29422_, _29421_, _12281_);
  or (_29423_, _29422_, _29398_);
  and (_29424_, _29423_, _12134_);
  or (_29425_, _29424_, _29394_);
  and (_29427_, _29425_, _12131_);
  or (_29428_, _12131_, _12146_);
  nand (_29429_, _29428_, _12292_);
  or (_29430_, _29429_, _29427_);
  or (_29431_, _29374_, _12292_);
  and (_29432_, _29431_, _06229_);
  and (_29433_, _29432_, _29430_);
  or (_29434_, _29433_, _29392_);
  and (_29435_, _29434_, _12300_);
  or (_29436_, _29373_, _12300_);
  nand (_29438_, _29436_, _12306_);
  or (_29439_, _29438_, _29435_);
  or (_29440_, _12306_, _29376_);
  and (_29441_, _29440_, _12125_);
  and (_29442_, _29441_, _29439_);
  nand (_29443_, _12120_, _11965_);
  or (_29444_, _29383_, _12120_);
  and (_29445_, _29444_, _29443_);
  and (_29446_, _29445_, _12126_);
  or (_29447_, _29446_, _26862_);
  or (_29449_, _29447_, _29442_);
  and (_29450_, _29449_, _29391_);
  and (_29451_, _29450_, _29387_);
  or (_29452_, _29451_, _06295_);
  and (_29453_, _29383_, _12347_);
  and (_29454_, _12346_, _11966_);
  or (_29455_, _29454_, _12317_);
  or (_29456_, _29455_, _29453_);
  and (_29457_, _29456_, _11925_);
  and (_29458_, _29457_, _29452_);
  and (_29460_, _29374_, _11924_);
  or (_29461_, _29460_, _29458_);
  and (_29462_, _29461_, _12363_);
  nor (_29463_, _12363_, _12146_);
  or (_29464_, _29463_, _29462_);
  and (_29465_, _29464_, _12369_);
  nor (_29466_, _29373_, _12369_);
  or (_29467_, _29466_, _12376_);
  or (_29468_, _29467_, _29465_);
  or (_29469_, _12375_, _29376_);
  and (_29471_, _29469_, _12381_);
  and (_29472_, _29471_, _29468_);
  nor (_29473_, _29373_, _12381_);
  or (_29474_, _29473_, _12386_);
  or (_29475_, _29474_, _29472_);
  or (_29476_, _29376_, _12385_);
  and (_29477_, _29476_, _05805_);
  and (_29478_, _29477_, _29475_);
  or (_29479_, _29373_, _05805_);
  nand (_29480_, _29479_, _12395_);
  or (_29482_, _29480_, _29478_);
  or (_29483_, _12395_, _29376_);
  and (_29484_, _29483_, _11296_);
  and (_29485_, _29484_, _29482_);
  nand (_29486_, _11966_, _06293_);
  nand (_29487_, _29486_, _06133_);
  or (_29488_, _29487_, _29485_);
  or (_29489_, _29376_, _06133_);
  and (_29490_, _29489_, _06114_);
  and (_29491_, _29490_, _29488_);
  nand (_29493_, _11966_, _05787_);
  nand (_29494_, _29493_, _11922_);
  or (_29495_, _29494_, _29491_);
  or (_29496_, _29374_, _11922_);
  and (_29497_, _29496_, _12410_);
  and (_29498_, _29497_, _29495_);
  or (_29499_, _29498_, _29380_);
  and (_29500_, _29499_, _12417_);
  nor (_29501_, _29417_, _12417_);
  or (_29502_, _29501_, _08788_);
  or (_29504_, _29502_, _29500_);
  or (_29505_, _29376_, _08787_);
  and (_29506_, _29505_, _06111_);
  and (_29507_, _29506_, _29504_);
  and (_29508_, _11966_, _06110_);
  or (_29509_, _29508_, _29507_);
  and (_29510_, _29509_, _10752_);
  and (_29511_, _29376_, _10751_);
  or (_29512_, _29511_, _12431_);
  or (_29513_, _29512_, _29510_);
  nor (_29515_, _12463_, \oc8051_golden_model_1.DPH [6]);
  or (_29516_, _12464_, _12432_);
  or (_29517_, _29516_, _29515_);
  and (_29518_, _29517_, _12469_);
  and (_29519_, _29518_, _29513_);
  nor (_29520_, _12469_, _12146_);
  or (_29521_, _29520_, _12473_);
  or (_29522_, _29521_, _29519_);
  nor (_29523_, _29417_, _11101_);
  or (_29524_, _12146_, _12480_);
  nand (_29525_, _29524_, _12473_);
  or (_29526_, _29525_, _29523_);
  and (_29527_, _29526_, _11919_);
  and (_29528_, _29527_, _29522_);
  nor (_29529_, _29373_, _11919_);
  or (_29530_, _29529_, _11917_);
  or (_29531_, _29530_, _29528_);
  or (_29532_, _29376_, _11916_);
  and (_29533_, _29532_, _07127_);
  and (_29534_, _29533_, _29531_);
  nand (_29537_, _11966_, _06297_);
  nand (_29538_, _29537_, _12493_);
  or (_29539_, _29538_, _29534_);
  and (_29540_, _29539_, _29379_);
  or (_29541_, _29540_, _12496_);
  nor (_29542_, _29417_, _12480_);
  or (_29543_, _12146_, _11101_);
  nand (_29544_, _29543_, _12496_);
  or (_29545_, _29544_, _29542_);
  and (_29546_, _29545_, _11914_);
  and (_29548_, _29546_, _29541_);
  nor (_29549_, _29373_, _11914_);
  or (_29550_, _29549_, _10822_);
  or (_29551_, _29550_, _29548_);
  or (_29552_, _29376_, _10821_);
  and (_29553_, _29552_, _07132_);
  and (_29554_, _29553_, _29551_);
  nand (_29555_, _11966_, _06306_);
  nand (_29556_, _29555_, _12514_);
  or (_29557_, _29556_, _29554_);
  and (_29559_, _29557_, _29378_);
  or (_29560_, _29559_, _12517_);
  nor (_29561_, _29417_, \oc8051_golden_model_1.PSW [7]);
  or (_29562_, _12146_, _10693_);
  nand (_29563_, _29562_, _12517_);
  or (_29564_, _29563_, _29561_);
  and (_29565_, _29564_, _11912_);
  and (_29566_, _29565_, _29560_);
  nor (_29567_, _29373_, _11912_);
  or (_29568_, _29567_, _10850_);
  or (_29570_, _29568_, _29566_);
  or (_29571_, _29376_, _10849_);
  and (_29572_, _29571_, _08819_);
  and (_29573_, _29572_, _29570_);
  nand (_29574_, _11966_, _06303_);
  nand (_29575_, _29574_, _12535_);
  or (_29576_, _29575_, _29573_);
  and (_29577_, _29576_, _29377_);
  or (_29578_, _29577_, _12538_);
  or (_29579_, _29417_, _10693_);
  or (_29581_, _12146_, \oc8051_golden_model_1.PSW [7]);
  and (_29582_, _29581_, _12538_);
  and (_29583_, _29582_, _29579_);
  nor (_29584_, _29583_, _12547_);
  and (_29585_, _29584_, _29578_);
  nor (_29586_, _29373_, _11907_);
  or (_29587_, _29586_, _10897_);
  or (_29588_, _29587_, _29585_);
  or (_29589_, _29376_, _10896_);
  and (_29590_, _29589_, _10926_);
  and (_29592_, _29590_, _29588_);
  and (_29593_, _29374_, _10925_);
  or (_29594_, _29593_, _06417_);
  or (_29595_, _29594_, _29592_);
  or (_29596_, _08347_, _12558_);
  and (_29597_, _29596_, _05846_);
  and (_29598_, _29597_, _29595_);
  nor (_29599_, _12146_, _05846_);
  or (_29600_, _29599_, _06301_);
  or (_29601_, _29600_, _29598_);
  nor (_29603_, _11965_, _12682_);
  and (_29604_, _29383_, _12682_);
  or (_29605_, _29604_, _06421_);
  or (_29606_, _29605_, _29603_);
  and (_29607_, _29606_, _11905_);
  and (_29608_, _29607_, _29601_);
  nor (_29609_, _29373_, _11905_);
  or (_29610_, _29609_, _12691_);
  or (_29611_, _29610_, _29608_);
  or (_29612_, _12690_, _29376_);
  and (_29614_, _29612_, _12693_);
  and (_29615_, _29614_, _29611_);
  or (_29616_, _29615_, _29375_);
  and (_29617_, _29616_, _06168_);
  and (_29618_, _08347_, _06167_);
  or (_29619_, _29618_, _05826_);
  or (_29620_, _29619_, _29617_);
  nand (_29621_, _12146_, _05826_);
  and (_29622_, _29621_, _06166_);
  and (_29623_, _29622_, _29620_);
  nand (_29625_, _11965_, _12682_);
  or (_29626_, _29383_, _12682_);
  and (_29627_, _29626_, _29625_);
  and (_29628_, _29627_, _06165_);
  or (_29629_, _29628_, _29623_);
  and (_29630_, _29629_, _12711_);
  nor (_29631_, _29373_, _12711_);
  or (_29632_, _29631_, _29630_);
  and (_29633_, _29632_, _06829_);
  nand (_29634_, _29376_, _06433_);
  nand (_29636_, _29634_, _12719_);
  or (_29637_, _29636_, _29633_);
  or (_29638_, _29374_, _12719_);
  and (_29639_, _29638_, _12723_);
  and (_29640_, _29639_, _29637_);
  and (_29641_, _06310_, _06203_);
  or (_29642_, _29641_, _05823_);
  or (_29643_, _29642_, _29640_);
  nand (_29644_, _12146_, _05823_);
  and (_29645_, _29644_, _05749_);
  and (_29647_, _29645_, _29643_);
  and (_29648_, _29627_, _05748_);
  or (_29649_, _29648_, _12737_);
  or (_29650_, _29649_, _29647_);
  or (_29651_, _29374_, _12735_);
  and (_29652_, _29651_, _06444_);
  and (_29653_, _29652_, _29650_);
  nand (_29654_, _29376_, _06440_);
  nand (_29655_, _29654_, _12744_);
  or (_29656_, _29655_, _29653_);
  or (_29658_, _29374_, _12744_);
  and (_29659_, _29658_, _12747_);
  and (_29660_, _29659_, _29656_);
  nor (_29661_, _29660_, _29370_);
  and (_29662_, _12146_, _05821_);
  nor (_29663_, _29662_, _29661_);
  or (_29664_, _29663_, _12754_);
  nand (_29665_, _29373_, _12754_);
  and (_29666_, _29665_, _29664_);
  nand (_29667_, _29666_, _01317_);
  or (_29669_, _01317_, \oc8051_golden_model_1.PC [14]);
  and (_29670_, _29669_, _43100_);
  and (_43703_, _29670_, _29667_);
  not (_29671_, _12768_);
  and (_29672_, _29671_, \oc8051_golden_model_1.P2 [0]);
  or (_29673_, _12858_, \oc8051_golden_model_1.ACC [0]);
  nand (_29674_, _12858_, \oc8051_golden_model_1.ACC [0]);
  and (_29675_, _29674_, _29673_);
  and (_29676_, _29675_, _12768_);
  or (_29677_, _29676_, _29672_);
  and (_29679_, _29677_, _06402_);
  and (_29680_, _12768_, _07049_);
  or (_29681_, _29680_, _29672_);
  or (_29682_, _29681_, _06132_);
  nor (_29683_, _12858_, _29671_);
  or (_29684_, _29683_, _29672_);
  or (_29685_, _29684_, _06161_);
  and (_29686_, _12768_, \oc8051_golden_model_1.ACC [0]);
  or (_29687_, _29686_, _29672_);
  and (_29688_, _29687_, _07056_);
  and (_29690_, _07057_, \oc8051_golden_model_1.P2 [0]);
  or (_29691_, _29690_, _06160_);
  or (_29692_, _29691_, _29688_);
  and (_29693_, _29692_, _06157_);
  and (_29694_, _29693_, _29685_);
  not (_29695_, _12773_);
  and (_29696_, _29695_, \oc8051_golden_model_1.P2 [0]);
  and (_29697_, _07847_, \oc8051_golden_model_1.P0 [0]);
  and (_29698_, _12773_, \oc8051_golden_model_1.P2 [0]);
  or (_29699_, _29698_, _29697_);
  and (_29701_, _12778_, \oc8051_golden_model_1.P1 [0]);
  and (_29702_, _12780_, \oc8051_golden_model_1.P3 [0]);
  or (_29703_, _29702_, _29701_);
  or (_29704_, _29703_, _29699_);
  or (_29705_, _14169_, _29704_);
  and (_29706_, _29705_, _12773_);
  or (_29707_, _29706_, _29696_);
  and (_29708_, _29707_, _06156_);
  or (_29709_, _29708_, _29694_);
  and (_29710_, _29709_, _07075_);
  and (_29712_, _29681_, _06217_);
  or (_29713_, _29712_, _06220_);
  or (_29714_, _29713_, _29710_);
  or (_29715_, _29687_, _06229_);
  and (_29716_, _29715_, _06153_);
  and (_29717_, _29716_, _29714_);
  and (_29718_, _29672_, _06152_);
  or (_29719_, _29718_, _06145_);
  or (_29720_, _29719_, _29717_);
  or (_29721_, _29684_, _06146_);
  and (_29723_, _29721_, _06140_);
  and (_29724_, _29723_, _29720_);
  or (_29725_, _29696_, _14170_);
  and (_29726_, _29725_, _06139_);
  and (_29727_, _29726_, _29707_);
  or (_29728_, _29727_, _09842_);
  or (_29729_, _29728_, _29724_);
  and (_29730_, _29729_, _29682_);
  or (_29731_, _29730_, _06116_);
  and (_29732_, _12768_, _09160_);
  or (_29734_, _29672_, _06117_);
  or (_29735_, _29734_, _29732_);
  and (_29736_, _29735_, _06114_);
  and (_29737_, _29736_, _29731_);
  and (_29738_, _12918_, \oc8051_golden_model_1.P1 [0]);
  and (_29739_, _12916_, \oc8051_golden_model_1.P0 [0]);
  and (_29740_, _12920_, \oc8051_golden_model_1.P2 [0]);
  and (_29741_, _12922_, \oc8051_golden_model_1.P3 [0]);
  or (_29742_, _29741_, _29740_);
  or (_29743_, _29742_, _29739_);
  or (_29745_, _29743_, _29738_);
  or (_29746_, _29745_, _14260_);
  and (_29747_, _29746_, _12768_);
  or (_29748_, _29747_, _29672_);
  and (_29749_, _29748_, _05787_);
  or (_29750_, _29749_, _29737_);
  or (_29751_, _29750_, _11136_);
  or (_29752_, _12858_, _08708_);
  and (_29753_, _12858_, _08708_);
  not (_29754_, _29753_);
  and (_29756_, _29754_, _29752_);
  and (_29757_, _29756_, _12768_);
  or (_29758_, _29672_, _07127_);
  or (_29759_, _29758_, _29757_);
  and (_29760_, _12768_, _08708_);
  or (_29761_, _29760_, _29672_);
  or (_29762_, _29761_, _06111_);
  and (_29763_, _29762_, _07125_);
  and (_29764_, _29763_, _29759_);
  and (_29765_, _29764_, _29751_);
  or (_29767_, _29765_, _29679_);
  and (_29768_, _29767_, _07132_);
  nand (_29769_, _29761_, _06306_);
  nor (_29770_, _29769_, _29683_);
  or (_29771_, _29770_, _29768_);
  and (_29772_, _29771_, _07130_);
  or (_29773_, _29672_, _12858_);
  and (_29774_, _29687_, _06411_);
  and (_29775_, _29774_, _29773_);
  or (_29776_, _29775_, _06303_);
  or (_29778_, _29776_, _29772_);
  and (_29779_, _29752_, _12768_);
  or (_29780_, _29672_, _08819_);
  or (_29781_, _29780_, _29779_);
  and (_29782_, _29781_, _08824_);
  and (_29783_, _29782_, _29778_);
  and (_29784_, _29673_, _12768_);
  or (_29785_, _29784_, _29672_);
  and (_29786_, _29785_, _06396_);
  or (_29787_, _29786_, _06433_);
  or (_29789_, _29787_, _29783_);
  or (_29790_, _29684_, _06829_);
  and (_29791_, _29790_, _05749_);
  and (_29792_, _29791_, _29789_);
  and (_29793_, _29672_, _05748_);
  or (_29794_, _29793_, _06440_);
  or (_29795_, _29794_, _29792_);
  or (_29796_, _29684_, _06444_);
  and (_29797_, _29796_, _01317_);
  and (_29798_, _29797_, _29795_);
  nor (_29799_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_29800_, _29799_, _00000_);
  or (_43705_, _29800_, _29798_);
  nor (_29801_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_29802_, _29801_, _00000_);
  and (_29803_, _07847_, \oc8051_golden_model_1.P0 [1]);
  and (_29804_, _12778_, \oc8051_golden_model_1.P1 [1]);
  or (_29805_, _29804_, _29803_);
  and (_29806_, _12773_, \oc8051_golden_model_1.P2 [1]);
  and (_29807_, _12780_, \oc8051_golden_model_1.P3 [1]);
  or (_29810_, _29807_, _29806_);
  or (_29811_, _29810_, _29805_);
  or (_29812_, _29811_, _12627_);
  nand (_29813_, _29812_, _07781_);
  or (_29814_, _14367_, _29811_);
  and (_29815_, _29814_, _12773_);
  and (_29816_, _29815_, _29813_);
  and (_29817_, _29695_, \oc8051_golden_model_1.P2 [1]);
  or (_29818_, _29817_, _06146_);
  or (_29819_, _29818_, _29816_);
  or (_29821_, _12768_, \oc8051_golden_model_1.P2 [1]);
  not (_29822_, _12977_);
  and (_29823_, _29822_, _12859_);
  and (_29824_, _29823_, _12768_);
  not (_29825_, _29824_);
  and (_29826_, _29825_, _29821_);
  or (_29827_, _29826_, _06161_);
  nand (_29828_, _12768_, _05887_);
  and (_29829_, _29828_, _29821_);
  and (_29830_, _29829_, _07056_);
  and (_29832_, _07057_, \oc8051_golden_model_1.P2 [1]);
  or (_29833_, _29832_, _06160_);
  or (_29834_, _29833_, _29830_);
  and (_29835_, _29834_, _06157_);
  and (_29836_, _29835_, _29827_);
  or (_29837_, _29817_, _06217_);
  or (_29838_, _29837_, _29815_);
  and (_29839_, _29838_, _13860_);
  or (_29840_, _29839_, _29836_);
  and (_29841_, _29671_, \oc8051_golden_model_1.P2 [1]);
  and (_29843_, _12768_, _07306_);
  or (_29844_, _29843_, _29841_);
  or (_29845_, _29844_, _07075_);
  and (_29846_, _29845_, _29840_);
  or (_29847_, _29846_, _06220_);
  or (_29848_, _29829_, _06229_);
  and (_29849_, _29848_, _06153_);
  and (_29850_, _29849_, _29847_);
  and (_29851_, _29812_, _14348_);
  and (_29852_, _29851_, _12773_);
  or (_29854_, _29852_, _29817_);
  and (_29855_, _29854_, _06152_);
  or (_29856_, _29855_, _06145_);
  or (_29857_, _29856_, _29850_);
  and (_29858_, _29857_, _29819_);
  and (_29859_, _29858_, _06140_);
  or (_29860_, _29851_, _14350_);
  and (_29861_, _29860_, _12773_);
  or (_29862_, _29817_, _29861_);
  and (_29863_, _29862_, _06139_);
  or (_29865_, _29863_, _09842_);
  or (_29866_, _29865_, _29859_);
  or (_29867_, _29844_, _06132_);
  and (_29868_, _29867_, _29866_);
  or (_29869_, _29868_, _06116_);
  and (_29870_, _12768_, _09115_);
  or (_29871_, _29841_, _06117_);
  or (_29872_, _29871_, _29870_);
  and (_29873_, _29872_, _06114_);
  and (_29874_, _29873_, _29869_);
  and (_29876_, _12916_, \oc8051_golden_model_1.P0 [1]);
  and (_29877_, _12918_, \oc8051_golden_model_1.P1 [1]);
  and (_29878_, _12920_, \oc8051_golden_model_1.P2 [1]);
  and (_29879_, _12922_, \oc8051_golden_model_1.P3 [1]);
  or (_29880_, _29879_, _29878_);
  or (_29881_, _29880_, _29877_);
  or (_29882_, _29881_, _29876_);
  or (_29883_, _29882_, _14442_);
  and (_29884_, _29883_, _12768_);
  or (_29885_, _29884_, _29841_);
  and (_29887_, _29885_, _05787_);
  or (_29888_, _29887_, _29874_);
  and (_29889_, _29888_, _06298_);
  nand (_29890_, _12768_, _06945_);
  and (_29891_, _29821_, _06110_);
  and (_29892_, _29891_, _29890_);
  or (_29893_, _12850_, _08763_);
  and (_29894_, _29893_, _12768_);
  or (_29895_, _29894_, _29841_);
  and (_29896_, _12850_, _08763_);
  not (_29898_, _29896_);
  or (_29899_, _29898_, _29841_);
  and (_29900_, _29899_, _06297_);
  and (_29901_, _29900_, _29895_);
  or (_29902_, _29901_, _29892_);
  or (_29903_, _29902_, _29889_);
  and (_29904_, _29903_, _07125_);
  or (_29905_, _12850_, \oc8051_golden_model_1.ACC [1]);
  and (_29906_, _29905_, _12768_);
  or (_29907_, _29906_, _29841_);
  nand (_29909_, _12850_, \oc8051_golden_model_1.ACC [1]);
  or (_29910_, _29909_, _29841_);
  and (_29911_, _29910_, _06402_);
  and (_29912_, _29911_, _29907_);
  or (_29913_, _29912_, _29904_);
  and (_29914_, _29913_, _07132_);
  or (_29915_, _29896_, _29671_);
  and (_29916_, _29821_, _06306_);
  and (_29917_, _29916_, _29915_);
  or (_29918_, _29917_, _29914_);
  and (_29920_, _29918_, _07130_);
  or (_29921_, _29841_, _12850_);
  and (_29922_, _29829_, _06411_);
  and (_29923_, _29922_, _29921_);
  or (_29924_, _29923_, _06303_);
  or (_29925_, _29924_, _29920_);
  or (_29926_, _29895_, _08819_);
  and (_29927_, _29926_, _08824_);
  and (_29928_, _29927_, _29925_);
  and (_29929_, _29907_, _06396_);
  or (_29931_, _29929_, _06433_);
  or (_29932_, _29931_, _29928_);
  or (_29933_, _29826_, _06829_);
  and (_29934_, _29933_, _05749_);
  and (_29935_, _29934_, _29932_);
  and (_29936_, _29854_, _05748_);
  or (_29937_, _29936_, _06440_);
  or (_29938_, _29937_, _29935_);
  or (_29939_, _29841_, _06444_);
  or (_29940_, _29939_, _29824_);
  and (_29942_, _29940_, _01317_);
  and (_29943_, _29942_, _29938_);
  or (_43706_, _29943_, _29802_);
  and (_29944_, _29671_, \oc8051_golden_model_1.P2 [2]);
  or (_29945_, _12842_, _08768_);
  and (_29946_, _29945_, _12768_);
  or (_29947_, _29946_, _29944_);
  nand (_29948_, _12842_, _08768_);
  or (_29949_, _29948_, _29944_);
  and (_29950_, _29949_, _06297_);
  and (_29952_, _29950_, _29947_);
  and (_29953_, _12859_, _12842_);
  or (_29954_, _29953_, _12860_);
  and (_29955_, _29954_, _12768_);
  or (_29956_, _29955_, _29944_);
  or (_29957_, _29956_, _06161_);
  and (_29958_, _12768_, \oc8051_golden_model_1.ACC [2]);
  or (_29959_, _29958_, _29944_);
  and (_29960_, _29959_, _07056_);
  and (_29961_, _07057_, \oc8051_golden_model_1.P2 [2]);
  or (_29963_, _29961_, _06160_);
  or (_29964_, _29963_, _29960_);
  and (_29965_, _29964_, _06157_);
  and (_29966_, _29965_, _29957_);
  and (_29967_, _29695_, \oc8051_golden_model_1.P2 [2]);
  and (_29968_, _07847_, \oc8051_golden_model_1.P0 [2]);
  and (_29969_, _12773_, \oc8051_golden_model_1.P2 [2]);
  or (_29970_, _29969_, _29968_);
  and (_29971_, _12778_, \oc8051_golden_model_1.P1 [2]);
  and (_29972_, _12780_, \oc8051_golden_model_1.P3 [2]);
  or (_29974_, _29972_, _29971_);
  or (_29975_, _29974_, _29970_);
  or (_29976_, _14538_, _29975_);
  and (_29977_, _29976_, _12773_);
  or (_29978_, _29977_, _29967_);
  and (_29979_, _29978_, _06156_);
  or (_29980_, _29979_, _06217_);
  or (_29981_, _29980_, _29966_);
  and (_29982_, _12768_, _07708_);
  or (_29983_, _29982_, _29944_);
  or (_29985_, _29983_, _07075_);
  and (_29986_, _29985_, _29981_);
  or (_29987_, _29986_, _06220_);
  or (_29988_, _29959_, _06229_);
  and (_29989_, _29988_, _06153_);
  and (_29990_, _29989_, _29987_);
  or (_29991_, _29975_, _12644_);
  and (_29992_, _29991_, _14535_);
  and (_29993_, _29992_, _12773_);
  or (_29994_, _29993_, _29967_);
  and (_29996_, _29994_, _06152_);
  or (_29997_, _29996_, _06145_);
  or (_29998_, _29997_, _29990_);
  nand (_29999_, _29991_, _07848_);
  or (_30000_, _29967_, _29999_);
  and (_30001_, _30000_, _29978_);
  or (_30002_, _30001_, _06146_);
  and (_30003_, _30002_, _06140_);
  and (_30004_, _30003_, _29998_);
  or (_30005_, _29992_, _14582_);
  and (_30007_, _30005_, _12773_);
  or (_30008_, _30007_, _29967_);
  and (_30009_, _30008_, _06139_);
  or (_30010_, _30009_, _09842_);
  or (_30011_, _30010_, _30004_);
  or (_30012_, _29983_, _06132_);
  and (_30013_, _30012_, _30011_);
  or (_30014_, _30013_, _06116_);
  and (_30015_, _12768_, _09211_);
  or (_30016_, _29944_, _06117_);
  or (_30018_, _30016_, _30015_);
  and (_30019_, _30018_, _06114_);
  and (_30020_, _30019_, _30014_);
  and (_30021_, _12916_, \oc8051_golden_model_1.P0 [2]);
  and (_30022_, _12918_, \oc8051_golden_model_1.P1 [2]);
  and (_30023_, _12920_, \oc8051_golden_model_1.P2 [2]);
  and (_30024_, _12922_, \oc8051_golden_model_1.P3 [2]);
  or (_30025_, _30024_, _30023_);
  or (_30026_, _30025_, _30022_);
  or (_30027_, _30026_, _30021_);
  or (_30029_, _30027_, _14630_);
  and (_30030_, _30029_, _12768_);
  or (_30031_, _30030_, _29944_);
  and (_30032_, _30031_, _05787_);
  or (_30033_, _30032_, _06110_);
  or (_30034_, _30033_, _30020_);
  and (_30035_, _12768_, _08768_);
  or (_30036_, _30035_, _29944_);
  or (_30037_, _30036_, _06111_);
  and (_30038_, _30037_, _07127_);
  and (_30040_, _30038_, _30034_);
  or (_30041_, _30040_, _29952_);
  and (_30042_, _30041_, _07125_);
  or (_30043_, _12842_, \oc8051_golden_model_1.ACC [2]);
  and (_30044_, _30043_, _12768_);
  or (_30045_, _30044_, _29944_);
  nand (_30046_, _12842_, \oc8051_golden_model_1.ACC [2]);
  or (_30047_, _30046_, _29944_);
  and (_30048_, _30047_, _06402_);
  and (_30049_, _30048_, _30045_);
  or (_30051_, _30049_, _30042_);
  and (_30052_, _30051_, _07132_);
  or (_30053_, _29944_, _12842_);
  and (_30054_, _30036_, _06306_);
  and (_30055_, _30054_, _30053_);
  or (_30056_, _30055_, _30052_);
  and (_30057_, _30056_, _07130_);
  and (_30058_, _29959_, _06411_);
  and (_30059_, _30058_, _30053_);
  or (_30060_, _30059_, _06303_);
  or (_30062_, _30060_, _30057_);
  or (_30063_, _29947_, _08819_);
  and (_30064_, _30063_, _08824_);
  and (_30065_, _30064_, _30062_);
  and (_30066_, _30045_, _06396_);
  or (_30067_, _30066_, _06433_);
  or (_30068_, _30067_, _30065_);
  or (_30069_, _29956_, _06829_);
  and (_30070_, _30069_, _05749_);
  and (_30071_, _30070_, _30068_);
  and (_30073_, _29994_, _05748_);
  or (_30074_, _30073_, _06440_);
  or (_30075_, _30074_, _30071_);
  nor (_30076_, _12977_, _12842_);
  nor (_30077_, _30076_, _12978_);
  and (_30078_, _30077_, _12768_);
  or (_30079_, _29944_, _06444_);
  or (_30080_, _30079_, _30078_);
  and (_30081_, _30080_, _01317_);
  and (_30082_, _30081_, _30075_);
  nor (_30084_, \oc8051_golden_model_1.P2 [2], rst);
  nor (_30085_, _30084_, _00000_);
  or (_43707_, _30085_, _30082_);
  and (_30086_, _29671_, \oc8051_golden_model_1.P2 [3]);
  and (_30087_, _12768_, _07544_);
  or (_30088_, _30087_, _30086_);
  or (_30089_, _30088_, _06132_);
  and (_30090_, _29695_, \oc8051_golden_model_1.P2 [3]);
  and (_30091_, _07847_, \oc8051_golden_model_1.P0 [3]);
  and (_30092_, _12778_, \oc8051_golden_model_1.P1 [3]);
  or (_30094_, _30092_, _30091_);
  and (_30095_, _12773_, \oc8051_golden_model_1.P2 [3]);
  and (_30096_, _12780_, \oc8051_golden_model_1.P3 [3]);
  or (_30097_, _30096_, _30095_);
  or (_30098_, _30097_, _30094_);
  or (_30099_, _30098_, _12595_);
  and (_30100_, _30099_, _14730_);
  and (_30101_, _30100_, _12773_);
  or (_30102_, _30101_, _30090_);
  and (_30103_, _30102_, _06152_);
  and (_30105_, _12861_, _12834_);
  or (_30106_, _30105_, _12862_);
  and (_30107_, _30106_, _12768_);
  or (_30108_, _30107_, _30086_);
  or (_30109_, _30108_, _06161_);
  and (_30110_, _12768_, \oc8051_golden_model_1.ACC [3]);
  or (_30111_, _30110_, _30086_);
  and (_30112_, _30111_, _07056_);
  and (_30113_, _07057_, \oc8051_golden_model_1.P2 [3]);
  or (_30114_, _30113_, _06160_);
  or (_30116_, _30114_, _30112_);
  and (_30117_, _30116_, _06157_);
  and (_30118_, _30117_, _30109_);
  or (_30119_, _14735_, _30098_);
  and (_30120_, _30119_, _12773_);
  or (_30121_, _30120_, _30090_);
  and (_30122_, _30121_, _06156_);
  or (_30123_, _30122_, _06217_);
  or (_30124_, _30123_, _30118_);
  or (_30125_, _30088_, _07075_);
  and (_30127_, _30125_, _30124_);
  or (_30128_, _30127_, _06220_);
  or (_30129_, _30111_, _06229_);
  and (_30130_, _30129_, _06153_);
  and (_30131_, _30130_, _30128_);
  or (_30132_, _30131_, _30103_);
  and (_30133_, _30132_, _06146_);
  nand (_30134_, _30099_, _07851_);
  or (_30135_, _30090_, _30134_);
  and (_30136_, _30121_, _06145_);
  and (_30138_, _30136_, _30135_);
  or (_30139_, _30138_, _30133_);
  and (_30140_, _30139_, _06140_);
  or (_30141_, _30100_, _14729_);
  and (_30142_, _30141_, _12773_);
  or (_30143_, _30142_, _30090_);
  and (_30144_, _30143_, _06139_);
  or (_30145_, _30144_, _09842_);
  or (_30146_, _30145_, _30140_);
  and (_30147_, _30146_, _30089_);
  or (_30149_, _30147_, _06116_);
  and (_30150_, _12768_, _09210_);
  or (_30151_, _30086_, _06117_);
  or (_30152_, _30151_, _30150_);
  and (_30153_, _30152_, _06114_);
  and (_30154_, _30153_, _30149_);
  and (_30155_, _12916_, \oc8051_golden_model_1.P0 [3]);
  and (_30156_, _12918_, \oc8051_golden_model_1.P1 [3]);
  and (_30157_, _12920_, \oc8051_golden_model_1.P2 [3]);
  and (_30158_, _12922_, \oc8051_golden_model_1.P3 [3]);
  or (_30160_, _30158_, _30157_);
  or (_30161_, _30160_, _30156_);
  or (_30162_, _30161_, _30155_);
  or (_30163_, _30162_, _14825_);
  and (_30164_, _30163_, _12768_);
  or (_30165_, _30164_, _30086_);
  and (_30166_, _30165_, _05787_);
  or (_30167_, _30166_, _06110_);
  or (_30168_, _30167_, _30154_);
  and (_30169_, _12768_, _08712_);
  or (_30171_, _30169_, _30086_);
  or (_30172_, _30171_, _06111_);
  and (_30173_, _30172_, _07127_);
  and (_30174_, _30173_, _30168_);
  or (_30175_, _12834_, _08712_);
  and (_30176_, _30175_, _12768_);
  or (_30177_, _30176_, _30086_);
  nand (_30178_, _12834_, _08712_);
  or (_30179_, _30178_, _30086_);
  and (_30180_, _30179_, _06297_);
  and (_30182_, _30180_, _30177_);
  or (_30183_, _30182_, _30174_);
  and (_30184_, _30183_, _07125_);
  or (_30185_, _12834_, \oc8051_golden_model_1.ACC [3]);
  and (_30186_, _30185_, _12768_);
  or (_30187_, _30186_, _30086_);
  nand (_30188_, _12834_, \oc8051_golden_model_1.ACC [3]);
  or (_30189_, _30188_, _30086_);
  and (_30190_, _30189_, _06402_);
  and (_30191_, _30190_, _30187_);
  or (_30193_, _30191_, _30184_);
  and (_30194_, _30193_, _07132_);
  or (_30195_, _30086_, _12834_);
  and (_30196_, _30171_, _06306_);
  and (_30197_, _30196_, _30195_);
  or (_30198_, _30197_, _30194_);
  and (_30199_, _30198_, _07130_);
  and (_30200_, _30111_, _06411_);
  and (_30201_, _30200_, _30195_);
  or (_30202_, _30201_, _06303_);
  or (_30204_, _30202_, _30199_);
  or (_30205_, _30177_, _08819_);
  and (_30206_, _30205_, _08824_);
  and (_30207_, _30206_, _30204_);
  and (_30208_, _30187_, _06396_);
  or (_30209_, _30208_, _06433_);
  or (_30210_, _30209_, _30207_);
  or (_30211_, _30108_, _06829_);
  and (_30212_, _30211_, _05749_);
  and (_30213_, _30212_, _30210_);
  and (_30215_, _30102_, _05748_);
  or (_30216_, _30215_, _06440_);
  or (_30217_, _30216_, _30213_);
  nor (_30218_, _12978_, _12834_);
  nor (_30219_, _30218_, _12979_);
  and (_30220_, _30219_, _12768_);
  or (_30221_, _30086_, _06444_);
  or (_30222_, _30221_, _30220_);
  and (_30223_, _30222_, _01317_);
  and (_30224_, _30223_, _30217_);
  nor (_30226_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_30227_, _30226_, _00000_);
  or (_43708_, _30227_, _30224_);
  and (_30228_, _29671_, \oc8051_golden_model_1.P2 [4]);
  and (_30229_, _12768_, _08336_);
  or (_30230_, _30229_, _30228_);
  or (_30231_, _30230_, _06132_);
  and (_30232_, _29695_, \oc8051_golden_model_1.P2 [4]);
  and (_30233_, _07847_, \oc8051_golden_model_1.P0 [4]);
  and (_30234_, _12778_, \oc8051_golden_model_1.P1 [4]);
  or (_30236_, _30234_, _30233_);
  and (_30237_, _12773_, \oc8051_golden_model_1.P2 [4]);
  and (_30238_, _12780_, \oc8051_golden_model_1.P3 [4]);
  or (_30239_, _30238_, _30237_);
  nor (_30240_, _30239_, _30236_);
  nand (_30241_, _30240_, _12676_);
  and (_30242_, _30241_, _12678_);
  and (_30243_, _30242_, _12773_);
  or (_30244_, _30243_, _30232_);
  and (_30245_, _30244_, _06152_);
  and (_30247_, _12863_, _12826_);
  or (_30248_, _30247_, _12864_);
  and (_30249_, _30248_, _12768_);
  or (_30250_, _30249_, _30228_);
  or (_30251_, _30250_, _06161_);
  and (_30252_, _12768_, \oc8051_golden_model_1.ACC [4]);
  or (_30253_, _30252_, _30228_);
  and (_30254_, _30253_, _07056_);
  and (_30255_, _07057_, \oc8051_golden_model_1.P2 [4]);
  or (_30256_, _30255_, _06160_);
  or (_30258_, _30256_, _30254_);
  and (_30259_, _30258_, _06157_);
  and (_30260_, _30259_, _30251_);
  or (_30261_, _30241_, _12677_);
  and (_30262_, _30261_, _12773_);
  or (_30263_, _30262_, _30232_);
  and (_30264_, _30263_, _06156_);
  or (_30265_, _30264_, _06217_);
  or (_30266_, _30265_, _30260_);
  or (_30267_, _30230_, _07075_);
  and (_30269_, _30267_, _30266_);
  or (_30270_, _30269_, _06220_);
  or (_30271_, _30253_, _06229_);
  and (_30272_, _30271_, _06153_);
  and (_30273_, _30272_, _30270_);
  or (_30274_, _30273_, _30245_);
  and (_30275_, _30274_, _06146_);
  nand (_30276_, _30241_, _12677_);
  or (_30277_, _30232_, _30276_);
  and (_30278_, _30263_, _06145_);
  and (_30280_, _30278_, _30277_);
  or (_30281_, _30280_, _30275_);
  and (_30282_, _30281_, _06140_);
  or (_30283_, _30242_, _14965_);
  and (_30284_, _30283_, _12773_);
  or (_30285_, _30284_, _30232_);
  and (_30286_, _30285_, _06139_);
  or (_30287_, _30286_, _09842_);
  or (_30288_, _30287_, _30282_);
  and (_30289_, _30288_, _30231_);
  or (_30291_, _30289_, _06116_);
  and (_30292_, _12768_, _09209_);
  or (_30293_, _30228_, _06117_);
  or (_30294_, _30293_, _30292_);
  and (_30295_, _30294_, _06114_);
  and (_30296_, _30295_, _30291_);
  and (_30297_, _12918_, \oc8051_golden_model_1.P1 [4]);
  and (_30298_, _12916_, \oc8051_golden_model_1.P0 [4]);
  and (_30299_, _12920_, \oc8051_golden_model_1.P2 [4]);
  and (_30300_, _12922_, \oc8051_golden_model_1.P3 [4]);
  or (_30302_, _30300_, _30299_);
  or (_30303_, _30302_, _30298_);
  or (_30304_, _30303_, _30297_);
  or (_30305_, _30304_, _15013_);
  and (_30306_, _30305_, _12768_);
  or (_30307_, _30306_, _30228_);
  and (_30308_, _30307_, _05787_);
  or (_30309_, _30308_, _06110_);
  or (_30310_, _30309_, _30296_);
  and (_30311_, _12768_, _08715_);
  or (_30313_, _30311_, _30228_);
  or (_30314_, _30313_, _06111_);
  and (_30315_, _30314_, _07127_);
  and (_30316_, _30315_, _30310_);
  or (_30317_, _12826_, _08715_);
  and (_30318_, _30317_, _12768_);
  or (_30319_, _30318_, _30228_);
  nand (_30320_, _12826_, _08715_);
  or (_30321_, _30320_, _30228_);
  and (_30322_, _30321_, _06297_);
  and (_30324_, _30322_, _30319_);
  or (_30325_, _30324_, _30316_);
  and (_30326_, _30325_, _07125_);
  or (_30327_, _12826_, \oc8051_golden_model_1.ACC [4]);
  and (_30328_, _30327_, _12768_);
  or (_30329_, _30328_, _30228_);
  nand (_30330_, _12826_, \oc8051_golden_model_1.ACC [4]);
  or (_30331_, _30330_, _30228_);
  and (_30332_, _30331_, _06402_);
  and (_30333_, _30332_, _30329_);
  or (_30335_, _30333_, _30326_);
  and (_30336_, _30335_, _07132_);
  or (_30337_, _30228_, _12826_);
  and (_30338_, _30313_, _06306_);
  and (_30339_, _30338_, _30337_);
  or (_30340_, _30339_, _30336_);
  and (_30341_, _30340_, _07130_);
  and (_30342_, _30253_, _06411_);
  and (_30343_, _30342_, _30337_);
  or (_30344_, _30343_, _06303_);
  or (_30346_, _30344_, _30341_);
  or (_30347_, _30319_, _08819_);
  and (_30348_, _30347_, _08824_);
  and (_30349_, _30348_, _30346_);
  and (_30350_, _30329_, _06396_);
  or (_30351_, _30350_, _06433_);
  or (_30352_, _30351_, _30349_);
  or (_30353_, _30250_, _06829_);
  and (_30354_, _30353_, _05749_);
  and (_30355_, _30354_, _30352_);
  and (_30357_, _30244_, _05748_);
  or (_30358_, _30357_, _06440_);
  or (_30359_, _30358_, _30355_);
  nor (_30360_, _12979_, _12826_);
  nor (_30361_, _30360_, _12980_);
  and (_30362_, _30361_, _12768_);
  or (_30363_, _30228_, _06444_);
  or (_30364_, _30363_, _30362_);
  and (_30365_, _30364_, _01317_);
  and (_30366_, _30365_, _30359_);
  nor (_30368_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_30369_, _30368_, _00000_);
  or (_43709_, _30369_, _30366_);
  nor (_30370_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_30371_, _30370_, _00000_);
  and (_30372_, _29671_, \oc8051_golden_model_1.P2 [5]);
  and (_30373_, _12768_, _08101_);
  or (_30374_, _30373_, _30372_);
  or (_30375_, _30374_, _06132_);
  and (_30376_, _12865_, _12818_);
  or (_30378_, _30376_, _12866_);
  and (_30379_, _30378_, _12768_);
  or (_30380_, _30379_, _30372_);
  or (_30381_, _30380_, _06161_);
  and (_30382_, _12768_, \oc8051_golden_model_1.ACC [5]);
  or (_30383_, _30382_, _30372_);
  and (_30384_, _30383_, _07056_);
  and (_30385_, _07057_, \oc8051_golden_model_1.P2 [5]);
  or (_30386_, _30385_, _06160_);
  or (_30387_, _30386_, _30384_);
  and (_30389_, _30387_, _06157_);
  and (_30390_, _30389_, _30381_);
  and (_30391_, _29695_, \oc8051_golden_model_1.P2 [5]);
  and (_30392_, _07847_, \oc8051_golden_model_1.P0 [5]);
  and (_30393_, _12773_, \oc8051_golden_model_1.P2 [5]);
  or (_30394_, _30393_, _30392_);
  and (_30395_, _12778_, \oc8051_golden_model_1.P1 [5]);
  and (_30396_, _12780_, \oc8051_golden_model_1.P3 [5]);
  or (_30397_, _30396_, _30395_);
  or (_30398_, _30397_, _30394_);
  or (_30400_, _15123_, _30398_);
  and (_30401_, _30400_, _12773_);
  or (_30402_, _30401_, _30391_);
  and (_30403_, _30402_, _06156_);
  or (_30404_, _30403_, _06217_);
  or (_30405_, _30404_, _30390_);
  or (_30406_, _30374_, _07075_);
  and (_30407_, _30406_, _30405_);
  or (_30408_, _30407_, _06220_);
  or (_30409_, _30383_, _06229_);
  and (_30411_, _30409_, _06153_);
  and (_30412_, _30411_, _30408_);
  or (_30413_, _30398_, _12611_);
  and (_30414_, _30413_, _15103_);
  and (_30415_, _30414_, _12773_);
  or (_30416_, _30415_, _30391_);
  and (_30417_, _30416_, _06152_);
  or (_30418_, _30417_, _06145_);
  or (_30419_, _30418_, _30412_);
  nand (_30420_, _30413_, _12612_);
  or (_30421_, _30391_, _30420_);
  and (_30422_, _30421_, _30402_);
  or (_30423_, _30422_, _06146_);
  and (_30424_, _30423_, _06140_);
  and (_30425_, _30424_, _30419_);
  or (_30426_, _30414_, _15154_);
  and (_30427_, _30426_, _12773_);
  or (_30428_, _30427_, _30391_);
  and (_30429_, _30428_, _06139_);
  or (_30430_, _30429_, _09842_);
  or (_30433_, _30430_, _30425_);
  and (_30434_, _30433_, _30375_);
  or (_30435_, _30434_, _06116_);
  and (_30436_, _12768_, _09208_);
  or (_30437_, _30372_, _06117_);
  or (_30438_, _30437_, _30436_);
  and (_30439_, _30438_, _06114_);
  and (_30440_, _30439_, _30435_);
  and (_30441_, _12918_, \oc8051_golden_model_1.P1 [5]);
  and (_30442_, _12916_, \oc8051_golden_model_1.P0 [5]);
  and (_30444_, _12920_, \oc8051_golden_model_1.P2 [5]);
  and (_30445_, _12922_, \oc8051_golden_model_1.P3 [5]);
  or (_30446_, _30445_, _30444_);
  or (_30447_, _30446_, _30442_);
  or (_30448_, _30447_, _30441_);
  or (_30449_, _30448_, _15203_);
  and (_30450_, _30449_, _12768_);
  or (_30451_, _30450_, _30372_);
  and (_30452_, _30451_, _05787_);
  or (_30453_, _30452_, _06110_);
  or (_30455_, _30453_, _30440_);
  and (_30456_, _12768_, _08736_);
  or (_30457_, _30456_, _30372_);
  or (_30458_, _30457_, _06111_);
  and (_30459_, _30458_, _07127_);
  and (_30460_, _30459_, _30455_);
  or (_30461_, _12818_, _08736_);
  and (_30462_, _30461_, _12768_);
  or (_30463_, _30462_, _30372_);
  nand (_30464_, _12818_, _08736_);
  or (_30466_, _30464_, _30372_);
  and (_30467_, _30466_, _06297_);
  and (_30468_, _30467_, _30463_);
  or (_30469_, _30468_, _30460_);
  and (_30470_, _30469_, _07125_);
  or (_30471_, _12818_, \oc8051_golden_model_1.ACC [5]);
  and (_30472_, _30471_, _12768_);
  or (_30473_, _30472_, _30372_);
  nand (_30474_, _12818_, \oc8051_golden_model_1.ACC [5]);
  or (_30475_, _30474_, _30372_);
  and (_30477_, _30475_, _06402_);
  and (_30478_, _30477_, _30473_);
  or (_30479_, _30478_, _30470_);
  and (_30480_, _30479_, _07132_);
  or (_30481_, _30372_, _12818_);
  and (_30482_, _30457_, _06306_);
  and (_30483_, _30482_, _30481_);
  or (_30484_, _30483_, _30480_);
  and (_30485_, _30484_, _07130_);
  and (_30486_, _30383_, _06411_);
  and (_30488_, _30486_, _30481_);
  or (_30489_, _30488_, _06303_);
  or (_30490_, _30489_, _30485_);
  or (_30491_, _30463_, _08819_);
  and (_30492_, _30491_, _08824_);
  and (_30493_, _30492_, _30490_);
  and (_30494_, _30473_, _06396_);
  or (_30495_, _30494_, _06433_);
  or (_30496_, _30495_, _30493_);
  or (_30497_, _30380_, _06829_);
  and (_30499_, _30497_, _05749_);
  and (_30500_, _30499_, _30496_);
  and (_30501_, _30416_, _05748_);
  or (_30502_, _30501_, _06440_);
  or (_30503_, _30502_, _30500_);
  nor (_30504_, _12980_, _12818_);
  nor (_30505_, _30504_, _12981_);
  and (_30506_, _30505_, _12768_);
  or (_30507_, _30372_, _06444_);
  or (_30508_, _30507_, _30506_);
  and (_30510_, _30508_, _01317_);
  and (_30511_, _30510_, _30503_);
  or (_43710_, _30511_, _30371_);
  and (_30512_, _29671_, \oc8051_golden_model_1.P2 [6]);
  and (_30513_, _12768_, _08012_);
  or (_30514_, _30513_, _30512_);
  or (_30515_, _30514_, _06132_);
  and (_30516_, _29695_, \oc8051_golden_model_1.P2 [6]);
  and (_30517_, _07847_, \oc8051_golden_model_1.P0 [6]);
  and (_30518_, _12773_, \oc8051_golden_model_1.P2 [6]);
  or (_30520_, _30518_, _30517_);
  and (_30521_, _12778_, \oc8051_golden_model_1.P1 [6]);
  and (_30522_, _12780_, \oc8051_golden_model_1.P3 [6]);
  or (_30523_, _30522_, _30521_);
  or (_30524_, _30523_, _30520_);
  or (_30525_, _30524_, _12579_);
  and (_30526_, _30525_, _15296_);
  and (_30527_, _30526_, _12773_);
  or (_30528_, _30527_, _30516_);
  and (_30529_, _30528_, _06152_);
  and (_30531_, _12867_, _12810_);
  or (_30532_, _30531_, _12868_);
  and (_30533_, _30532_, _12768_);
  or (_30534_, _30533_, _30512_);
  or (_30535_, _30534_, _06161_);
  and (_30536_, _12768_, \oc8051_golden_model_1.ACC [6]);
  or (_30537_, _30536_, _30512_);
  and (_30538_, _30537_, _07056_);
  and (_30539_, _07057_, \oc8051_golden_model_1.P2 [6]);
  or (_30540_, _30539_, _06160_);
  or (_30542_, _30540_, _30538_);
  and (_30543_, _30542_, _06157_);
  and (_30544_, _30543_, _30535_);
  or (_30545_, _15316_, _30524_);
  and (_30546_, _30545_, _12773_);
  or (_30547_, _30546_, _30516_);
  and (_30548_, _30547_, _06156_);
  or (_30549_, _30548_, _06217_);
  or (_30550_, _30549_, _30544_);
  or (_30551_, _30514_, _07075_);
  and (_30553_, _30551_, _30550_);
  or (_30554_, _30553_, _06220_);
  or (_30555_, _30537_, _06229_);
  and (_30556_, _30555_, _06153_);
  and (_30557_, _30556_, _30554_);
  or (_30558_, _30557_, _30529_);
  and (_30559_, _30558_, _06146_);
  nand (_30560_, _30525_, _12580_);
  or (_30561_, _30516_, _30560_);
  and (_30562_, _30547_, _06145_);
  and (_30564_, _30562_, _30561_);
  or (_30565_, _30564_, _30559_);
  and (_30566_, _30565_, _06140_);
  or (_30567_, _30526_, _15347_);
  and (_30568_, _30567_, _12773_);
  or (_30569_, _30568_, _30516_);
  and (_30570_, _30569_, _06139_);
  or (_30571_, _30570_, _09842_);
  or (_30572_, _30571_, _30566_);
  and (_30573_, _30572_, _30515_);
  or (_30575_, _30573_, _06116_);
  and (_30576_, _12768_, _09207_);
  or (_30577_, _30512_, _06117_);
  or (_30578_, _30577_, _30576_);
  and (_30579_, _30578_, _06114_);
  and (_30580_, _30579_, _30575_);
  and (_30581_, _12916_, \oc8051_golden_model_1.P0 [6]);
  and (_30582_, _12918_, \oc8051_golden_model_1.P1 [6]);
  and (_30583_, _12920_, \oc8051_golden_model_1.P2 [6]);
  and (_30584_, _12922_, \oc8051_golden_model_1.P3 [6]);
  or (_30586_, _30584_, _30583_);
  or (_30587_, _30586_, _30582_);
  or (_30588_, _30587_, _30581_);
  or (_30589_, _30588_, _15395_);
  and (_30590_, _30589_, _12768_);
  or (_30591_, _30590_, _30512_);
  and (_30592_, _30591_, _05787_);
  or (_30593_, _30592_, _06110_);
  or (_30594_, _30593_, _30580_);
  and (_30595_, _12768_, _15402_);
  or (_30597_, _30595_, _30512_);
  or (_30598_, _30597_, _06111_);
  and (_30599_, _30598_, _07127_);
  and (_30600_, _30599_, _30594_);
  or (_30601_, _12810_, _15402_);
  and (_30602_, _30601_, _12768_);
  or (_30603_, _30602_, _30512_);
  nand (_30604_, _12810_, _15402_);
  or (_30605_, _30604_, _30512_);
  and (_30606_, _30605_, _06297_);
  and (_30608_, _30606_, _30603_);
  or (_30609_, _30608_, _06402_);
  or (_30610_, _30609_, _30600_);
  or (_30611_, _12810_, \oc8051_golden_model_1.ACC [6]);
  nand (_30612_, _12810_, \oc8051_golden_model_1.ACC [6]);
  and (_30613_, _30612_, _30611_);
  and (_30614_, _30613_, _12768_);
  or (_30615_, _30512_, _07125_);
  or (_30616_, _30615_, _30614_);
  and (_30617_, _30616_, _07132_);
  and (_30619_, _30617_, _30610_);
  or (_30620_, _30512_, _12810_);
  and (_30621_, _30597_, _06306_);
  and (_30622_, _30621_, _30620_);
  or (_30623_, _30622_, _30619_);
  and (_30624_, _30623_, _07130_);
  and (_30625_, _30537_, _06411_);
  and (_30626_, _30625_, _30620_);
  or (_30627_, _30626_, _06303_);
  or (_30628_, _30627_, _30624_);
  or (_30630_, _30603_, _08819_);
  and (_30631_, _30630_, _08824_);
  and (_30632_, _30631_, _30628_);
  and (_30633_, _30611_, _12768_);
  or (_30634_, _30633_, _30512_);
  and (_30635_, _30634_, _06396_);
  or (_30636_, _30635_, _06433_);
  or (_30637_, _30636_, _30632_);
  or (_30638_, _30534_, _06829_);
  and (_30639_, _30638_, _05749_);
  and (_30641_, _30639_, _30637_);
  and (_30642_, _30528_, _05748_);
  or (_30643_, _30642_, _06440_);
  or (_30644_, _30643_, _30641_);
  or (_30645_, _12981_, _12810_);
  and (_30646_, _30645_, _12982_);
  and (_30647_, _30646_, _12768_);
  or (_30648_, _30512_, _06444_);
  or (_30649_, _30648_, _30647_);
  and (_30650_, _30649_, _01317_);
  and (_30652_, _30650_, _30644_);
  nor (_30653_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_30654_, _30653_, _00000_);
  or (_43711_, _30654_, _30652_);
  and (_30655_, _12996_, \oc8051_golden_model_1.P3 [0]);
  and (_30656_, _29705_, _12780_);
  or (_30657_, _30656_, _30655_);
  or (_30658_, _30657_, _06157_);
  and (_30659_, _12991_, \oc8051_golden_model_1.P3 [0]);
  nor (_30660_, _12858_, _12991_);
  or (_30662_, _30660_, _30659_);
  and (_30663_, _30662_, _06160_);
  and (_30664_, _07057_, \oc8051_golden_model_1.P3 [0]);
  and (_30665_, _12797_, \oc8051_golden_model_1.ACC [0]);
  or (_30666_, _30665_, _30659_);
  and (_30667_, _30666_, _07056_);
  or (_30668_, _30667_, _30664_);
  and (_30669_, _30668_, _06161_);
  or (_30670_, _30669_, _06156_);
  or (_30671_, _30670_, _30663_);
  and (_30673_, _30671_, _30658_);
  and (_30674_, _30673_, _07075_);
  and (_30675_, _12797_, _07049_);
  or (_30676_, _30675_, _30659_);
  and (_30677_, _30676_, _06217_);
  or (_30678_, _30677_, _06220_);
  or (_30679_, _30678_, _30674_);
  or (_30680_, _30666_, _06229_);
  and (_30681_, _30680_, _06153_);
  and (_30682_, _30681_, _30679_);
  and (_30684_, _30659_, _06152_);
  or (_30685_, _30684_, _06145_);
  or (_30686_, _30685_, _30682_);
  or (_30687_, _30662_, _06146_);
  and (_30688_, _30687_, _06140_);
  and (_30689_, _30688_, _30686_);
  or (_30690_, _30655_, _14170_);
  and (_30691_, _30690_, _06139_);
  and (_30692_, _30691_, _30657_);
  or (_30693_, _30692_, _09842_);
  or (_30695_, _30693_, _30689_);
  or (_30696_, _30676_, _06132_);
  and (_30697_, _30696_, _30695_);
  or (_30698_, _30697_, _06116_);
  and (_30699_, _12797_, _09160_);
  or (_30700_, _30659_, _06117_);
  or (_30701_, _30700_, _30699_);
  and (_30702_, _30701_, _06114_);
  and (_30703_, _30702_, _30698_);
  and (_30704_, _29746_, _12797_);
  or (_30706_, _30704_, _30659_);
  and (_30707_, _30706_, _05787_);
  or (_30708_, _30707_, _06110_);
  or (_30709_, _30708_, _30703_);
  and (_30710_, _12797_, _08708_);
  or (_30711_, _30710_, _30659_);
  or (_30712_, _30711_, _06111_);
  and (_30713_, _30712_, _07127_);
  and (_30714_, _30713_, _30709_);
  and (_30715_, _29752_, _12797_);
  or (_30717_, _30715_, _30659_);
  or (_30718_, _30659_, _29754_);
  and (_30719_, _30718_, _06297_);
  and (_30720_, _30719_, _30717_);
  or (_30721_, _30720_, _06402_);
  or (_30722_, _30721_, _30714_);
  and (_30723_, _29675_, _12797_);
  or (_30724_, _30659_, _07125_);
  or (_30725_, _30724_, _30723_);
  and (_30726_, _30725_, _07132_);
  and (_30728_, _30726_, _30722_);
  nand (_30729_, _30711_, _06306_);
  nor (_30730_, _30729_, _30660_);
  or (_30731_, _30730_, _30728_);
  and (_30732_, _30731_, _07130_);
  or (_30733_, _30659_, _12858_);
  and (_30734_, _30666_, _06411_);
  and (_30735_, _30734_, _30733_);
  or (_30736_, _30735_, _06303_);
  or (_30737_, _30736_, _30732_);
  or (_30739_, _30717_, _08819_);
  and (_30740_, _30739_, _08824_);
  and (_30741_, _30740_, _30737_);
  and (_30742_, _29673_, _12797_);
  or (_30743_, _30742_, _30659_);
  and (_30744_, _30743_, _06396_);
  or (_30745_, _30744_, _06433_);
  or (_30746_, _30745_, _30741_);
  or (_30747_, _30662_, _06829_);
  and (_30748_, _30747_, _05749_);
  and (_30750_, _30748_, _30746_);
  and (_30751_, _30659_, _05748_);
  or (_30752_, _30751_, _06440_);
  or (_30753_, _30752_, _30750_);
  or (_30754_, _30662_, _06444_);
  and (_30755_, _30754_, _01317_);
  and (_30756_, _30755_, _30753_);
  nor (_30757_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_30758_, _30757_, _00000_);
  or (_43713_, _30758_, _30756_);
  nor (_30760_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_30761_, _30760_, _00000_);
  or (_30762_, _29883_, _12991_);
  or (_30763_, _12797_, \oc8051_golden_model_1.P3 [1]);
  and (_30764_, _30763_, _05787_);
  and (_30765_, _30764_, _30762_);
  and (_30766_, _29814_, _12780_);
  and (_30767_, _30766_, _29813_);
  and (_30768_, _12996_, \oc8051_golden_model_1.P3 [1]);
  or (_30769_, _30768_, _06146_);
  or (_30771_, _30769_, _30767_);
  and (_30772_, _29823_, _12797_);
  not (_30773_, _30772_);
  and (_30774_, _30773_, _30763_);
  or (_30775_, _30774_, _06161_);
  nand (_30776_, _12797_, _05887_);
  and (_30777_, _30776_, _30763_);
  and (_30778_, _30777_, _07056_);
  and (_30779_, _07057_, \oc8051_golden_model_1.P3 [1]);
  or (_30780_, _30779_, _06160_);
  or (_30782_, _30780_, _30778_);
  and (_30783_, _30782_, _06157_);
  and (_30784_, _30783_, _30775_);
  or (_30785_, _30768_, _06217_);
  or (_30786_, _30785_, _30766_);
  and (_30787_, _30786_, _13860_);
  or (_30788_, _30787_, _30784_);
  and (_30789_, _12991_, \oc8051_golden_model_1.P3 [1]);
  and (_30790_, _12797_, _07306_);
  or (_30791_, _30790_, _30789_);
  or (_30793_, _30791_, _07075_);
  and (_30794_, _30793_, _30788_);
  or (_30795_, _30794_, _06220_);
  or (_30796_, _30777_, _06229_);
  and (_30797_, _30796_, _06153_);
  and (_30798_, _30797_, _30795_);
  and (_30799_, _29851_, _12780_);
  or (_30800_, _30799_, _30768_);
  and (_30801_, _30800_, _06152_);
  or (_30802_, _30801_, _06145_);
  or (_30804_, _30802_, _30798_);
  and (_30805_, _30804_, _30771_);
  and (_30806_, _30805_, _06140_);
  and (_30807_, _29860_, _12780_);
  or (_30808_, _30768_, _30807_);
  and (_30809_, _30808_, _06139_);
  or (_30810_, _30809_, _09842_);
  or (_30811_, _30810_, _30806_);
  or (_30812_, _30791_, _06132_);
  and (_30813_, _30812_, _30811_);
  or (_30815_, _30813_, _06116_);
  and (_30816_, _12797_, _09115_);
  or (_30817_, _30789_, _06117_);
  or (_30818_, _30817_, _30816_);
  and (_30819_, _30818_, _06114_);
  and (_30820_, _30819_, _30815_);
  or (_30821_, _30820_, _30765_);
  and (_30822_, _30821_, _06298_);
  and (_30823_, _29898_, _29893_);
  or (_30824_, _30823_, _12991_);
  and (_30826_, _30824_, _06297_);
  nand (_30827_, _12797_, _06945_);
  and (_30828_, _30827_, _06110_);
  or (_30829_, _30828_, _30826_);
  and (_30830_, _30829_, _30763_);
  or (_30831_, _30830_, _30822_);
  and (_30832_, _30831_, _07125_);
  and (_30833_, _29909_, _29905_);
  or (_30834_, _30833_, _12991_);
  and (_30835_, _30763_, _06402_);
  and (_30837_, _30835_, _30834_);
  or (_30838_, _30837_, _30832_);
  and (_30839_, _30838_, _07132_);
  or (_30840_, _29896_, _12991_);
  and (_30841_, _30763_, _06306_);
  and (_30842_, _30841_, _30840_);
  or (_30843_, _30842_, _30839_);
  and (_30844_, _30843_, _07130_);
  or (_30845_, _30789_, _12850_);
  and (_30846_, _30777_, _06411_);
  and (_30848_, _30846_, _30845_);
  or (_30849_, _30848_, _30844_);
  and (_30850_, _30849_, _06397_);
  or (_30851_, _30827_, _12850_);
  and (_30852_, _30763_, _06303_);
  and (_30853_, _30852_, _30851_);
  or (_30854_, _30776_, _12850_);
  and (_30855_, _30763_, _06396_);
  and (_30856_, _30855_, _30854_);
  or (_30857_, _30856_, _06433_);
  or (_30859_, _30857_, _30853_);
  or (_30860_, _30859_, _30850_);
  or (_30861_, _30774_, _06829_);
  and (_30862_, _30861_, _05749_);
  and (_30863_, _30862_, _30860_);
  and (_30864_, _30800_, _05748_);
  or (_30865_, _30864_, _06440_);
  or (_30866_, _30865_, _30863_);
  or (_30867_, _30789_, _06444_);
  or (_30868_, _30867_, _30772_);
  and (_30870_, _30868_, _01317_);
  and (_30871_, _30870_, _30866_);
  or (_43714_, _30871_, _30761_);
  and (_30872_, _12991_, \oc8051_golden_model_1.P3 [2]);
  and (_30873_, _29954_, _12797_);
  or (_30874_, _30873_, _30872_);
  or (_30875_, _30874_, _06161_);
  and (_30876_, _12797_, \oc8051_golden_model_1.ACC [2]);
  or (_30877_, _30876_, _30872_);
  and (_30878_, _30877_, _07056_);
  and (_30880_, _07057_, \oc8051_golden_model_1.P3 [2]);
  or (_30881_, _30880_, _06160_);
  or (_30882_, _30881_, _30878_);
  and (_30883_, _30882_, _06157_);
  and (_30884_, _30883_, _30875_);
  and (_30885_, _12996_, \oc8051_golden_model_1.P3 [2]);
  and (_30886_, _29976_, _12780_);
  or (_30887_, _30886_, _30885_);
  and (_30888_, _30887_, _06156_);
  or (_30889_, _30888_, _06217_);
  or (_30891_, _30889_, _30884_);
  and (_30892_, _12797_, _07708_);
  or (_30893_, _30892_, _30872_);
  or (_30894_, _30893_, _07075_);
  and (_30895_, _30894_, _30891_);
  or (_30896_, _30895_, _06220_);
  or (_30897_, _30877_, _06229_);
  and (_30898_, _30897_, _06153_);
  and (_30899_, _30898_, _30896_);
  and (_30900_, _29992_, _12780_);
  or (_30902_, _30900_, _30885_);
  and (_30903_, _30902_, _06152_);
  or (_30904_, _30903_, _06145_);
  or (_30905_, _30904_, _30899_);
  or (_30906_, _30885_, _29999_);
  and (_30907_, _30906_, _30887_);
  or (_30908_, _30907_, _06146_);
  and (_30909_, _30908_, _06140_);
  and (_30910_, _30909_, _30905_);
  and (_30911_, _30005_, _12780_);
  or (_30913_, _30911_, _30885_);
  and (_30914_, _30913_, _06139_);
  or (_30915_, _30914_, _09842_);
  or (_30916_, _30915_, _30910_);
  or (_30917_, _30893_, _06132_);
  and (_30918_, _30917_, _30916_);
  or (_30919_, _30918_, _06116_);
  and (_30920_, _12797_, _09211_);
  or (_30921_, _30872_, _06117_);
  or (_30922_, _30921_, _30920_);
  and (_30924_, _30922_, _06114_);
  and (_30925_, _30924_, _30919_);
  and (_30926_, _30029_, _12797_);
  or (_30927_, _30926_, _30872_);
  and (_30928_, _30927_, _05787_);
  or (_30929_, _30928_, _06110_);
  or (_30930_, _30929_, _30925_);
  and (_30931_, _12797_, _08768_);
  or (_30932_, _30931_, _30872_);
  or (_30933_, _30932_, _06111_);
  and (_30935_, _30933_, _07127_);
  and (_30936_, _30935_, _30930_);
  and (_30937_, _29945_, _12797_);
  or (_30938_, _30937_, _30872_);
  or (_30939_, _30872_, _29948_);
  and (_30940_, _30939_, _06297_);
  and (_30941_, _30940_, _30938_);
  or (_30942_, _30941_, _30936_);
  and (_30943_, _30942_, _07125_);
  and (_30944_, _30043_, _12797_);
  or (_30946_, _30944_, _30872_);
  or (_30947_, _30872_, _30046_);
  and (_30948_, _30947_, _06402_);
  and (_30949_, _30948_, _30946_);
  or (_30950_, _30949_, _30943_);
  and (_30951_, _30950_, _07132_);
  or (_30952_, _30872_, _12842_);
  and (_30953_, _30932_, _06306_);
  and (_30954_, _30953_, _30952_);
  or (_30955_, _30954_, _30951_);
  and (_30957_, _30955_, _07130_);
  and (_30958_, _30877_, _06411_);
  and (_30959_, _30958_, _30952_);
  or (_30960_, _30959_, _06303_);
  or (_30961_, _30960_, _30957_);
  or (_30962_, _30938_, _08819_);
  and (_30963_, _30962_, _08824_);
  and (_30964_, _30963_, _30961_);
  and (_30965_, _30946_, _06396_);
  or (_30966_, _30965_, _06433_);
  or (_30968_, _30966_, _30964_);
  or (_30969_, _30874_, _06829_);
  and (_30970_, _30969_, _05749_);
  and (_30971_, _30970_, _30968_);
  and (_30972_, _30902_, _05748_);
  or (_30973_, _30972_, _06440_);
  or (_30974_, _30973_, _30971_);
  and (_30975_, _30077_, _12797_);
  or (_30976_, _30872_, _06444_);
  or (_30977_, _30976_, _30975_);
  and (_30979_, _30977_, _01317_);
  and (_30980_, _30979_, _30974_);
  nor (_30981_, \oc8051_golden_model_1.P3 [2], rst);
  nor (_30982_, _30981_, _00000_);
  or (_43715_, _30982_, _30980_);
  and (_30983_, _12991_, \oc8051_golden_model_1.P3 [3]);
  and (_30984_, _12797_, _07544_);
  or (_30985_, _30984_, _30983_);
  or (_30986_, _30985_, _06132_);
  and (_30987_, _12996_, \oc8051_golden_model_1.P3 [3]);
  and (_30989_, _30100_, _12780_);
  or (_30990_, _30989_, _30987_);
  and (_30991_, _30990_, _06152_);
  and (_30992_, _30106_, _12797_);
  or (_30993_, _30992_, _30983_);
  or (_30994_, _30993_, _06161_);
  and (_30995_, _12797_, \oc8051_golden_model_1.ACC [3]);
  or (_30996_, _30995_, _30983_);
  and (_30997_, _30996_, _07056_);
  and (_30998_, _07057_, \oc8051_golden_model_1.P3 [3]);
  or (_31000_, _30998_, _06160_);
  or (_31001_, _31000_, _30997_);
  and (_31002_, _31001_, _06157_);
  and (_31003_, _31002_, _30994_);
  and (_31004_, _30119_, _12780_);
  or (_31005_, _31004_, _30987_);
  and (_31006_, _31005_, _06156_);
  or (_31007_, _31006_, _06217_);
  or (_31008_, _31007_, _31003_);
  or (_31009_, _30985_, _07075_);
  and (_31011_, _31009_, _31008_);
  or (_31012_, _31011_, _06220_);
  or (_31013_, _30996_, _06229_);
  and (_31014_, _31013_, _06153_);
  and (_31015_, _31014_, _31012_);
  or (_31016_, _31015_, _30991_);
  and (_31017_, _31016_, _06146_);
  or (_31018_, _30987_, _30134_);
  and (_31019_, _31005_, _06145_);
  and (_31020_, _31019_, _31018_);
  or (_31022_, _31020_, _31017_);
  and (_31023_, _31022_, _06140_);
  and (_31024_, _30141_, _12780_);
  or (_31025_, _31024_, _30987_);
  and (_31026_, _31025_, _06139_);
  or (_31027_, _31026_, _09842_);
  or (_31028_, _31027_, _31023_);
  and (_31029_, _31028_, _30986_);
  or (_31030_, _31029_, _06116_);
  and (_31031_, _12797_, _09210_);
  or (_31033_, _30983_, _06117_);
  or (_31034_, _31033_, _31031_);
  and (_31035_, _31034_, _06114_);
  and (_31036_, _31035_, _31030_);
  and (_31037_, _30163_, _12797_);
  or (_31038_, _31037_, _30983_);
  and (_31039_, _31038_, _05787_);
  or (_31040_, _31039_, _11136_);
  or (_31041_, _31040_, _31036_);
  and (_31042_, _30178_, _30175_);
  and (_31044_, _31042_, _12797_);
  or (_31045_, _30983_, _07127_);
  or (_31046_, _31045_, _31044_);
  and (_31047_, _12797_, _08712_);
  or (_31048_, _31047_, _30983_);
  or (_31049_, _31048_, _06111_);
  and (_31050_, _31049_, _07125_);
  and (_31051_, _31050_, _31046_);
  and (_31052_, _31051_, _31041_);
  and (_31053_, _30188_, _30185_);
  and (_31055_, _31053_, _12797_);
  or (_31056_, _31055_, _30983_);
  and (_31057_, _31056_, _06402_);
  or (_31058_, _31057_, _31052_);
  and (_31059_, _31058_, _07132_);
  or (_31060_, _30983_, _12834_);
  and (_31061_, _31048_, _06306_);
  and (_31062_, _31061_, _31060_);
  or (_31063_, _31062_, _31059_);
  and (_31064_, _31063_, _07130_);
  and (_31066_, _30996_, _06411_);
  and (_31067_, _31066_, _31060_);
  or (_31068_, _31067_, _06303_);
  or (_31069_, _31068_, _31064_);
  and (_31070_, _30175_, _12797_);
  or (_31071_, _30983_, _08819_);
  or (_31072_, _31071_, _31070_);
  and (_31073_, _31072_, _08824_);
  and (_31074_, _31073_, _31069_);
  and (_31075_, _30185_, _12797_);
  or (_31077_, _31075_, _30983_);
  and (_31078_, _31077_, _06396_);
  or (_31079_, _31078_, _06433_);
  or (_31080_, _31079_, _31074_);
  or (_31081_, _30993_, _06829_);
  and (_31082_, _31081_, _05749_);
  and (_31083_, _31082_, _31080_);
  and (_31084_, _30990_, _05748_);
  or (_31085_, _31084_, _06440_);
  or (_31086_, _31085_, _31083_);
  and (_31088_, _30219_, _12797_);
  or (_31089_, _30983_, _06444_);
  or (_31090_, _31089_, _31088_);
  and (_31091_, _31090_, _01317_);
  and (_31092_, _31091_, _31086_);
  nor (_31093_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_31094_, _31093_, _00000_);
  or (_43716_, _31094_, _31092_);
  nor (_31095_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_31096_, _31095_, _00000_);
  and (_31098_, _12991_, \oc8051_golden_model_1.P3 [4]);
  and (_31099_, _12797_, _08336_);
  or (_31100_, _31099_, _31098_);
  or (_31101_, _31100_, _06132_);
  and (_31102_, _12996_, \oc8051_golden_model_1.P3 [4]);
  and (_31103_, _30242_, _12780_);
  or (_31104_, _31103_, _31102_);
  and (_31105_, _31104_, _06152_);
  and (_31106_, _30248_, _12797_);
  or (_31107_, _31106_, _31098_);
  or (_31109_, _31107_, _06161_);
  and (_31110_, _12797_, \oc8051_golden_model_1.ACC [4]);
  or (_31111_, _31110_, _31098_);
  and (_31112_, _31111_, _07056_);
  and (_31113_, _07057_, \oc8051_golden_model_1.P3 [4]);
  or (_31114_, _31113_, _06160_);
  or (_31115_, _31114_, _31112_);
  and (_31116_, _31115_, _06157_);
  and (_31117_, _31116_, _31109_);
  and (_31118_, _30261_, _12780_);
  or (_31120_, _31118_, _31102_);
  and (_31121_, _31120_, _06156_);
  or (_31122_, _31121_, _06217_);
  or (_31123_, _31122_, _31117_);
  or (_31124_, _31100_, _07075_);
  and (_31125_, _31124_, _31123_);
  or (_31126_, _31125_, _06220_);
  or (_31127_, _31111_, _06229_);
  and (_31128_, _31127_, _06153_);
  and (_31129_, _31128_, _31126_);
  or (_31131_, _31129_, _31105_);
  and (_31132_, _31131_, _06146_);
  or (_31133_, _31102_, _30276_);
  and (_31134_, _31120_, _06145_);
  and (_31135_, _31134_, _31133_);
  or (_31136_, _31135_, _31132_);
  and (_31137_, _31136_, _06140_);
  and (_31138_, _30283_, _12780_);
  or (_31139_, _31138_, _31102_);
  and (_31140_, _31139_, _06139_);
  or (_31143_, _31140_, _09842_);
  or (_31144_, _31143_, _31137_);
  and (_31145_, _31144_, _31101_);
  or (_31146_, _31145_, _06116_);
  and (_31147_, _12797_, _09209_);
  or (_31148_, _31098_, _06117_);
  or (_31149_, _31148_, _31147_);
  and (_31150_, _31149_, _06114_);
  and (_31151_, _31150_, _31146_);
  and (_31152_, _30305_, _12797_);
  or (_31154_, _31152_, _31098_);
  and (_31155_, _31154_, _05787_);
  or (_31156_, _31155_, _06110_);
  or (_31157_, _31156_, _31151_);
  and (_31158_, _12797_, _08715_);
  or (_31159_, _31158_, _31098_);
  or (_31160_, _31159_, _06111_);
  and (_31161_, _31160_, _07127_);
  and (_31162_, _31161_, _31157_);
  and (_31163_, _30317_, _12797_);
  or (_31166_, _31163_, _31098_);
  or (_31167_, _31098_, _30320_);
  and (_31168_, _31167_, _06297_);
  and (_31169_, _31168_, _31166_);
  or (_31170_, _31169_, _06402_);
  or (_31171_, _31170_, _31162_);
  and (_31172_, _30330_, _30327_);
  and (_31173_, _31172_, _12797_);
  or (_31174_, _31098_, _07125_);
  or (_31175_, _31174_, _31173_);
  and (_31177_, _31175_, _07132_);
  and (_31178_, _31177_, _31171_);
  or (_31179_, _31098_, _12826_);
  and (_31180_, _31159_, _06306_);
  and (_31181_, _31180_, _31179_);
  or (_31182_, _31181_, _31178_);
  and (_31183_, _31182_, _07130_);
  and (_31184_, _31111_, _06411_);
  and (_31185_, _31184_, _31179_);
  or (_31186_, _31185_, _06303_);
  or (_31189_, _31186_, _31183_);
  or (_31190_, _31166_, _08819_);
  and (_31191_, _31190_, _08824_);
  and (_31192_, _31191_, _31189_);
  and (_31193_, _30327_, _12797_);
  or (_31194_, _31193_, _31098_);
  and (_31195_, _31194_, _06396_);
  or (_31196_, _31195_, _06433_);
  or (_31197_, _31196_, _31192_);
  or (_31198_, _31107_, _06829_);
  and (_31200_, _31198_, _05749_);
  and (_31201_, _31200_, _31197_);
  and (_31202_, _31104_, _05748_);
  or (_31203_, _31202_, _06440_);
  or (_31204_, _31203_, _31201_);
  and (_31205_, _30361_, _12797_);
  or (_31206_, _31098_, _06444_);
  or (_31207_, _31206_, _31205_);
  and (_31208_, _31207_, _01317_);
  and (_31209_, _31208_, _31204_);
  or (_43717_, _31209_, _31096_);
  and (_31212_, _12991_, \oc8051_golden_model_1.P3 [5]);
  and (_31213_, _12797_, _08101_);
  or (_31214_, _31213_, _31212_);
  or (_31215_, _31214_, _06132_);
  and (_31216_, _30378_, _12797_);
  or (_31217_, _31216_, _31212_);
  or (_31218_, _31217_, _06161_);
  and (_31219_, _12797_, \oc8051_golden_model_1.ACC [5]);
  or (_31220_, _31219_, _31212_);
  and (_31222_, _31220_, _07056_);
  and (_31223_, _07057_, \oc8051_golden_model_1.P3 [5]);
  or (_31224_, _31223_, _06160_);
  or (_31225_, _31224_, _31222_);
  and (_31226_, _31225_, _06157_);
  and (_31227_, _31226_, _31218_);
  and (_31228_, _12996_, \oc8051_golden_model_1.P3 [5]);
  and (_31229_, _30400_, _12780_);
  or (_31230_, _31229_, _31228_);
  and (_31231_, _31230_, _06156_);
  or (_31233_, _31231_, _06217_);
  or (_31234_, _31233_, _31227_);
  or (_31235_, _31214_, _07075_);
  and (_31236_, _31235_, _31234_);
  or (_31237_, _31236_, _06220_);
  or (_31238_, _31220_, _06229_);
  and (_31239_, _31238_, _06153_);
  and (_31240_, _31239_, _31237_);
  and (_31241_, _30414_, _12780_);
  or (_31242_, _31241_, _31228_);
  and (_31244_, _31242_, _06152_);
  or (_31245_, _31244_, _06145_);
  or (_31246_, _31245_, _31240_);
  or (_31247_, _31228_, _30420_);
  and (_31248_, _31247_, _31230_);
  or (_31249_, _31248_, _06146_);
  and (_31250_, _31249_, _06140_);
  and (_31251_, _31250_, _31246_);
  and (_31252_, _30426_, _12780_);
  or (_31253_, _31252_, _31228_);
  and (_31254_, _31253_, _06139_);
  or (_31255_, _31254_, _09842_);
  or (_31256_, _31255_, _31251_);
  and (_31257_, _31256_, _31215_);
  or (_31258_, _31257_, _06116_);
  and (_31259_, _12797_, _09208_);
  or (_31260_, _31212_, _06117_);
  or (_31261_, _31260_, _31259_);
  and (_31262_, _31261_, _06114_);
  and (_31263_, _31262_, _31258_);
  and (_31266_, _30449_, _12797_);
  or (_31267_, _31266_, _31212_);
  and (_31268_, _31267_, _05787_);
  or (_31269_, _31268_, _06110_);
  or (_31270_, _31269_, _31263_);
  and (_31271_, _12797_, _08736_);
  or (_31272_, _31271_, _31212_);
  or (_31273_, _31272_, _06111_);
  and (_31274_, _31273_, _07127_);
  and (_31275_, _31274_, _31270_);
  and (_31276_, _30461_, _12797_);
  or (_31277_, _31276_, _31212_);
  or (_31278_, _31212_, _30464_);
  and (_31279_, _31278_, _06297_);
  and (_31280_, _31279_, _31277_);
  or (_31281_, _31280_, _31275_);
  and (_31282_, _31281_, _07125_);
  and (_31283_, _30471_, _12797_);
  or (_31284_, _31283_, _31212_);
  or (_31285_, _31212_, _30474_);
  and (_31288_, _31285_, _06402_);
  and (_31289_, _31288_, _31284_);
  or (_31290_, _31289_, _31282_);
  and (_31291_, _31290_, _07132_);
  or (_31292_, _31212_, _12818_);
  and (_31293_, _31272_, _06306_);
  and (_31294_, _31293_, _31292_);
  or (_31295_, _31294_, _31291_);
  and (_31296_, _31295_, _07130_);
  and (_31297_, _31220_, _06411_);
  and (_31298_, _31297_, _31292_);
  or (_31299_, _31298_, _06303_);
  or (_31300_, _31299_, _31296_);
  or (_31301_, _31277_, _08819_);
  and (_31302_, _31301_, _08824_);
  and (_31303_, _31302_, _31300_);
  and (_31304_, _31284_, _06396_);
  or (_31305_, _31304_, _06433_);
  or (_31306_, _31305_, _31303_);
  or (_31307_, _31217_, _06829_);
  and (_31310_, _31307_, _05749_);
  and (_31311_, _31310_, _31306_);
  and (_31312_, _31242_, _05748_);
  or (_31313_, _31312_, _06440_);
  or (_31314_, _31313_, _31311_);
  and (_31315_, _30505_, _12797_);
  or (_31316_, _31212_, _06444_);
  or (_31317_, _31316_, _31315_);
  and (_31318_, _31317_, _01317_);
  and (_31319_, _31318_, _31314_);
  nor (_31320_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_31321_, _31320_, _00000_);
  or (_43719_, _31321_, _31319_);
  and (_31322_, _12991_, \oc8051_golden_model_1.P3 [6]);
  and (_31323_, _12797_, _08012_);
  or (_31324_, _31323_, _31322_);
  or (_31325_, _31324_, _06132_);
  and (_31326_, _12996_, \oc8051_golden_model_1.P3 [6]);
  and (_31327_, _30526_, _12780_);
  or (_31328_, _31327_, _31326_);
  and (_31331_, _31328_, _06152_);
  and (_31332_, _30532_, _12797_);
  or (_31333_, _31332_, _31322_);
  or (_31334_, _31333_, _06161_);
  and (_31335_, _12797_, \oc8051_golden_model_1.ACC [6]);
  or (_31336_, _31335_, _31322_);
  and (_31337_, _31336_, _07056_);
  and (_31338_, _07057_, \oc8051_golden_model_1.P3 [6]);
  or (_31339_, _31338_, _06160_);
  or (_31340_, _31339_, _31337_);
  and (_31341_, _31340_, _06157_);
  and (_31342_, _31341_, _31334_);
  and (_31343_, _30545_, _12780_);
  or (_31344_, _31343_, _31326_);
  and (_31345_, _31344_, _06156_);
  or (_31346_, _31345_, _06217_);
  or (_31347_, _31346_, _31342_);
  or (_31348_, _31324_, _07075_);
  and (_31349_, _31348_, _31347_);
  or (_31350_, _31349_, _06220_);
  or (_31353_, _31336_, _06229_);
  and (_31354_, _31353_, _06153_);
  and (_31355_, _31354_, _31350_);
  or (_31356_, _31355_, _31331_);
  and (_31357_, _31356_, _06146_);
  or (_31358_, _31326_, _30560_);
  and (_31359_, _31344_, _06145_);
  and (_31360_, _31359_, _31358_);
  or (_31361_, _31360_, _31357_);
  and (_31362_, _31361_, _06140_);
  and (_31363_, _30567_, _12780_);
  or (_31364_, _31363_, _31326_);
  and (_31365_, _31364_, _06139_);
  or (_31366_, _31365_, _09842_);
  or (_31367_, _31366_, _31362_);
  and (_31368_, _31367_, _31325_);
  or (_31369_, _31368_, _06116_);
  and (_31370_, _12797_, _09207_);
  or (_31371_, _31322_, _06117_);
  or (_31372_, _31371_, _31370_);
  and (_31375_, _31372_, _06114_);
  and (_31376_, _31375_, _31369_);
  and (_31377_, _30589_, _12797_);
  or (_31378_, _31377_, _31322_);
  and (_31379_, _31378_, _05787_);
  or (_31380_, _31379_, _06110_);
  or (_31381_, _31380_, _31376_);
  and (_31382_, _12797_, _15402_);
  or (_31383_, _31382_, _31322_);
  or (_31384_, _31383_, _06111_);
  and (_31385_, _31384_, _07127_);
  and (_31386_, _31385_, _31381_);
  and (_31387_, _30601_, _12797_);
  or (_31388_, _31387_, _31322_);
  or (_31389_, _31322_, _30604_);
  and (_31390_, _31389_, _06297_);
  and (_31391_, _31390_, _31388_);
  or (_31392_, _31391_, _06402_);
  or (_31393_, _31392_, _31386_);
  and (_31394_, _30613_, _12797_);
  or (_31396_, _31322_, _07125_);
  or (_31397_, _31396_, _31394_);
  and (_31398_, _31397_, _07132_);
  and (_31399_, _31398_, _31393_);
  or (_31400_, _31322_, _12810_);
  and (_31401_, _31383_, _06306_);
  and (_31402_, _31401_, _31400_);
  or (_31403_, _31402_, _31399_);
  and (_31404_, _31403_, _07130_);
  and (_31405_, _31336_, _06411_);
  and (_31406_, _31405_, _31400_);
  or (_31407_, _31406_, _06303_);
  or (_31408_, _31407_, _31404_);
  or (_31409_, _31388_, _08819_);
  and (_31410_, _31409_, _08824_);
  and (_31411_, _31410_, _31408_);
  and (_31412_, _30611_, _12797_);
  or (_31413_, _31412_, _31322_);
  and (_31414_, _31413_, _06396_);
  or (_31415_, _31414_, _06433_);
  or (_31418_, _31415_, _31411_);
  or (_31419_, _31333_, _06829_);
  and (_31420_, _31419_, _05749_);
  and (_31421_, _31420_, _31418_);
  and (_31422_, _31328_, _05748_);
  or (_31423_, _31422_, _06440_);
  or (_31424_, _31423_, _31421_);
  and (_31425_, _30646_, _12797_);
  or (_31426_, _31322_, _06444_);
  or (_31427_, _31426_, _31425_);
  and (_31428_, _31427_, _01317_);
  and (_31429_, _31428_, _31424_);
  nor (_31430_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_31431_, _31430_, _00000_);
  or (_43720_, _31431_, _31429_);
  nor (_31432_, \oc8051_golden_model_1.P0 [0], rst);
  nor (_31433_, _31432_, _00000_);
  and (_31434_, _13096_, \oc8051_golden_model_1.P0 [0]);
  and (_31435_, _29675_, _12789_);
  or (_31436_, _31435_, _31434_);
  and (_31439_, _31436_, _06402_);
  and (_31440_, _12789_, _07049_);
  or (_31441_, _31440_, _31434_);
  or (_31442_, _31441_, _06132_);
  and (_31443_, _13101_, \oc8051_golden_model_1.P0 [0]);
  and (_31444_, _29705_, _07847_);
  or (_31445_, _31444_, _31443_);
  or (_31446_, _31445_, _06157_);
  nor (_31447_, _12858_, _13096_);
  or (_31448_, _31447_, _31434_);
  and (_31449_, _31448_, _06160_);
  and (_31450_, _07057_, \oc8051_golden_model_1.P0 [0]);
  and (_31451_, _12789_, \oc8051_golden_model_1.ACC [0]);
  or (_31452_, _31451_, _31434_);
  and (_31453_, _31452_, _07056_);
  or (_31454_, _31453_, _31450_);
  and (_31455_, _31454_, _06161_);
  or (_31456_, _31455_, _06156_);
  or (_31457_, _31456_, _31449_);
  and (_31458_, _31457_, _31446_);
  and (_31461_, _31458_, _07075_);
  and (_31462_, _31441_, _06217_);
  or (_31463_, _31462_, _06220_);
  or (_31464_, _31463_, _31461_);
  or (_31465_, _31452_, _06229_);
  and (_31466_, _31465_, _06153_);
  and (_31467_, _31466_, _31464_);
  and (_31468_, _31434_, _06152_);
  or (_31469_, _31468_, _06145_);
  or (_31470_, _31469_, _31467_);
  or (_31471_, _31448_, _06146_);
  and (_31472_, _31471_, _06140_);
  and (_31473_, _31472_, _31470_);
  or (_31474_, _31443_, _14170_);
  and (_31475_, _31474_, _06139_);
  and (_31476_, _31475_, _31445_);
  or (_31477_, _31476_, _09842_);
  or (_31478_, _31477_, _31473_);
  and (_31479_, _31478_, _31442_);
  or (_31480_, _31479_, _06116_);
  and (_31483_, _12789_, _09160_);
  or (_31484_, _31434_, _06117_);
  or (_31485_, _31484_, _31483_);
  and (_31486_, _31485_, _06114_);
  and (_31487_, _31486_, _31480_);
  and (_31488_, _29746_, _12789_);
  or (_31489_, _31488_, _31434_);
  and (_31490_, _31489_, _05787_);
  or (_31491_, _31490_, _31487_);
  or (_31492_, _31491_, _11136_);
  and (_31493_, _29756_, _12789_);
  or (_31494_, _31434_, _07127_);
  or (_31495_, _31494_, _31493_);
  and (_31496_, _12789_, _08708_);
  or (_31497_, _31496_, _31434_);
  or (_31498_, _31497_, _06111_);
  and (_31499_, _31498_, _07125_);
  and (_31500_, _31499_, _31495_);
  and (_31501_, _31500_, _31492_);
  or (_31502_, _31501_, _31439_);
  and (_31505_, _31502_, _07132_);
  nand (_31506_, _31497_, _06306_);
  nor (_31507_, _31506_, _31447_);
  or (_31508_, _31507_, _31505_);
  and (_31509_, _31508_, _07130_);
  or (_31510_, _31434_, _12858_);
  and (_31511_, _31452_, _06411_);
  and (_31512_, _31511_, _31510_);
  or (_31513_, _31512_, _06303_);
  or (_31514_, _31513_, _31509_);
  and (_31515_, _29752_, _12789_);
  or (_31516_, _31434_, _08819_);
  or (_31517_, _31516_, _31515_);
  and (_31518_, _31517_, _08824_);
  and (_31519_, _31518_, _31514_);
  and (_31520_, _29673_, _12789_);
  or (_31521_, _31520_, _31434_);
  and (_31522_, _31521_, _06396_);
  or (_31523_, _31522_, _06433_);
  or (_31524_, _31523_, _31519_);
  or (_31527_, _31448_, _06829_);
  and (_31528_, _31527_, _05749_);
  and (_31529_, _31528_, _31524_);
  and (_31530_, _31434_, _05748_);
  or (_31531_, _31530_, _06440_);
  or (_31532_, _31531_, _31529_);
  or (_31533_, _31448_, _06444_);
  and (_31534_, _31533_, _01317_);
  and (_31535_, _31534_, _31532_);
  or (_43721_, _31535_, _31433_);
  nor (_31536_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_31537_, _31536_, _00000_);
  or (_31538_, _29883_, _13096_);
  or (_31539_, _12789_, \oc8051_golden_model_1.P0 [1]);
  and (_31540_, _31539_, _05787_);
  and (_31541_, _31540_, _31538_);
  and (_31542_, _29814_, _07847_);
  and (_31543_, _31542_, _29813_);
  and (_31544_, _13101_, \oc8051_golden_model_1.P0 [1]);
  or (_31545_, _31544_, _06146_);
  or (_31548_, _31545_, _31543_);
  and (_31549_, _29823_, _12789_);
  not (_31550_, _31549_);
  and (_31551_, _31550_, _31539_);
  or (_31552_, _31551_, _06161_);
  nand (_31553_, _12789_, _05887_);
  and (_31554_, _31553_, _31539_);
  and (_31555_, _31554_, _07056_);
  and (_31556_, _07057_, \oc8051_golden_model_1.P0 [1]);
  or (_31557_, _31556_, _06160_);
  or (_31558_, _31557_, _31555_);
  and (_31559_, _31558_, _06157_);
  and (_31560_, _31559_, _31552_);
  or (_31561_, _31544_, _06217_);
  or (_31562_, _31561_, _31542_);
  and (_31563_, _31562_, _13860_);
  or (_31564_, _31563_, _31560_);
  and (_31565_, _13096_, \oc8051_golden_model_1.P0 [1]);
  and (_31566_, _12789_, _07306_);
  or (_31567_, _31566_, _31565_);
  or (_31570_, _31567_, _07075_);
  and (_31571_, _31570_, _31564_);
  or (_31572_, _31571_, _06220_);
  or (_31573_, _31554_, _06229_);
  and (_31574_, _31573_, _06153_);
  and (_31575_, _31574_, _31572_);
  and (_31576_, _29851_, _07847_);
  or (_31577_, _31576_, _31544_);
  and (_31578_, _31577_, _06152_);
  or (_31579_, _31578_, _06145_);
  or (_31580_, _31579_, _31575_);
  and (_31581_, _31580_, _31548_);
  and (_31582_, _31581_, _06140_);
  and (_31583_, _29860_, _07847_);
  or (_31584_, _31544_, _31583_);
  and (_31585_, _31584_, _06139_);
  or (_31586_, _31585_, _09842_);
  or (_31587_, _31586_, _31582_);
  or (_31588_, _31567_, _06132_);
  and (_31589_, _31588_, _31587_);
  or (_31592_, _31589_, _06116_);
  and (_31593_, _12789_, _09115_);
  or (_31594_, _31565_, _06117_);
  or (_31595_, _31594_, _31593_);
  and (_31596_, _31595_, _06114_);
  and (_31597_, _31596_, _31592_);
  or (_31598_, _31597_, _31541_);
  and (_31599_, _31598_, _06298_);
  or (_31600_, _30823_, _13096_);
  and (_31601_, _31600_, _06297_);
  nand (_31602_, _12789_, _06945_);
  and (_31603_, _31602_, _06110_);
  or (_31604_, _31603_, _31601_);
  and (_31605_, _31604_, _31539_);
  or (_31606_, _31605_, _31599_);
  and (_31607_, _31606_, _07125_);
  or (_31608_, _30833_, _13096_);
  and (_31609_, _31539_, _06402_);
  and (_31610_, _31609_, _31608_);
  or (_31611_, _31610_, _31607_);
  and (_31614_, _31611_, _07132_);
  or (_31615_, _29896_, _13096_);
  and (_31616_, _31539_, _06306_);
  and (_31617_, _31616_, _31615_);
  or (_31618_, _31617_, _31614_);
  and (_31619_, _31618_, _07130_);
  or (_31620_, _31565_, _12850_);
  and (_31621_, _31554_, _06411_);
  and (_31622_, _31621_, _31620_);
  or (_31623_, _31622_, _31619_);
  and (_31624_, _31623_, _06397_);
  or (_31625_, _31602_, _12850_);
  and (_31626_, _31539_, _06303_);
  and (_31627_, _31626_, _31625_);
  or (_31628_, _31553_, _12850_);
  and (_31629_, _31539_, _06396_);
  and (_31630_, _31629_, _31628_);
  or (_31631_, _31630_, _06433_);
  or (_31632_, _31631_, _31627_);
  or (_31633_, _31632_, _31624_);
  or (_31636_, _31551_, _06829_);
  and (_31637_, _31636_, _05749_);
  and (_31638_, _31637_, _31633_);
  and (_31639_, _31577_, _05748_);
  or (_31640_, _31639_, _06440_);
  or (_31641_, _31640_, _31638_);
  or (_31642_, _31565_, _06444_);
  or (_31643_, _31642_, _31549_);
  and (_31644_, _31643_, _01317_);
  and (_31645_, _31644_, _31641_);
  or (_43723_, _31645_, _31537_);
  nor (_31646_, \oc8051_golden_model_1.P0 [2], rst);
  nor (_31647_, _31646_, _00000_);
  and (_31648_, _13096_, \oc8051_golden_model_1.P0 [2]);
  and (_31649_, _12789_, _07708_);
  or (_31650_, _31649_, _31648_);
  or (_31651_, _31650_, _06132_);
  and (_31652_, _29954_, _12789_);
  or (_31653_, _31652_, _31648_);
  or (_31654_, _31653_, _06161_);
  and (_31657_, _12789_, \oc8051_golden_model_1.ACC [2]);
  or (_31658_, _31657_, _31648_);
  and (_31659_, _31658_, _07056_);
  and (_31660_, _07057_, \oc8051_golden_model_1.P0 [2]);
  or (_31661_, _31660_, _06160_);
  or (_31662_, _31661_, _31659_);
  and (_31663_, _31662_, _06157_);
  and (_31664_, _31663_, _31654_);
  and (_31665_, _13101_, \oc8051_golden_model_1.P0 [2]);
  and (_31666_, _29976_, _07847_);
  or (_31667_, _31666_, _31665_);
  and (_31668_, _31667_, _06156_);
  or (_31669_, _31668_, _06217_);
  or (_31670_, _31669_, _31664_);
  or (_31671_, _31650_, _07075_);
  and (_31672_, _31671_, _31670_);
  or (_31673_, _31672_, _06220_);
  or (_31674_, _31658_, _06229_);
  and (_31675_, _31674_, _06153_);
  and (_31676_, _31675_, _31673_);
  and (_31679_, _29992_, _07847_);
  or (_31680_, _31679_, _31665_);
  and (_31681_, _31680_, _06152_);
  or (_31682_, _31681_, _06145_);
  or (_31683_, _31682_, _31676_);
  or (_31684_, _31665_, _29999_);
  and (_31685_, _31684_, _31667_);
  or (_31686_, _31685_, _06146_);
  and (_31687_, _31686_, _06140_);
  and (_31688_, _31687_, _31683_);
  and (_31689_, _30005_, _07847_);
  or (_31690_, _31689_, _31665_);
  and (_31691_, _31690_, _06139_);
  or (_31692_, _31691_, _09842_);
  or (_31693_, _31692_, _31688_);
  and (_31694_, _31693_, _31651_);
  or (_31695_, _31694_, _06116_);
  and (_31696_, _12789_, _09211_);
  or (_31697_, _31648_, _06117_);
  or (_31698_, _31697_, _31696_);
  and (_31701_, _31698_, _06114_);
  and (_31702_, _31701_, _31695_);
  and (_31703_, _30029_, _12789_);
  or (_31704_, _31648_, _31703_);
  and (_31705_, _31704_, _05787_);
  or (_31706_, _31705_, _31702_);
  or (_31707_, _31706_, _11136_);
  and (_31708_, _29948_, _29945_);
  and (_31709_, _31708_, _12789_);
  or (_31710_, _31648_, _07127_);
  or (_31711_, _31710_, _31709_);
  and (_31712_, _12789_, _08768_);
  or (_31713_, _31712_, _31648_);
  or (_31714_, _31713_, _06111_);
  and (_31715_, _31714_, _07125_);
  and (_31716_, _31715_, _31711_);
  and (_31717_, _31716_, _31707_);
  and (_31718_, _30043_, _12789_);
  and (_31719_, _31718_, _30046_);
  or (_31720_, _31719_, _31648_);
  and (_31723_, _31720_, _06402_);
  or (_31724_, _31723_, _31717_);
  and (_31725_, _31724_, _07132_);
  or (_31726_, _31648_, _12842_);
  and (_31727_, _31713_, _06306_);
  and (_31728_, _31727_, _31726_);
  or (_31729_, _31728_, _31725_);
  and (_31730_, _31729_, _07130_);
  and (_31731_, _31658_, _06411_);
  and (_31732_, _31731_, _31726_);
  or (_31733_, _31732_, _06303_);
  or (_31734_, _31733_, _31730_);
  and (_31735_, _29945_, _12789_);
  or (_31736_, _31648_, _08819_);
  or (_31737_, _31736_, _31735_);
  and (_31738_, _31737_, _08824_);
  and (_31739_, _31738_, _31734_);
  or (_31740_, _31718_, _31648_);
  and (_31741_, _31740_, _06396_);
  or (_31742_, _31741_, _06433_);
  or (_31745_, _31742_, _31739_);
  or (_31746_, _31653_, _06829_);
  and (_31747_, _31746_, _05749_);
  and (_31748_, _31747_, _31745_);
  and (_31749_, _31680_, _05748_);
  or (_31750_, _31749_, _06440_);
  or (_31751_, _31750_, _31748_);
  and (_31752_, _30077_, _12789_);
  or (_31753_, _31648_, _06444_);
  or (_31754_, _31753_, _31752_);
  and (_31755_, _31754_, _01317_);
  and (_31756_, _31755_, _31751_);
  or (_43724_, _31756_, _31647_);
  and (_31757_, _13096_, \oc8051_golden_model_1.P0 [3]);
  and (_31758_, _12789_, _07544_);
  or (_31759_, _31758_, _31757_);
  or (_31760_, _31759_, _06132_);
  and (_31761_, _13101_, \oc8051_golden_model_1.P0 [3]);
  and (_31762_, _30100_, _07847_);
  or (_31763_, _31762_, _31761_);
  and (_31766_, _31763_, _06152_);
  and (_31767_, _30106_, _12789_);
  or (_31768_, _31767_, _31757_);
  or (_31769_, _31768_, _06161_);
  and (_31770_, _12789_, \oc8051_golden_model_1.ACC [3]);
  or (_31771_, _31770_, _31757_);
  and (_31772_, _31771_, _07056_);
  and (_31773_, _07057_, \oc8051_golden_model_1.P0 [3]);
  or (_31774_, _31773_, _06160_);
  or (_31775_, _31774_, _31772_);
  and (_31776_, _31775_, _06157_);
  and (_31777_, _31776_, _31769_);
  and (_31778_, _30119_, _07847_);
  or (_31779_, _31778_, _31761_);
  and (_31780_, _31779_, _06156_);
  or (_31781_, _31780_, _06217_);
  or (_31782_, _31781_, _31777_);
  or (_31783_, _31759_, _07075_);
  and (_31784_, _31783_, _31782_);
  or (_31785_, _31784_, _06220_);
  or (_31788_, _31771_, _06229_);
  and (_31789_, _31788_, _06153_);
  and (_31790_, _31789_, _31785_);
  or (_31791_, _31790_, _31766_);
  and (_31792_, _31791_, _06146_);
  or (_31793_, _31761_, _30134_);
  and (_31794_, _31779_, _06145_);
  and (_31795_, _31794_, _31793_);
  or (_31796_, _31795_, _31792_);
  and (_31797_, _31796_, _06140_);
  and (_31798_, _30141_, _07847_);
  or (_31799_, _31798_, _31761_);
  and (_31800_, _31799_, _06139_);
  or (_31801_, _31800_, _09842_);
  or (_31802_, _31801_, _31797_);
  and (_31803_, _31802_, _31760_);
  or (_31804_, _31803_, _06116_);
  and (_31805_, _12789_, _09210_);
  or (_31806_, _31757_, _06117_);
  or (_31807_, _31806_, _31805_);
  and (_31810_, _31807_, _06114_);
  and (_31811_, _31810_, _31804_);
  and (_31812_, _30163_, _12789_);
  or (_31813_, _31812_, _31757_);
  and (_31814_, _31813_, _05787_);
  or (_31815_, _31814_, _11136_);
  or (_31816_, _31815_, _31811_);
  and (_31817_, _31042_, _12789_);
  or (_31818_, _31757_, _07127_);
  or (_31819_, _31818_, _31817_);
  and (_31820_, _12789_, _08712_);
  or (_31821_, _31820_, _31757_);
  or (_31822_, _31821_, _06111_);
  and (_31823_, _31822_, _07125_);
  and (_31824_, _31823_, _31819_);
  and (_31825_, _31824_, _31816_);
  and (_31826_, _31053_, _12789_);
  or (_31827_, _31826_, _31757_);
  and (_31828_, _31827_, _06402_);
  or (_31829_, _31828_, _31825_);
  and (_31832_, _31829_, _07132_);
  or (_31833_, _31757_, _12834_);
  and (_31834_, _31821_, _06306_);
  and (_31835_, _31834_, _31833_);
  or (_31836_, _31835_, _31832_);
  and (_31837_, _31836_, _07130_);
  and (_31838_, _31771_, _06411_);
  and (_31839_, _31838_, _31833_);
  or (_31840_, _31839_, _06303_);
  or (_31841_, _31840_, _31837_);
  and (_31842_, _30175_, _12789_);
  or (_31843_, _31757_, _08819_);
  or (_31844_, _31843_, _31842_);
  and (_31845_, _31844_, _08824_);
  and (_31846_, _31845_, _31841_);
  and (_31847_, _30185_, _12789_);
  or (_31848_, _31847_, _31757_);
  and (_31849_, _31848_, _06396_);
  or (_31850_, _31849_, _06433_);
  or (_31851_, _31850_, _31846_);
  or (_31854_, _31768_, _06829_);
  and (_31855_, _31854_, _05749_);
  and (_31856_, _31855_, _31851_);
  and (_31857_, _31763_, _05748_);
  or (_31858_, _31857_, _06440_);
  or (_31859_, _31858_, _31856_);
  and (_31860_, _30219_, _12789_);
  or (_31861_, _31757_, _06444_);
  or (_31862_, _31861_, _31860_);
  and (_31863_, _31862_, _01317_);
  and (_31865_, _31863_, _31859_);
  nor (_31866_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_31867_, _31866_, _00000_);
  or (_43725_, _31867_, _31865_);
  and (_31868_, _13096_, \oc8051_golden_model_1.P0 [4]);
  and (_31869_, _12789_, _08336_);
  or (_31870_, _31869_, _31868_);
  or (_31871_, _31870_, _06132_);
  and (_31872_, _13101_, \oc8051_golden_model_1.P0 [4]);
  and (_31873_, _30242_, _07847_);
  or (_31875_, _31873_, _31872_);
  and (_31876_, _31875_, _06152_);
  and (_31877_, _30248_, _12789_);
  or (_31878_, _31877_, _31868_);
  or (_31879_, _31878_, _06161_);
  and (_31880_, _12789_, \oc8051_golden_model_1.ACC [4]);
  or (_31881_, _31880_, _31868_);
  and (_31882_, _31881_, _07056_);
  and (_31883_, _07057_, \oc8051_golden_model_1.P0 [4]);
  or (_31884_, _31883_, _06160_);
  or (_31886_, _31884_, _31882_);
  and (_31887_, _31886_, _06157_);
  and (_31888_, _31887_, _31879_);
  and (_31889_, _30261_, _07847_);
  or (_31890_, _31889_, _31872_);
  and (_31891_, _31890_, _06156_);
  or (_31892_, _31891_, _06217_);
  or (_31893_, _31892_, _31888_);
  or (_31894_, _31870_, _07075_);
  and (_31895_, _31894_, _31893_);
  or (_31897_, _31895_, _06220_);
  or (_31898_, _31881_, _06229_);
  and (_31899_, _31898_, _06153_);
  and (_31900_, _31899_, _31897_);
  or (_31901_, _31900_, _31876_);
  and (_31902_, _31901_, _06146_);
  or (_31903_, _31872_, _30276_);
  and (_31904_, _31890_, _06145_);
  and (_31905_, _31904_, _31903_);
  or (_31906_, _31905_, _31902_);
  and (_31908_, _31906_, _06140_);
  and (_31909_, _30283_, _07847_);
  or (_31910_, _31909_, _31872_);
  and (_31911_, _31910_, _06139_);
  or (_31912_, _31911_, _09842_);
  or (_31913_, _31912_, _31908_);
  and (_31914_, _31913_, _31871_);
  or (_31915_, _31914_, _06116_);
  and (_31916_, _12789_, _09209_);
  or (_31917_, _31868_, _06117_);
  or (_31919_, _31917_, _31916_);
  and (_31920_, _31919_, _06114_);
  and (_31921_, _31920_, _31915_);
  and (_31922_, _30305_, _12789_);
  or (_31923_, _31922_, _31868_);
  and (_31924_, _31923_, _05787_);
  or (_31925_, _31924_, _11136_);
  or (_31926_, _31925_, _31921_);
  and (_31927_, _30317_, _12789_);
  and (_31928_, _31927_, _30320_);
  or (_31930_, _31868_, _07127_);
  or (_31931_, _31930_, _31928_);
  and (_31932_, _12789_, _08715_);
  or (_31933_, _31932_, _31868_);
  or (_31934_, _31933_, _06111_);
  and (_31935_, _31934_, _07125_);
  and (_31936_, _31935_, _31931_);
  and (_31937_, _31936_, _31926_);
  and (_31938_, _31172_, _12789_);
  or (_31939_, _31938_, _31868_);
  and (_31941_, _31939_, _06402_);
  or (_31942_, _31941_, _31937_);
  and (_31943_, _31942_, _07132_);
  or (_31944_, _31868_, _12826_);
  and (_31945_, _31933_, _06306_);
  and (_31946_, _31945_, _31944_);
  or (_31947_, _31946_, _31943_);
  and (_31948_, _31947_, _07130_);
  and (_31949_, _31881_, _06411_);
  and (_31950_, _31949_, _31944_);
  or (_31951_, _31950_, _06303_);
  or (_31952_, _31951_, _31948_);
  or (_31953_, _31868_, _08819_);
  or (_31954_, _31953_, _31927_);
  and (_31955_, _31954_, _08824_);
  and (_31956_, _31955_, _31952_);
  and (_31957_, _30327_, _12789_);
  or (_31958_, _31957_, _31868_);
  and (_31959_, _31958_, _06396_);
  or (_31960_, _31959_, _06433_);
  or (_31962_, _31960_, _31956_);
  or (_31963_, _31878_, _06829_);
  and (_31964_, _31963_, _05749_);
  and (_31965_, _31964_, _31962_);
  and (_31966_, _31875_, _05748_);
  or (_31967_, _31966_, _06440_);
  or (_31968_, _31967_, _31965_);
  and (_31969_, _30361_, _12789_);
  or (_31970_, _31868_, _06444_);
  or (_31971_, _31970_, _31969_);
  and (_31973_, _31971_, _01317_);
  and (_31974_, _31973_, _31968_);
  nor (_31975_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_31976_, _31975_, _00000_);
  or (_43726_, _31976_, _31974_);
  and (_31977_, _13096_, \oc8051_golden_model_1.P0 [5]);
  and (_31978_, _12789_, _08101_);
  or (_31979_, _31978_, _31977_);
  or (_31980_, _31979_, _06132_);
  and (_31981_, _30378_, _12789_);
  or (_31983_, _31981_, _31977_);
  or (_31984_, _31983_, _06161_);
  and (_31985_, _12789_, \oc8051_golden_model_1.ACC [5]);
  or (_31986_, _31985_, _31977_);
  and (_31987_, _31986_, _07056_);
  and (_31988_, _07057_, \oc8051_golden_model_1.P0 [5]);
  or (_31989_, _31988_, _06160_);
  or (_31990_, _31989_, _31987_);
  and (_31991_, _31990_, _06157_);
  and (_31992_, _31991_, _31984_);
  and (_31994_, _13101_, \oc8051_golden_model_1.P0 [5]);
  and (_31995_, _30400_, _07847_);
  or (_31996_, _31995_, _31994_);
  and (_31997_, _31996_, _06156_);
  or (_31998_, _31997_, _06217_);
  or (_31999_, _31998_, _31992_);
  or (_32000_, _31979_, _07075_);
  and (_32001_, _32000_, _31999_);
  or (_32002_, _32001_, _06220_);
  or (_32003_, _31986_, _06229_);
  and (_32005_, _32003_, _06153_);
  and (_32006_, _32005_, _32002_);
  and (_32007_, _30414_, _07847_);
  or (_32008_, _32007_, _31994_);
  and (_32009_, _32008_, _06152_);
  or (_32010_, _32009_, _06145_);
  or (_32011_, _32010_, _32006_);
  or (_32012_, _31994_, _30420_);
  and (_32013_, _32012_, _31996_);
  or (_32014_, _32013_, _06146_);
  and (_32016_, _32014_, _06140_);
  and (_32017_, _32016_, _32011_);
  and (_32018_, _30426_, _07847_);
  or (_32019_, _32018_, _31994_);
  and (_32020_, _32019_, _06139_);
  or (_32021_, _32020_, _09842_);
  or (_32022_, _32021_, _32017_);
  and (_32023_, _32022_, _31980_);
  or (_32024_, _32023_, _06116_);
  and (_32025_, _12789_, _09208_);
  or (_32027_, _31977_, _06117_);
  or (_32028_, _32027_, _32025_);
  and (_32029_, _32028_, _06114_);
  and (_32030_, _32029_, _32024_);
  and (_32031_, _30449_, _12789_);
  or (_32032_, _32031_, _31977_);
  and (_32033_, _32032_, _05787_);
  or (_32034_, _32033_, _11136_);
  or (_32035_, _32034_, _32030_);
  and (_32036_, _30464_, _30461_);
  and (_32038_, _32036_, _12789_);
  or (_32039_, _31977_, _07127_);
  or (_32040_, _32039_, _32038_);
  and (_32041_, _12789_, _08736_);
  or (_32042_, _32041_, _31977_);
  or (_32043_, _32042_, _06111_);
  and (_32044_, _32043_, _07125_);
  and (_32045_, _32044_, _32040_);
  and (_32046_, _32045_, _32035_);
  and (_32047_, _30474_, _30471_);
  and (_32049_, _32047_, _12789_);
  or (_32050_, _32049_, _31977_);
  and (_32051_, _32050_, _06402_);
  or (_32052_, _32051_, _32046_);
  and (_32053_, _32052_, _07132_);
  or (_32054_, _31977_, _12818_);
  and (_32055_, _32042_, _06306_);
  and (_32056_, _32055_, _32054_);
  or (_32057_, _32056_, _32053_);
  and (_32058_, _32057_, _07130_);
  and (_32060_, _31986_, _06411_);
  and (_32061_, _32060_, _32054_);
  or (_32062_, _32061_, _06303_);
  or (_32063_, _32062_, _32058_);
  and (_32064_, _30461_, _12789_);
  or (_32065_, _31977_, _08819_);
  or (_32066_, _32065_, _32064_);
  and (_32067_, _32066_, _08824_);
  and (_32068_, _32067_, _32063_);
  and (_32069_, _30471_, _12789_);
  or (_32071_, _32069_, _31977_);
  and (_32072_, _32071_, _06396_);
  or (_32073_, _32072_, _06433_);
  or (_32074_, _32073_, _32068_);
  or (_32075_, _31983_, _06829_);
  and (_32076_, _32075_, _05749_);
  and (_32077_, _32076_, _32074_);
  and (_32078_, _32008_, _05748_);
  or (_32079_, _32078_, _06440_);
  or (_32080_, _32079_, _32077_);
  and (_32082_, _30505_, _12789_);
  or (_32083_, _31977_, _06444_);
  or (_32084_, _32083_, _32082_);
  and (_32085_, _32084_, _01317_);
  and (_32086_, _32085_, _32080_);
  nor (_32087_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_32088_, _32087_, _00000_);
  or (_43727_, _32088_, _32086_);
  nor (_32089_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_32090_, _32089_, _00000_);
  and (_32092_, _13096_, \oc8051_golden_model_1.P0 [6]);
  and (_32093_, _12789_, _08012_);
  or (_32094_, _32093_, _32092_);
  or (_32095_, _32094_, _06132_);
  and (_32096_, _13101_, \oc8051_golden_model_1.P0 [6]);
  and (_32097_, _30526_, _07847_);
  or (_32098_, _32097_, _32096_);
  and (_32099_, _32098_, _06152_);
  and (_32100_, _30532_, _12789_);
  or (_32101_, _32100_, _32092_);
  or (_32103_, _32101_, _06161_);
  and (_32104_, _12789_, \oc8051_golden_model_1.ACC [6]);
  or (_32105_, _32104_, _32092_);
  and (_32106_, _32105_, _07056_);
  and (_32107_, _07057_, \oc8051_golden_model_1.P0 [6]);
  or (_32108_, _32107_, _06160_);
  or (_32109_, _32108_, _32106_);
  and (_32110_, _32109_, _06157_);
  and (_32111_, _32110_, _32103_);
  and (_32112_, _30545_, _07847_);
  or (_32114_, _32112_, _32096_);
  and (_32115_, _32114_, _06156_);
  or (_32116_, _32115_, _06217_);
  or (_32117_, _32116_, _32111_);
  or (_32118_, _32094_, _07075_);
  and (_32119_, _32118_, _32117_);
  or (_32120_, _32119_, _06220_);
  or (_32121_, _32105_, _06229_);
  and (_32122_, _32121_, _06153_);
  and (_32123_, _32122_, _32120_);
  or (_32125_, _32123_, _32099_);
  and (_32126_, _32125_, _06146_);
  or (_32127_, _32096_, _30560_);
  and (_32128_, _32114_, _06145_);
  and (_32129_, _32128_, _32127_);
  or (_32130_, _32129_, _32126_);
  and (_32131_, _32130_, _06140_);
  and (_32132_, _30567_, _07847_);
  or (_32133_, _32132_, _32096_);
  and (_32134_, _32133_, _06139_);
  or (_32136_, _32134_, _09842_);
  or (_32137_, _32136_, _32131_);
  and (_32138_, _32137_, _32095_);
  or (_32139_, _32138_, _06116_);
  and (_32140_, _12789_, _09207_);
  or (_32141_, _32092_, _06117_);
  or (_32142_, _32141_, _32140_);
  and (_32143_, _32142_, _06114_);
  and (_32144_, _32143_, _32139_);
  and (_32145_, _30589_, _12789_);
  or (_32147_, _32145_, _32092_);
  and (_32148_, _32147_, _05787_);
  or (_32149_, _32148_, _11136_);
  or (_32150_, _32149_, _32144_);
  and (_32151_, _30604_, _30601_);
  and (_32152_, _32151_, _12789_);
  or (_32153_, _32092_, _07127_);
  or (_32154_, _32153_, _32152_);
  and (_32155_, _12789_, _15402_);
  or (_32156_, _32155_, _32092_);
  or (_32158_, _32156_, _06111_);
  and (_32159_, _32158_, _07125_);
  and (_32160_, _32159_, _32154_);
  and (_32161_, _32160_, _32150_);
  and (_32162_, _30613_, _12789_);
  or (_32163_, _32162_, _32092_);
  and (_32164_, _32163_, _06402_);
  or (_32165_, _32164_, _32161_);
  and (_32166_, _32165_, _07132_);
  or (_32167_, _32092_, _12810_);
  and (_32169_, _32156_, _06306_);
  and (_32170_, _32169_, _32167_);
  or (_32171_, _32170_, _32166_);
  and (_32172_, _32171_, _07130_);
  and (_32173_, _32105_, _06411_);
  and (_32174_, _32173_, _32167_);
  or (_32175_, _32174_, _06303_);
  or (_32176_, _32175_, _32172_);
  and (_32177_, _30601_, _12789_);
  or (_32178_, _32092_, _08819_);
  or (_32180_, _32178_, _32177_);
  and (_32181_, _32180_, _08824_);
  and (_32182_, _32181_, _32176_);
  and (_32183_, _30611_, _12789_);
  or (_32184_, _32183_, _32092_);
  and (_32185_, _32184_, _06396_);
  or (_32186_, _32185_, _06433_);
  or (_32187_, _32186_, _32182_);
  or (_32188_, _32101_, _06829_);
  and (_32189_, _32188_, _05749_);
  and (_32191_, _32189_, _32187_);
  and (_32192_, _32098_, _05748_);
  or (_32193_, _32192_, _06440_);
  or (_32194_, _32193_, _32191_);
  and (_32195_, _30646_, _12789_);
  or (_32196_, _32092_, _06444_);
  or (_32197_, _32196_, _32195_);
  and (_32198_, _32197_, _01317_);
  and (_32199_, _32198_, _32194_);
  or (_43728_, _32199_, _32090_);
  nor (_32201_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_32202_, _32201_, _00000_);
  and (_32203_, _13196_, \oc8051_golden_model_1.P1 [0]);
  and (_32204_, _29675_, _12792_);
  or (_32205_, _32204_, _32203_);
  and (_32206_, _32205_, _06402_);
  and (_32207_, _12792_, _07049_);
  or (_32208_, _32207_, _32203_);
  or (_32209_, _32208_, _06132_);
  and (_32210_, _13201_, \oc8051_golden_model_1.P1 [0]);
  and (_32212_, _29705_, _12778_);
  or (_32213_, _32212_, _32210_);
  or (_32214_, _32213_, _06157_);
  nor (_32215_, _12858_, _13196_);
  or (_32216_, _32215_, _32203_);
  and (_32217_, _32216_, _06160_);
  and (_32218_, _07057_, \oc8051_golden_model_1.P1 [0]);
  and (_32219_, _12792_, \oc8051_golden_model_1.ACC [0]);
  or (_32220_, _32219_, _32203_);
  and (_32221_, _32220_, _07056_);
  or (_32223_, _32221_, _32218_);
  and (_32224_, _32223_, _06161_);
  or (_32225_, _32224_, _06156_);
  or (_32226_, _32225_, _32217_);
  and (_32227_, _32226_, _32214_);
  and (_32228_, _32227_, _07075_);
  and (_32229_, _32208_, _06217_);
  or (_32230_, _32229_, _06220_);
  or (_32231_, _32230_, _32228_);
  or (_32232_, _32220_, _06229_);
  and (_32234_, _32232_, _06153_);
  and (_32235_, _32234_, _32231_);
  and (_32236_, _32203_, _06152_);
  or (_32237_, _32236_, _06145_);
  or (_32238_, _32237_, _32235_);
  or (_32239_, _32216_, _06146_);
  and (_32240_, _32239_, _06140_);
  and (_32241_, _32240_, _32238_);
  or (_32242_, _32210_, _14170_);
  and (_32243_, _32242_, _06139_);
  and (_32245_, _32243_, _32213_);
  or (_32246_, _32245_, _09842_);
  or (_32247_, _32246_, _32241_);
  and (_32248_, _32247_, _32209_);
  or (_32249_, _32248_, _06116_);
  and (_32250_, _12792_, _09160_);
  or (_32251_, _32203_, _06117_);
  or (_32252_, _32251_, _32250_);
  and (_32253_, _32252_, _06114_);
  and (_32254_, _32253_, _32249_);
  and (_32256_, _29746_, _12792_);
  or (_32257_, _32256_, _32203_);
  and (_32258_, _32257_, _05787_);
  or (_32259_, _32258_, _32254_);
  or (_32260_, _32259_, _11136_);
  and (_32261_, _29756_, _12792_);
  or (_32262_, _32203_, _07127_);
  or (_32263_, _32262_, _32261_);
  and (_32264_, _12792_, _08708_);
  or (_32265_, _32264_, _32203_);
  or (_32267_, _32265_, _06111_);
  and (_32268_, _32267_, _07125_);
  and (_32269_, _32268_, _32263_);
  and (_32270_, _32269_, _32260_);
  or (_32271_, _32270_, _32206_);
  and (_32272_, _32271_, _07132_);
  nand (_32273_, _32265_, _06306_);
  nor (_32274_, _32273_, _32215_);
  or (_32275_, _32274_, _32272_);
  and (_32276_, _32275_, _07130_);
  or (_32278_, _32203_, _12858_);
  and (_32279_, _32220_, _06411_);
  and (_32280_, _32279_, _32278_);
  or (_32281_, _32280_, _06303_);
  or (_32282_, _32281_, _32276_);
  and (_32283_, _29752_, _12792_);
  or (_32284_, _32203_, _08819_);
  or (_32285_, _32284_, _32283_);
  and (_32286_, _32285_, _08824_);
  and (_32287_, _32286_, _32282_);
  and (_32289_, _29673_, _12792_);
  or (_32290_, _32289_, _32203_);
  and (_32291_, _32290_, _06396_);
  or (_32292_, _32291_, _06433_);
  or (_32293_, _32292_, _32287_);
  or (_32294_, _32216_, _06829_);
  and (_32295_, _32294_, _05749_);
  and (_32296_, _32295_, _32293_);
  and (_32297_, _32203_, _05748_);
  or (_32298_, _32297_, _06440_);
  or (_32300_, _32298_, _32296_);
  or (_32301_, _32216_, _06444_);
  and (_32302_, _32301_, _01317_);
  and (_32303_, _32302_, _32300_);
  or (_43730_, _32303_, _32202_);
  and (_32304_, _29814_, _12778_);
  and (_32305_, _32304_, _29813_);
  and (_32306_, _13201_, \oc8051_golden_model_1.P1 [1]);
  or (_32307_, _32306_, _06146_);
  or (_32308_, _32307_, _32305_);
  or (_32310_, _12792_, \oc8051_golden_model_1.P1 [1]);
  and (_32311_, _29823_, _12792_);
  not (_32312_, _32311_);
  and (_32313_, _32312_, _32310_);
  or (_32314_, _32313_, _06161_);
  nand (_32315_, _12792_, _05887_);
  and (_32316_, _32315_, _32310_);
  and (_32317_, _32316_, _07056_);
  and (_32318_, _07057_, \oc8051_golden_model_1.P1 [1]);
  or (_32319_, _32318_, _06160_);
  or (_32321_, _32319_, _32317_);
  and (_32322_, _32321_, _06157_);
  and (_32323_, _32322_, _32314_);
  or (_32324_, _32306_, _06217_);
  or (_32325_, _32324_, _32304_);
  and (_32326_, _32325_, _13860_);
  or (_32327_, _32326_, _32323_);
  and (_32328_, _13196_, \oc8051_golden_model_1.P1 [1]);
  and (_32329_, _12792_, _07306_);
  or (_32330_, _32329_, _32328_);
  or (_32332_, _32330_, _07075_);
  and (_32333_, _32332_, _32327_);
  or (_32334_, _32333_, _06220_);
  or (_32335_, _32316_, _06229_);
  and (_32336_, _32335_, _06153_);
  and (_32337_, _32336_, _32334_);
  and (_32338_, _29851_, _12778_);
  or (_32339_, _32338_, _32306_);
  and (_32340_, _32339_, _06152_);
  or (_32341_, _32340_, _06145_);
  or (_32343_, _32341_, _32337_);
  and (_32344_, _32343_, _32308_);
  and (_32345_, _32344_, _06140_);
  and (_32346_, _29860_, _12778_);
  or (_32347_, _32306_, _32346_);
  and (_32348_, _32347_, _06139_);
  or (_32349_, _32348_, _09842_);
  or (_32350_, _32349_, _32345_);
  or (_32351_, _32330_, _06132_);
  and (_32352_, _32351_, _32350_);
  or (_32354_, _32352_, _06116_);
  and (_32355_, _12792_, _09115_);
  or (_32356_, _32328_, _06117_);
  or (_32357_, _32356_, _32355_);
  and (_32358_, _32357_, _06114_);
  and (_32359_, _32358_, _32354_);
  and (_32360_, _29883_, _12792_);
  or (_32361_, _32360_, _32328_);
  and (_32362_, _32361_, _05787_);
  or (_32363_, _32362_, _32359_);
  and (_32365_, _32363_, _06298_);
  or (_32366_, _30823_, _13196_);
  and (_32367_, _32366_, _06297_);
  nand (_32368_, _12792_, _06945_);
  and (_32369_, _32368_, _06110_);
  or (_32370_, _32369_, _32367_);
  and (_32371_, _32370_, _32310_);
  or (_32372_, _32371_, _32365_);
  and (_32373_, _32372_, _07125_);
  or (_32374_, _30833_, _13196_);
  and (_32376_, _32310_, _06402_);
  and (_32377_, _32376_, _32374_);
  or (_32378_, _32377_, _32373_);
  and (_32379_, _32378_, _07132_);
  or (_32380_, _29896_, _13196_);
  and (_32381_, _32310_, _06306_);
  and (_32382_, _32381_, _32380_);
  or (_32383_, _32382_, _32379_);
  and (_32384_, _32383_, _07130_);
  or (_32385_, _32328_, _12850_);
  and (_32387_, _32316_, _06411_);
  and (_32388_, _32387_, _32385_);
  or (_32389_, _32388_, _32384_);
  and (_32390_, _32389_, _06397_);
  or (_32391_, _32368_, _12850_);
  and (_32392_, _32310_, _06303_);
  and (_32393_, _32392_, _32391_);
  or (_32394_, _32315_, _12850_);
  and (_32395_, _32310_, _06396_);
  and (_32396_, _32395_, _32394_);
  or (_32398_, _32396_, _06433_);
  or (_32399_, _32398_, _32393_);
  or (_32400_, _32399_, _32390_);
  or (_32401_, _32313_, _06829_);
  and (_32402_, _32401_, _05749_);
  and (_32403_, _32402_, _32400_);
  and (_32404_, _32339_, _05748_);
  or (_32405_, _32404_, _06440_);
  or (_32406_, _32405_, _32403_);
  or (_32407_, _32328_, _06444_);
  or (_32409_, _32407_, _32311_);
  and (_32410_, _32409_, _01317_);
  and (_32411_, _32410_, _32406_);
  nor (_32412_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_32413_, _32412_, _00000_);
  or (_43731_, _32413_, _32411_);
  and (_32414_, _13196_, \oc8051_golden_model_1.P1 [2]);
  and (_32415_, _12792_, _07708_);
  or (_32416_, _32415_, _32414_);
  or (_32417_, _32416_, _06132_);
  and (_32419_, _29954_, _12792_);
  or (_32420_, _32419_, _32414_);
  or (_32421_, _32420_, _06161_);
  and (_32422_, _12792_, \oc8051_golden_model_1.ACC [2]);
  or (_32423_, _32422_, _32414_);
  and (_32424_, _32423_, _07056_);
  and (_32425_, _07057_, \oc8051_golden_model_1.P1 [2]);
  or (_32426_, _32425_, _06160_);
  or (_32427_, _32426_, _32424_);
  and (_32428_, _32427_, _06157_);
  and (_32430_, _32428_, _32421_);
  and (_32431_, _13201_, \oc8051_golden_model_1.P1 [2]);
  and (_32432_, _29976_, _12778_);
  or (_32433_, _32432_, _32431_);
  and (_32434_, _32433_, _06156_);
  or (_32435_, _32434_, _06217_);
  or (_32436_, _32435_, _32430_);
  or (_32437_, _32416_, _07075_);
  and (_32438_, _32437_, _32436_);
  or (_32439_, _32438_, _06220_);
  or (_32441_, _32423_, _06229_);
  and (_32442_, _32441_, _06153_);
  and (_32443_, _32442_, _32439_);
  and (_32444_, _29992_, _12778_);
  or (_32445_, _32444_, _32431_);
  and (_32446_, _32445_, _06152_);
  or (_32447_, _32446_, _06145_);
  or (_32448_, _32447_, _32443_);
  or (_32449_, _32431_, _29999_);
  and (_32450_, _32449_, _32433_);
  or (_32452_, _32450_, _06146_);
  and (_32453_, _32452_, _06140_);
  and (_32454_, _32453_, _32448_);
  and (_32455_, _30005_, _12778_);
  or (_32456_, _32455_, _32431_);
  and (_32457_, _32456_, _06139_);
  or (_32458_, _32457_, _09842_);
  or (_32459_, _32458_, _32454_);
  and (_32460_, _32459_, _32417_);
  or (_32461_, _32460_, _06116_);
  and (_32463_, _12792_, _09211_);
  or (_32464_, _32414_, _06117_);
  or (_32465_, _32464_, _32463_);
  and (_32466_, _32465_, _06114_);
  and (_32467_, _32466_, _32461_);
  and (_32468_, _30029_, _12792_);
  or (_32469_, _32414_, _32468_);
  and (_32470_, _32469_, _05787_);
  or (_32471_, _32470_, _32467_);
  or (_32472_, _32471_, _11136_);
  and (_32474_, _31708_, _12792_);
  or (_32475_, _32414_, _07127_);
  or (_32476_, _32475_, _32474_);
  and (_32477_, _12792_, _08768_);
  or (_32478_, _32477_, _32414_);
  or (_32479_, _32478_, _06111_);
  and (_32480_, _32479_, _07125_);
  and (_32481_, _32480_, _32476_);
  and (_32482_, _32481_, _32472_);
  and (_32483_, _30043_, _12792_);
  or (_32485_, _32483_, _32414_);
  or (_32486_, _32414_, _30046_);
  and (_32487_, _32486_, _06402_);
  and (_32488_, _32487_, _32485_);
  or (_32489_, _32488_, _32482_);
  and (_32490_, _32489_, _07132_);
  or (_32491_, _32414_, _12842_);
  and (_32492_, _32478_, _06306_);
  and (_32493_, _32492_, _32491_);
  or (_32494_, _32493_, _32490_);
  and (_32496_, _32494_, _07130_);
  and (_32497_, _32423_, _06411_);
  and (_32498_, _32497_, _32491_);
  or (_32499_, _32498_, _06303_);
  or (_32500_, _32499_, _32496_);
  and (_32501_, _29945_, _12792_);
  or (_32502_, _32414_, _08819_);
  or (_32503_, _32502_, _32501_);
  and (_32504_, _32503_, _08824_);
  and (_32505_, _32504_, _32500_);
  and (_32507_, _32485_, _06396_);
  or (_32508_, _32507_, _06433_);
  or (_32509_, _32508_, _32505_);
  or (_32510_, _32420_, _06829_);
  and (_32511_, _32510_, _05749_);
  and (_32512_, _32511_, _32509_);
  and (_32513_, _32445_, _05748_);
  or (_32514_, _32513_, _06440_);
  or (_32515_, _32514_, _32512_);
  and (_32516_, _30077_, _12792_);
  or (_32518_, _32414_, _06444_);
  or (_32519_, _32518_, _32516_);
  and (_32520_, _32519_, _01317_);
  and (_32521_, _32520_, _32515_);
  nor (_32522_, \oc8051_golden_model_1.P1 [2], rst);
  nor (_32523_, _32522_, _00000_);
  or (_43732_, _32523_, _32521_);
  nor (_32524_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_32525_, _32524_, _00000_);
  and (_32526_, _13196_, \oc8051_golden_model_1.P1 [3]);
  and (_32528_, _12792_, _07544_);
  or (_32529_, _32528_, _32526_);
  or (_32530_, _32529_, _06132_);
  and (_32531_, _13201_, \oc8051_golden_model_1.P1 [3]);
  and (_32532_, _30100_, _12778_);
  or (_32533_, _32532_, _32531_);
  and (_32534_, _32533_, _06152_);
  and (_32535_, _30106_, _12792_);
  or (_32536_, _32535_, _32526_);
  or (_32537_, _32536_, _06161_);
  and (_32539_, _12792_, \oc8051_golden_model_1.ACC [3]);
  or (_32540_, _32539_, _32526_);
  and (_32541_, _32540_, _07056_);
  and (_32542_, _07057_, \oc8051_golden_model_1.P1 [3]);
  or (_32543_, _32542_, _06160_);
  or (_32544_, _32543_, _32541_);
  and (_32545_, _32544_, _06157_);
  and (_32546_, _32545_, _32537_);
  and (_32547_, _30119_, _12778_);
  or (_32548_, _32547_, _32531_);
  and (_32550_, _32548_, _06156_);
  or (_32551_, _32550_, _06217_);
  or (_32552_, _32551_, _32546_);
  or (_32553_, _32529_, _07075_);
  and (_32554_, _32553_, _32552_);
  or (_32555_, _32554_, _06220_);
  or (_32556_, _32540_, _06229_);
  and (_32557_, _32556_, _06153_);
  and (_32558_, _32557_, _32555_);
  or (_32559_, _32558_, _32534_);
  and (_32561_, _32559_, _06146_);
  or (_32562_, _32531_, _30134_);
  and (_32563_, _32548_, _06145_);
  and (_32564_, _32563_, _32562_);
  or (_32565_, _32564_, _32561_);
  and (_32566_, _32565_, _06140_);
  and (_32567_, _30141_, _12778_);
  or (_32568_, _32567_, _32531_);
  and (_32569_, _32568_, _06139_);
  or (_32570_, _32569_, _09842_);
  or (_32572_, _32570_, _32566_);
  and (_32573_, _32572_, _32530_);
  or (_32574_, _32573_, _06116_);
  and (_32575_, _12792_, _09210_);
  or (_32576_, _32526_, _06117_);
  or (_32577_, _32576_, _32575_);
  and (_32578_, _32577_, _06114_);
  and (_32579_, _32578_, _32574_);
  and (_32580_, _30163_, _12792_);
  or (_32581_, _32580_, _32526_);
  and (_32583_, _32581_, _05787_);
  or (_32584_, _32583_, _11136_);
  or (_32585_, _32584_, _32579_);
  and (_32586_, _31042_, _12792_);
  or (_32587_, _32526_, _07127_);
  or (_32588_, _32587_, _32586_);
  and (_32589_, _12792_, _08712_);
  or (_32590_, _32589_, _32526_);
  or (_32591_, _32590_, _06111_);
  and (_32592_, _32591_, _07125_);
  and (_32594_, _32592_, _32588_);
  and (_32595_, _32594_, _32585_);
  and (_32596_, _31053_, _12792_);
  or (_32597_, _32596_, _32526_);
  and (_32598_, _32597_, _06402_);
  or (_32599_, _32598_, _32595_);
  and (_32600_, _32599_, _07132_);
  or (_32601_, _32526_, _12834_);
  and (_32602_, _32590_, _06306_);
  and (_32603_, _32602_, _32601_);
  or (_32605_, _32603_, _32600_);
  and (_32606_, _32605_, _07130_);
  and (_32607_, _32540_, _06411_);
  and (_32608_, _32607_, _32601_);
  or (_32609_, _32608_, _06303_);
  or (_32610_, _32609_, _32606_);
  and (_32611_, _30175_, _12792_);
  or (_32612_, _32526_, _08819_);
  or (_32613_, _32612_, _32611_);
  and (_32614_, _32613_, _08824_);
  and (_32616_, _32614_, _32610_);
  and (_32617_, _30185_, _12792_);
  or (_32618_, _32617_, _32526_);
  and (_32619_, _32618_, _06396_);
  or (_32620_, _32619_, _06433_);
  or (_32621_, _32620_, _32616_);
  or (_32622_, _32536_, _06829_);
  and (_32623_, _32622_, _05749_);
  and (_32624_, _32623_, _32621_);
  and (_32625_, _32533_, _05748_);
  or (_32627_, _32625_, _06440_);
  or (_32628_, _32627_, _32624_);
  and (_32629_, _30219_, _12792_);
  or (_32630_, _32526_, _06444_);
  or (_32631_, _32630_, _32629_);
  and (_32632_, _32631_, _01317_);
  and (_32633_, _32632_, _32628_);
  or (_43733_, _32633_, _32525_);
  and (_32634_, _13196_, \oc8051_golden_model_1.P1 [4]);
  and (_32635_, _12792_, _08336_);
  or (_32637_, _32635_, _32634_);
  or (_32638_, _32637_, _06132_);
  and (_32639_, _13201_, \oc8051_golden_model_1.P1 [4]);
  and (_32640_, _30242_, _12778_);
  or (_32641_, _32640_, _32639_);
  and (_32642_, _32641_, _06152_);
  and (_32643_, _30248_, _12792_);
  or (_32644_, _32643_, _32634_);
  or (_32645_, _32644_, _06161_);
  and (_32646_, _12792_, \oc8051_golden_model_1.ACC [4]);
  or (_32648_, _32646_, _32634_);
  and (_32649_, _32648_, _07056_);
  and (_32650_, _07057_, \oc8051_golden_model_1.P1 [4]);
  or (_32651_, _32650_, _06160_);
  or (_32652_, _32651_, _32649_);
  and (_32653_, _32652_, _06157_);
  and (_32654_, _32653_, _32645_);
  and (_32655_, _30261_, _12778_);
  or (_32656_, _32655_, _32639_);
  and (_32657_, _32656_, _06156_);
  or (_32659_, _32657_, _06217_);
  or (_32660_, _32659_, _32654_);
  or (_32661_, _32637_, _07075_);
  and (_32662_, _32661_, _32660_);
  or (_32663_, _32662_, _06220_);
  or (_32664_, _32648_, _06229_);
  and (_32665_, _32664_, _06153_);
  and (_32666_, _32665_, _32663_);
  or (_32667_, _32666_, _32642_);
  and (_32668_, _32667_, _06146_);
  or (_32670_, _32639_, _30276_);
  and (_32671_, _32656_, _06145_);
  and (_32672_, _32671_, _32670_);
  or (_32673_, _32672_, _32668_);
  and (_32674_, _32673_, _06140_);
  and (_32675_, _30283_, _12778_);
  or (_32676_, _32675_, _32639_);
  and (_32677_, _32676_, _06139_);
  or (_32678_, _32677_, _09842_);
  or (_32679_, _32678_, _32674_);
  and (_32681_, _32679_, _32638_);
  or (_32682_, _32681_, _06116_);
  and (_32683_, _12792_, _09209_);
  or (_32684_, _32634_, _06117_);
  or (_32685_, _32684_, _32683_);
  and (_32686_, _32685_, _06114_);
  and (_32687_, _32686_, _32682_);
  and (_32688_, _30305_, _12792_);
  or (_32689_, _32688_, _32634_);
  and (_32690_, _32689_, _05787_);
  or (_32691_, _32690_, _06110_);
  or (_32692_, _32691_, _32687_);
  and (_32693_, _12792_, _08715_);
  or (_32694_, _32693_, _32634_);
  or (_32695_, _32694_, _06111_);
  and (_32696_, _32695_, _07127_);
  and (_32697_, _32696_, _32692_);
  and (_32698_, _30317_, _12792_);
  or (_32699_, _32698_, _32634_);
  or (_32700_, _32634_, _30320_);
  and (_32702_, _32700_, _06297_);
  and (_32703_, _32702_, _32699_);
  or (_32704_, _32703_, _06402_);
  or (_32705_, _32704_, _32697_);
  and (_32706_, _31172_, _12792_);
  or (_32707_, _32634_, _07125_);
  or (_32708_, _32707_, _32706_);
  and (_32709_, _32708_, _07132_);
  and (_32710_, _32709_, _32705_);
  or (_32711_, _32634_, _12826_);
  and (_32713_, _32694_, _06306_);
  and (_32714_, _32713_, _32711_);
  or (_32715_, _32714_, _32710_);
  and (_32716_, _32715_, _07130_);
  and (_32717_, _32648_, _06411_);
  and (_32718_, _32717_, _32711_);
  or (_32719_, _32718_, _06303_);
  or (_32720_, _32719_, _32716_);
  or (_32721_, _32699_, _08819_);
  and (_32722_, _32721_, _08824_);
  and (_32724_, _32722_, _32720_);
  and (_32725_, _30327_, _12792_);
  or (_32726_, _32725_, _32634_);
  and (_32727_, _32726_, _06396_);
  or (_32728_, _32727_, _06433_);
  or (_32729_, _32728_, _32724_);
  or (_32730_, _32644_, _06829_);
  and (_32731_, _32730_, _05749_);
  and (_32732_, _32731_, _32729_);
  and (_32733_, _32641_, _05748_);
  or (_32735_, _32733_, _06440_);
  or (_32736_, _32735_, _32732_);
  and (_32737_, _30361_, _12792_);
  or (_32738_, _32634_, _06444_);
  or (_32739_, _32738_, _32737_);
  and (_32740_, _32739_, _01317_);
  and (_32741_, _32740_, _32736_);
  nor (_32742_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_32743_, _32742_, _00000_);
  or (_43734_, _32743_, _32741_);
  and (_32745_, _13196_, \oc8051_golden_model_1.P1 [5]);
  and (_32746_, _12792_, _08101_);
  or (_32747_, _32746_, _32745_);
  or (_32748_, _32747_, _06132_);
  and (_32749_, _30378_, _12792_);
  or (_32750_, _32749_, _32745_);
  or (_32751_, _32750_, _06161_);
  and (_32752_, _12792_, \oc8051_golden_model_1.ACC [5]);
  or (_32753_, _32752_, _32745_);
  and (_32754_, _32753_, _07056_);
  and (_32756_, _07057_, \oc8051_golden_model_1.P1 [5]);
  or (_32757_, _32756_, _06160_);
  or (_32758_, _32757_, _32754_);
  and (_32759_, _32758_, _06157_);
  and (_32760_, _32759_, _32751_);
  and (_32761_, _13201_, \oc8051_golden_model_1.P1 [5]);
  and (_32762_, _30400_, _12778_);
  or (_32763_, _32762_, _32761_);
  and (_32764_, _32763_, _06156_);
  or (_32765_, _32764_, _06217_);
  or (_32767_, _32765_, _32760_);
  or (_32768_, _32747_, _07075_);
  and (_32769_, _32768_, _32767_);
  or (_32770_, _32769_, _06220_);
  or (_32771_, _32753_, _06229_);
  and (_32772_, _32771_, _06153_);
  and (_32773_, _32772_, _32770_);
  and (_32774_, _30414_, _12778_);
  or (_32775_, _32774_, _32761_);
  and (_32776_, _32775_, _06152_);
  or (_32778_, _32776_, _06145_);
  or (_32779_, _32778_, _32773_);
  or (_32780_, _32761_, _30420_);
  and (_32781_, _32780_, _32763_);
  or (_32782_, _32781_, _06146_);
  and (_32783_, _32782_, _06140_);
  and (_32784_, _32783_, _32779_);
  and (_32785_, _30426_, _12778_);
  or (_32786_, _32785_, _32761_);
  and (_32787_, _32786_, _06139_);
  or (_32789_, _32787_, _09842_);
  or (_32790_, _32789_, _32784_);
  and (_32791_, _32790_, _32748_);
  or (_32792_, _32791_, _06116_);
  and (_32793_, _12792_, _09208_);
  or (_32794_, _32745_, _06117_);
  or (_32795_, _32794_, _32793_);
  and (_32796_, _32795_, _06114_);
  and (_32797_, _32796_, _32792_);
  and (_32798_, _30449_, _12792_);
  or (_32800_, _32798_, _32745_);
  and (_32801_, _32800_, _05787_);
  or (_32802_, _32801_, _11136_);
  or (_32803_, _32802_, _32797_);
  and (_32804_, _32036_, _12792_);
  or (_32805_, _32745_, _07127_);
  or (_32806_, _32805_, _32804_);
  and (_32807_, _12792_, _08736_);
  or (_32808_, _32807_, _32745_);
  or (_32809_, _32808_, _06111_);
  and (_32811_, _32809_, _07125_);
  and (_32812_, _32811_, _32806_);
  and (_32813_, _32812_, _32803_);
  and (_32814_, _32047_, _12792_);
  or (_32815_, _32814_, _32745_);
  and (_32816_, _32815_, _06402_);
  or (_32817_, _32816_, _32813_);
  and (_32818_, _32817_, _07132_);
  or (_32819_, _32745_, _12818_);
  and (_32820_, _32808_, _06306_);
  and (_32822_, _32820_, _32819_);
  or (_32823_, _32822_, _32818_);
  and (_32824_, _32823_, _07130_);
  and (_32825_, _32753_, _06411_);
  and (_32826_, _32825_, _32819_);
  or (_32827_, _32826_, _06303_);
  or (_32828_, _32827_, _32824_);
  and (_32829_, _30461_, _12792_);
  or (_32830_, _32745_, _08819_);
  or (_32831_, _32830_, _32829_);
  and (_32833_, _32831_, _08824_);
  and (_32834_, _32833_, _32828_);
  and (_32835_, _30471_, _12792_);
  or (_32836_, _32835_, _32745_);
  and (_32837_, _32836_, _06396_);
  or (_32838_, _32837_, _06433_);
  or (_32839_, _32838_, _32834_);
  or (_32840_, _32750_, _06829_);
  and (_32841_, _32840_, _05749_);
  and (_32842_, _32841_, _32839_);
  and (_32844_, _32775_, _05748_);
  or (_32845_, _32844_, _06440_);
  or (_32846_, _32845_, _32842_);
  and (_32847_, _30505_, _12792_);
  or (_32848_, _32745_, _06444_);
  or (_32849_, _32848_, _32847_);
  and (_32850_, _32849_, _01317_);
  and (_32851_, _32850_, _32846_);
  nor (_32852_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_32853_, _32852_, _00000_);
  or (_43735_, _32853_, _32851_);
  and (_32855_, _13196_, \oc8051_golden_model_1.P1 [6]);
  and (_32856_, _12792_, _08012_);
  or (_32857_, _32856_, _32855_);
  or (_32858_, _32857_, _06132_);
  and (_32859_, _13201_, \oc8051_golden_model_1.P1 [6]);
  and (_32860_, _30526_, _12778_);
  or (_32861_, _32860_, _32859_);
  and (_32862_, _32861_, _06152_);
  and (_32863_, _30532_, _12792_);
  or (_32865_, _32863_, _32855_);
  or (_32866_, _32865_, _06161_);
  and (_32867_, _12792_, \oc8051_golden_model_1.ACC [6]);
  or (_32868_, _32867_, _32855_);
  and (_32869_, _32868_, _07056_);
  and (_32870_, _07057_, \oc8051_golden_model_1.P1 [6]);
  or (_32871_, _32870_, _06160_);
  or (_32872_, _32871_, _32869_);
  and (_32873_, _32872_, _06157_);
  and (_32874_, _32873_, _32866_);
  and (_32876_, _30545_, _12778_);
  or (_32877_, _32876_, _32859_);
  and (_32878_, _32877_, _06156_);
  or (_32879_, _32878_, _06217_);
  or (_32880_, _32879_, _32874_);
  or (_32881_, _32857_, _07075_);
  and (_32882_, _32881_, _32880_);
  or (_32883_, _32882_, _06220_);
  or (_32884_, _32868_, _06229_);
  and (_32885_, _32884_, _06153_);
  and (_32887_, _32885_, _32883_);
  or (_32888_, _32887_, _32862_);
  and (_32889_, _32888_, _06146_);
  or (_32890_, _32859_, _30560_);
  and (_32891_, _32877_, _06145_);
  and (_32892_, _32891_, _32890_);
  or (_32893_, _32892_, _32889_);
  and (_32894_, _32893_, _06140_);
  and (_32895_, _30567_, _12778_);
  or (_32896_, _32895_, _32859_);
  and (_32898_, _32896_, _06139_);
  or (_32899_, _32898_, _09842_);
  or (_32900_, _32899_, _32894_);
  and (_32901_, _32900_, _32858_);
  or (_32902_, _32901_, _06116_);
  and (_32903_, _12792_, _09207_);
  or (_32904_, _32855_, _06117_);
  or (_32905_, _32904_, _32903_);
  and (_32906_, _32905_, _06114_);
  and (_32907_, _32906_, _32902_);
  and (_32909_, _30589_, _12792_);
  or (_32910_, _32909_, _32855_);
  and (_32911_, _32910_, _05787_);
  or (_32912_, _32911_, _11136_);
  or (_32913_, _32912_, _32907_);
  and (_32914_, _32151_, _12792_);
  or (_32915_, _32855_, _07127_);
  or (_32916_, _32915_, _32914_);
  and (_32917_, _12792_, _15402_);
  or (_32918_, _32917_, _32855_);
  or (_32920_, _32918_, _06111_);
  and (_32921_, _32920_, _07125_);
  and (_32922_, _32921_, _32916_);
  and (_32923_, _32922_, _32913_);
  and (_32924_, _30613_, _12792_);
  or (_32925_, _32924_, _32855_);
  and (_32926_, _32925_, _06402_);
  or (_32927_, _32926_, _32923_);
  and (_32928_, _32927_, _07132_);
  or (_32929_, _32855_, _12810_);
  and (_32931_, _32918_, _06306_);
  and (_32932_, _32931_, _32929_);
  or (_32933_, _32932_, _32928_);
  and (_32934_, _32933_, _07130_);
  and (_32935_, _32868_, _06411_);
  and (_32936_, _32935_, _32929_);
  or (_32937_, _32936_, _06303_);
  or (_32938_, _32937_, _32934_);
  and (_32939_, _30601_, _12792_);
  or (_32940_, _32855_, _08819_);
  or (_32942_, _32940_, _32939_);
  and (_32943_, _32942_, _08824_);
  and (_32944_, _32943_, _32938_);
  and (_32945_, _30611_, _12792_);
  or (_32946_, _32945_, _32855_);
  and (_32947_, _32946_, _06396_);
  or (_32948_, _32947_, _06433_);
  or (_32949_, _32948_, _32944_);
  or (_32950_, _32865_, _06829_);
  and (_32951_, _32950_, _05749_);
  and (_32953_, _32951_, _32949_);
  and (_32954_, _32861_, _05748_);
  or (_32955_, _32954_, _06440_);
  or (_32956_, _32955_, _32953_);
  and (_32957_, _30646_, _12792_);
  or (_32958_, _32855_, _06444_);
  or (_32959_, _32958_, _32957_);
  and (_32960_, _32959_, _01317_);
  and (_32961_, _32960_, _32956_);
  nor (_32962_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_32964_, _32962_, _00000_);
  or (_43736_, _32964_, _32961_);
  not (_32965_, \oc8051_golden_model_1.IP [0]);
  nor (_32966_, _01317_, _32965_);
  nand (_32967_, _10276_, _07830_);
  nor (_32968_, _07830_, _32965_);
  nor (_32969_, _32968_, _07130_);
  nand (_32970_, _32969_, _32967_);
  and (_32971_, _07830_, _07049_);
  or (_32972_, _32971_, _32968_);
  or (_32974_, _32972_, _06132_);
  nor (_32975_, _08211_, _13300_);
  or (_32976_, _32975_, _32968_);
  or (_32977_, _32976_, _06161_);
  and (_32978_, _07830_, \oc8051_golden_model_1.ACC [0]);
  or (_32979_, _32978_, _32968_);
  and (_32980_, _32979_, _07056_);
  nor (_32981_, _07056_, _32965_);
  or (_32982_, _32981_, _06160_);
  or (_32983_, _32982_, _32980_);
  and (_32985_, _32983_, _06157_);
  and (_32986_, _32985_, _32977_);
  nor (_32987_, _08415_, _32965_);
  and (_32988_, _14169_, _08415_);
  or (_32989_, _32988_, _32987_);
  and (_32990_, _32989_, _06156_);
  or (_32991_, _32990_, _32986_);
  and (_32992_, _32991_, _07075_);
  and (_32993_, _32972_, _06217_);
  or (_32994_, _32993_, _06220_);
  or (_32996_, _32994_, _32992_);
  or (_32997_, _32979_, _06229_);
  and (_32998_, _32997_, _06153_);
  and (_32999_, _32998_, _32996_);
  and (_33000_, _32968_, _06152_);
  or (_33001_, _33000_, _06145_);
  or (_33002_, _33001_, _32999_);
  or (_33003_, _32976_, _06146_);
  and (_33004_, _33003_, _06140_);
  and (_33005_, _33004_, _33002_);
  or (_33007_, _32987_, _14170_);
  and (_33008_, _33007_, _06139_);
  and (_33009_, _33008_, _32989_);
  or (_33010_, _33009_, _09842_);
  or (_33011_, _33010_, _33005_);
  and (_33012_, _33011_, _32974_);
  or (_33013_, _33012_, _06116_);
  and (_33014_, _09160_, _07830_);
  or (_33015_, _32968_, _06117_);
  or (_33016_, _33015_, _33014_);
  and (_33018_, _33016_, _06114_);
  and (_33019_, _33018_, _33013_);
  and (_33020_, _14260_, _07830_);
  or (_33021_, _33020_, _32968_);
  and (_33022_, _33021_, _05787_);
  or (_33023_, _33022_, _33019_);
  or (_33024_, _33023_, _11136_);
  and (_33025_, _14275_, _07830_);
  or (_33026_, _32968_, _07127_);
  or (_33027_, _33026_, _33025_);
  and (_33029_, _07830_, _08708_);
  or (_33030_, _33029_, _32968_);
  or (_33031_, _33030_, _06111_);
  and (_33032_, _33031_, _07125_);
  and (_33033_, _33032_, _33027_);
  and (_33034_, _33033_, _33024_);
  nor (_33035_, _12321_, _13300_);
  or (_33036_, _33035_, _32968_);
  and (_33037_, _32967_, _06402_);
  and (_33038_, _33037_, _33036_);
  or (_33040_, _33038_, _33034_);
  and (_33041_, _33040_, _07132_);
  nand (_33042_, _33030_, _06306_);
  nor (_33043_, _33042_, _32975_);
  or (_33044_, _33043_, _06411_);
  or (_33045_, _33044_, _33041_);
  and (_33046_, _33045_, _32970_);
  or (_33047_, _33046_, _06303_);
  and (_33048_, _14167_, _07830_);
  or (_33049_, _32968_, _08819_);
  or (_33051_, _33049_, _33048_);
  and (_33052_, _33051_, _08824_);
  and (_33053_, _33052_, _33047_);
  and (_33054_, _33036_, _06396_);
  or (_33055_, _33054_, _06433_);
  or (_33056_, _33055_, _33053_);
  or (_33057_, _32976_, _06829_);
  and (_33058_, _33057_, _33056_);
  or (_33059_, _33058_, _05748_);
  or (_33060_, _32968_, _05749_);
  and (_33062_, _33060_, _33059_);
  or (_33063_, _33062_, _06440_);
  or (_33064_, _32976_, _06444_);
  and (_33065_, _33064_, _01317_);
  and (_33066_, _33065_, _33063_);
  or (_33067_, _33066_, _32966_);
  and (_43738_, _33067_, _43100_);
  not (_33068_, \oc8051_golden_model_1.IP [1]);
  nor (_33069_, _01317_, _33068_);
  nor (_33070_, _07830_, _33068_);
  nor (_33072_, _10277_, _13300_);
  or (_33073_, _33072_, _33070_);
  or (_33074_, _33073_, _08824_);
  or (_33075_, _14442_, _13300_);
  or (_33076_, _07830_, \oc8051_golden_model_1.IP [1]);
  and (_33077_, _33076_, _05787_);
  and (_33078_, _33077_, _33075_);
  and (_33079_, _07830_, _07306_);
  or (_33080_, _33079_, _33070_);
  or (_33081_, _33080_, _07075_);
  and (_33083_, _14363_, _07830_);
  not (_33084_, _33083_);
  and (_33085_, _33084_, _33076_);
  or (_33086_, _33085_, _06161_);
  and (_33087_, _07830_, \oc8051_golden_model_1.ACC [1]);
  or (_33088_, _33087_, _33070_);
  and (_33089_, _33088_, _07056_);
  nor (_33090_, _07056_, _33068_);
  or (_33091_, _33090_, _06160_);
  or (_33092_, _33091_, _33089_);
  and (_33094_, _33092_, _06157_);
  and (_33095_, _33094_, _33086_);
  nor (_33096_, _08415_, _33068_);
  and (_33097_, _14367_, _08415_);
  or (_33098_, _33097_, _33096_);
  and (_33099_, _33098_, _06156_);
  or (_33100_, _33099_, _06217_);
  or (_33101_, _33100_, _33095_);
  and (_33102_, _33101_, _33081_);
  or (_33103_, _33102_, _06220_);
  or (_33105_, _33088_, _06229_);
  and (_33106_, _33105_, _06153_);
  and (_33107_, _33106_, _33103_);
  and (_33108_, _14349_, _08415_);
  or (_33109_, _33108_, _33096_);
  and (_33110_, _33109_, _06152_);
  or (_33111_, _33110_, _06145_);
  or (_33112_, _33111_, _33107_);
  and (_33113_, _33097_, _14382_);
  or (_33114_, _33096_, _06146_);
  or (_33116_, _33114_, _33113_);
  and (_33117_, _33116_, _33112_);
  and (_33118_, _33117_, _06140_);
  and (_33119_, _14351_, _08415_);
  or (_33120_, _33096_, _33119_);
  and (_33121_, _33120_, _06139_);
  or (_33122_, _33121_, _09842_);
  or (_33123_, _33122_, _33118_);
  or (_33124_, _33080_, _06132_);
  and (_33125_, _33124_, _33123_);
  or (_33127_, _33125_, _06116_);
  and (_33128_, _09115_, _07830_);
  or (_33129_, _33070_, _06117_);
  or (_33130_, _33129_, _33128_);
  and (_33131_, _33130_, _06114_);
  and (_33132_, _33131_, _33127_);
  or (_33133_, _33132_, _33078_);
  and (_33134_, _33133_, _06298_);
  or (_33135_, _14346_, _13300_);
  and (_33136_, _33135_, _06297_);
  nand (_33138_, _07830_, _06945_);
  and (_33139_, _33138_, _06110_);
  or (_33140_, _33139_, _33136_);
  and (_33141_, _33140_, _33076_);
  or (_33142_, _33141_, _06402_);
  or (_33143_, _33142_, _33134_);
  nand (_33144_, _10275_, _07830_);
  and (_33145_, _33144_, _33073_);
  or (_33146_, _33145_, _07125_);
  and (_33147_, _33146_, _07132_);
  and (_33149_, _33147_, _33143_);
  or (_33150_, _14344_, _13300_);
  and (_33151_, _33076_, _06306_);
  and (_33152_, _33151_, _33150_);
  or (_33153_, _33152_, _06411_);
  or (_33154_, _33153_, _33149_);
  nor (_33155_, _33070_, _07130_);
  nand (_33156_, _33155_, _33144_);
  and (_33157_, _33156_, _08819_);
  and (_33158_, _33157_, _33154_);
  or (_33160_, _33138_, _08176_);
  and (_33161_, _33076_, _06303_);
  and (_33162_, _33161_, _33160_);
  or (_33163_, _33162_, _06396_);
  or (_33164_, _33163_, _33158_);
  and (_33165_, _33164_, _33074_);
  or (_33166_, _33165_, _06433_);
  or (_33167_, _33085_, _06829_);
  and (_33168_, _33167_, _05749_);
  and (_33169_, _33168_, _33166_);
  and (_33171_, _33109_, _05748_);
  or (_33172_, _33171_, _06440_);
  or (_33173_, _33172_, _33169_);
  or (_33174_, _33070_, _06444_);
  or (_33175_, _33174_, _33083_);
  and (_33176_, _33175_, _01317_);
  and (_33177_, _33176_, _33173_);
  or (_33178_, _33177_, _33069_);
  and (_43739_, _33178_, _43100_);
  and (_33179_, _01321_, \oc8051_golden_model_1.IP [2]);
  and (_33181_, _13300_, \oc8051_golden_model_1.IP [2]);
  and (_33182_, _07830_, _07708_);
  or (_33183_, _33182_, _33181_);
  or (_33184_, _33183_, _06132_);
  or (_33185_, _33183_, _07075_);
  and (_33186_, _14542_, _07830_);
  or (_33187_, _33186_, _33181_);
  or (_33188_, _33187_, _06161_);
  and (_33189_, _07830_, \oc8051_golden_model_1.ACC [2]);
  or (_33190_, _33189_, _33181_);
  and (_33192_, _33190_, _07056_);
  and (_33193_, _07057_, \oc8051_golden_model_1.IP [2]);
  or (_33194_, _33193_, _06160_);
  or (_33195_, _33194_, _33192_);
  and (_33196_, _33195_, _06157_);
  and (_33197_, _33196_, _33188_);
  and (_33198_, _13305_, \oc8051_golden_model_1.IP [2]);
  and (_33199_, _14538_, _08415_);
  or (_33200_, _33199_, _33198_);
  and (_33201_, _33200_, _06156_);
  or (_33203_, _33201_, _06217_);
  or (_33204_, _33203_, _33197_);
  and (_33205_, _33204_, _33185_);
  or (_33206_, _33205_, _06220_);
  or (_33207_, _33190_, _06229_);
  and (_33208_, _33207_, _06153_);
  and (_33209_, _33208_, _33206_);
  and (_33210_, _14536_, _08415_);
  or (_33211_, _33210_, _33198_);
  and (_33212_, _33211_, _06152_);
  or (_33214_, _33212_, _06145_);
  or (_33215_, _33214_, _33209_);
  and (_33216_, _33199_, _14569_);
  or (_33217_, _33198_, _06146_);
  or (_33218_, _33217_, _33216_);
  and (_33219_, _33218_, _06140_);
  and (_33220_, _33219_, _33215_);
  and (_33221_, _14583_, _08415_);
  or (_33222_, _33221_, _33198_);
  and (_33223_, _33222_, _06139_);
  or (_33225_, _33223_, _09842_);
  or (_33226_, _33225_, _33220_);
  and (_33227_, _33226_, _33184_);
  or (_33228_, _33227_, _06116_);
  and (_33229_, _09211_, _07830_);
  or (_33230_, _33181_, _06117_);
  or (_33231_, _33230_, _33229_);
  and (_33232_, _33231_, _06114_);
  and (_33233_, _33232_, _33228_);
  and (_33234_, _14630_, _07830_);
  or (_33236_, _33181_, _33234_);
  and (_33237_, _33236_, _05787_);
  or (_33238_, _33237_, _33233_);
  or (_33239_, _33238_, _11136_);
  and (_33240_, _14646_, _07830_);
  or (_33241_, _33181_, _07127_);
  or (_33242_, _33241_, _33240_);
  and (_33243_, _07830_, _08768_);
  or (_33244_, _33243_, _33181_);
  or (_33245_, _33244_, _06111_);
  and (_33247_, _33245_, _07125_);
  and (_33248_, _33247_, _33242_);
  and (_33249_, _33248_, _33239_);
  and (_33250_, _10282_, _07830_);
  or (_33251_, _33250_, _33181_);
  and (_33252_, _33251_, _06402_);
  or (_33253_, _33252_, _33249_);
  and (_33254_, _33253_, _07132_);
  or (_33255_, _33181_, _08248_);
  and (_33256_, _33244_, _06306_);
  and (_33258_, _33256_, _33255_);
  or (_33259_, _33258_, _33254_);
  and (_33260_, _33259_, _07130_);
  and (_33261_, _33190_, _06411_);
  and (_33262_, _33261_, _33255_);
  or (_33263_, _33262_, _06303_);
  or (_33264_, _33263_, _33260_);
  and (_33265_, _14643_, _07830_);
  or (_33266_, _33181_, _08819_);
  or (_33267_, _33266_, _33265_);
  and (_33269_, _33267_, _08824_);
  and (_33270_, _33269_, _33264_);
  nor (_33271_, _10281_, _13300_);
  or (_33272_, _33271_, _33181_);
  and (_33273_, _33272_, _06396_);
  or (_33274_, _33273_, _06433_);
  or (_33275_, _33274_, _33270_);
  or (_33276_, _33187_, _06829_);
  and (_33277_, _33276_, _05749_);
  and (_33278_, _33277_, _33275_);
  and (_33280_, _33211_, _05748_);
  or (_33281_, _33280_, _06440_);
  or (_33282_, _33281_, _33278_);
  and (_33283_, _14710_, _07830_);
  or (_33284_, _33181_, _06444_);
  or (_33285_, _33284_, _33283_);
  and (_33286_, _33285_, _01317_);
  and (_33287_, _33286_, _33282_);
  or (_33288_, _33287_, _33179_);
  and (_43740_, _33288_, _43100_);
  and (_33290_, _01321_, \oc8051_golden_model_1.IP [3]);
  and (_33291_, _13300_, \oc8051_golden_model_1.IP [3]);
  and (_33292_, _07830_, _07544_);
  or (_33293_, _33292_, _33291_);
  or (_33294_, _33293_, _06132_);
  and (_33295_, _14738_, _07830_);
  or (_33296_, _33295_, _33291_);
  or (_33297_, _33296_, _06161_);
  and (_33298_, _07830_, \oc8051_golden_model_1.ACC [3]);
  or (_33299_, _33298_, _33291_);
  and (_33301_, _33299_, _07056_);
  and (_33302_, _07057_, \oc8051_golden_model_1.IP [3]);
  or (_33303_, _33302_, _06160_);
  or (_33304_, _33303_, _33301_);
  and (_33305_, _33304_, _06157_);
  and (_33306_, _33305_, _33297_);
  and (_33307_, _13305_, \oc8051_golden_model_1.IP [3]);
  and (_33308_, _14735_, _08415_);
  or (_33309_, _33308_, _33307_);
  and (_33310_, _33309_, _06156_);
  or (_33312_, _33310_, _06217_);
  or (_33313_, _33312_, _33306_);
  or (_33314_, _33293_, _07075_);
  and (_33315_, _33314_, _33313_);
  or (_33316_, _33315_, _06220_);
  or (_33317_, _33299_, _06229_);
  and (_33318_, _33317_, _06153_);
  and (_33319_, _33318_, _33316_);
  and (_33320_, _14731_, _08415_);
  or (_33321_, _33320_, _33307_);
  and (_33323_, _33321_, _06152_);
  or (_33324_, _33323_, _06145_);
  or (_33325_, _33324_, _33319_);
  or (_33326_, _33307_, _14764_);
  and (_33327_, _33326_, _33309_);
  or (_33328_, _33327_, _06146_);
  and (_33329_, _33328_, _06140_);
  and (_33330_, _33329_, _33325_);
  and (_33331_, _14732_, _08415_);
  or (_33332_, _33331_, _33307_);
  and (_33334_, _33332_, _06139_);
  or (_33335_, _33334_, _09842_);
  or (_33336_, _33335_, _33330_);
  and (_33337_, _33336_, _33294_);
  or (_33338_, _33337_, _06116_);
  and (_33339_, _09210_, _07830_);
  or (_33340_, _33291_, _06117_);
  or (_33341_, _33340_, _33339_);
  and (_33342_, _33341_, _06114_);
  and (_33343_, _33342_, _33338_);
  and (_33345_, _14825_, _07830_);
  or (_33346_, _33291_, _33345_);
  and (_33347_, _33346_, _05787_);
  or (_33348_, _33347_, _33343_);
  or (_33349_, _33348_, _11136_);
  and (_33350_, _14727_, _07830_);
  or (_33351_, _33291_, _07127_);
  or (_33352_, _33351_, _33350_);
  and (_33353_, _07830_, _08712_);
  or (_33354_, _33353_, _33291_);
  or (_33356_, _33354_, _06111_);
  and (_33357_, _33356_, _07125_);
  and (_33358_, _33357_, _33352_);
  and (_33359_, _33358_, _33349_);
  and (_33360_, _12318_, _07830_);
  or (_33361_, _33360_, _33291_);
  and (_33362_, _33361_, _06402_);
  or (_33363_, _33362_, _33359_);
  and (_33364_, _33363_, _07132_);
  or (_33365_, _33291_, _08140_);
  and (_33367_, _33354_, _06306_);
  and (_33368_, _33367_, _33365_);
  or (_33369_, _33368_, _33364_);
  and (_33370_, _33369_, _07130_);
  and (_33371_, _33299_, _06411_);
  and (_33372_, _33371_, _33365_);
  or (_33373_, _33372_, _06303_);
  or (_33374_, _33373_, _33370_);
  and (_33375_, _14724_, _07830_);
  or (_33376_, _33291_, _08819_);
  or (_33378_, _33376_, _33375_);
  and (_33379_, _33378_, _08824_);
  and (_33380_, _33379_, _33374_);
  nor (_33381_, _10273_, _13300_);
  or (_33382_, _33381_, _33291_);
  and (_33383_, _33382_, _06396_);
  or (_33384_, _33383_, _06433_);
  or (_33385_, _33384_, _33380_);
  or (_33386_, _33296_, _06829_);
  and (_33387_, _33386_, _05749_);
  and (_33389_, _33387_, _33385_);
  and (_33390_, _33321_, _05748_);
  or (_33391_, _33390_, _06440_);
  or (_33392_, _33391_, _33389_);
  and (_33393_, _14897_, _07830_);
  or (_33394_, _33291_, _06444_);
  or (_33395_, _33394_, _33393_);
  and (_33396_, _33395_, _01317_);
  and (_33397_, _33396_, _33392_);
  or (_33398_, _33397_, _33290_);
  and (_43742_, _33398_, _43100_);
  and (_33400_, _01321_, \oc8051_golden_model_1.IP [4]);
  and (_33401_, _13300_, \oc8051_golden_model_1.IP [4]);
  and (_33402_, _08336_, _07830_);
  or (_33403_, _33402_, _33401_);
  or (_33404_, _33403_, _06132_);
  and (_33405_, _13305_, \oc8051_golden_model_1.IP [4]);
  and (_33406_, _14942_, _08415_);
  or (_33407_, _33406_, _33405_);
  and (_33408_, _33407_, _06152_);
  and (_33410_, _14928_, _07830_);
  or (_33411_, _33410_, _33401_);
  or (_33412_, _33411_, _06161_);
  and (_33413_, _07830_, \oc8051_golden_model_1.ACC [4]);
  or (_33414_, _33413_, _33401_);
  and (_33415_, _33414_, _07056_);
  and (_33416_, _07057_, \oc8051_golden_model_1.IP [4]);
  or (_33417_, _33416_, _06160_);
  or (_33418_, _33417_, _33415_);
  and (_33419_, _33418_, _06157_);
  and (_33421_, _33419_, _33412_);
  and (_33422_, _14932_, _08415_);
  or (_33423_, _33422_, _33405_);
  and (_33424_, _33423_, _06156_);
  or (_33425_, _33424_, _06217_);
  or (_33426_, _33425_, _33421_);
  or (_33427_, _33403_, _07075_);
  and (_33428_, _33427_, _33426_);
  or (_33429_, _33428_, _06220_);
  or (_33430_, _33414_, _06229_);
  and (_33432_, _33430_, _06153_);
  and (_33433_, _33432_, _33429_);
  or (_33434_, _33433_, _33408_);
  and (_33435_, _33434_, _06146_);
  and (_33436_, _14950_, _08415_);
  or (_33437_, _33436_, _33405_);
  and (_33438_, _33437_, _06145_);
  or (_33439_, _33438_, _33435_);
  and (_33440_, _33439_, _06140_);
  and (_33441_, _14966_, _08415_);
  or (_33443_, _33441_, _33405_);
  and (_33444_, _33443_, _06139_);
  or (_33445_, _33444_, _09842_);
  or (_33446_, _33445_, _33440_);
  and (_33447_, _33446_, _33404_);
  or (_33448_, _33447_, _06116_);
  and (_33449_, _09209_, _07830_);
  or (_33450_, _33401_, _06117_);
  or (_33451_, _33450_, _33449_);
  and (_33452_, _33451_, _06114_);
  and (_33454_, _33452_, _33448_);
  and (_33455_, _15013_, _07830_);
  or (_33456_, _33455_, _33401_);
  and (_33457_, _33456_, _05787_);
  or (_33458_, _33457_, _11136_);
  or (_33459_, _33458_, _33454_);
  and (_33460_, _15029_, _07830_);
  or (_33461_, _33401_, _07127_);
  or (_33462_, _33461_, _33460_);
  and (_33463_, _08715_, _07830_);
  or (_33464_, _33463_, _33401_);
  or (_33465_, _33464_, _06111_);
  and (_33466_, _33465_, _07125_);
  and (_33467_, _33466_, _33462_);
  and (_33468_, _33467_, _33459_);
  and (_33469_, _10289_, _07830_);
  or (_33470_, _33469_, _33401_);
  and (_33471_, _33470_, _06402_);
  or (_33472_, _33471_, _33468_);
  and (_33473_, _33472_, _07132_);
  or (_33475_, _33401_, _08339_);
  and (_33476_, _33464_, _06306_);
  and (_33477_, _33476_, _33475_);
  or (_33478_, _33477_, _33473_);
  and (_33479_, _33478_, _07130_);
  and (_33480_, _33414_, _06411_);
  and (_33481_, _33480_, _33475_);
  or (_33482_, _33481_, _06303_);
  or (_33483_, _33482_, _33479_);
  and (_33484_, _15026_, _07830_);
  or (_33486_, _33401_, _08819_);
  or (_33487_, _33486_, _33484_);
  and (_33488_, _33487_, _08824_);
  and (_33489_, _33488_, _33483_);
  nor (_33490_, _10288_, _13300_);
  or (_33491_, _33490_, _33401_);
  and (_33492_, _33491_, _06396_);
  or (_33493_, _33492_, _06433_);
  or (_33494_, _33493_, _33489_);
  or (_33495_, _33411_, _06829_);
  and (_33497_, _33495_, _05749_);
  and (_33498_, _33497_, _33494_);
  and (_33499_, _33407_, _05748_);
  or (_33500_, _33499_, _06440_);
  or (_33501_, _33500_, _33498_);
  and (_33502_, _15087_, _07830_);
  or (_33503_, _33401_, _06444_);
  or (_33504_, _33503_, _33502_);
  and (_33505_, _33504_, _01317_);
  and (_33506_, _33505_, _33501_);
  or (_33508_, _33506_, _33400_);
  and (_43743_, _33508_, _43100_);
  and (_33509_, _01321_, \oc8051_golden_model_1.IP [5]);
  and (_33510_, _13300_, \oc8051_golden_model_1.IP [5]);
  and (_33511_, _15119_, _07830_);
  or (_33512_, _33511_, _33510_);
  or (_33513_, _33512_, _06161_);
  and (_33514_, _07830_, \oc8051_golden_model_1.ACC [5]);
  or (_33515_, _33514_, _33510_);
  and (_33516_, _33515_, _07056_);
  and (_33518_, _07057_, \oc8051_golden_model_1.IP [5]);
  or (_33519_, _33518_, _06160_);
  or (_33520_, _33519_, _33516_);
  and (_33521_, _33520_, _06157_);
  and (_33522_, _33521_, _33513_);
  and (_33523_, _13305_, \oc8051_golden_model_1.IP [5]);
  and (_33524_, _15123_, _08415_);
  or (_33525_, _33524_, _33523_);
  and (_33526_, _33525_, _06156_);
  or (_33527_, _33526_, _06217_);
  or (_33529_, _33527_, _33522_);
  and (_33530_, _08101_, _07830_);
  or (_33531_, _33530_, _33510_);
  or (_33532_, _33531_, _07075_);
  and (_33533_, _33532_, _33529_);
  or (_33534_, _33533_, _06220_);
  or (_33535_, _33515_, _06229_);
  and (_33536_, _33535_, _06153_);
  and (_33537_, _33536_, _33534_);
  and (_33538_, _15104_, _08415_);
  or (_33540_, _33538_, _33523_);
  and (_33541_, _33540_, _06152_);
  or (_33542_, _33541_, _06145_);
  or (_33543_, _33542_, _33537_);
  or (_33544_, _33523_, _15138_);
  and (_33545_, _33544_, _33525_);
  or (_33546_, _33545_, _06146_);
  and (_33547_, _33546_, _06140_);
  and (_33548_, _33547_, _33543_);
  and (_33549_, _15155_, _08415_);
  or (_33551_, _33549_, _33523_);
  and (_33552_, _33551_, _06139_);
  or (_33553_, _33552_, _09842_);
  or (_33554_, _33553_, _33548_);
  or (_33555_, _33531_, _06132_);
  and (_33556_, _33555_, _33554_);
  or (_33557_, _33556_, _06116_);
  and (_33558_, _09208_, _07830_);
  or (_33559_, _33510_, _06117_);
  or (_33560_, _33559_, _33558_);
  and (_33562_, _33560_, _06114_);
  and (_33563_, _33562_, _33557_);
  and (_33564_, _15203_, _07830_);
  or (_33565_, _33564_, _33510_);
  and (_33566_, _33565_, _05787_);
  or (_33567_, _33566_, _11136_);
  or (_33568_, _33567_, _33563_);
  and (_33569_, _15219_, _07830_);
  or (_33570_, _33510_, _07127_);
  or (_33571_, _33570_, _33569_);
  and (_33573_, _08736_, _07830_);
  or (_33574_, _33573_, _33510_);
  or (_33575_, _33574_, _06111_);
  and (_33576_, _33575_, _07125_);
  and (_33577_, _33576_, _33571_);
  and (_33578_, _33577_, _33568_);
  and (_33579_, _12325_, _07830_);
  or (_33580_, _33579_, _33510_);
  and (_33581_, _33580_, _06402_);
  or (_33582_, _33581_, _33578_);
  and (_33584_, _33582_, _07132_);
  or (_33585_, _33510_, _08104_);
  and (_33586_, _33574_, _06306_);
  and (_33587_, _33586_, _33585_);
  or (_33588_, _33587_, _33584_);
  and (_33589_, _33588_, _07130_);
  and (_33590_, _33515_, _06411_);
  and (_33591_, _33590_, _33585_);
  or (_33592_, _33591_, _06303_);
  or (_33593_, _33592_, _33589_);
  and (_33595_, _15216_, _07830_);
  or (_33596_, _33510_, _08819_);
  or (_33597_, _33596_, _33595_);
  and (_33598_, _33597_, _08824_);
  and (_33599_, _33598_, _33593_);
  nor (_33600_, _10269_, _13300_);
  or (_33601_, _33600_, _33510_);
  and (_33602_, _33601_, _06396_);
  or (_33603_, _33602_, _06433_);
  or (_33604_, _33603_, _33599_);
  or (_33606_, _33512_, _06829_);
  and (_33607_, _33606_, _05749_);
  and (_33608_, _33607_, _33604_);
  and (_33609_, _33540_, _05748_);
  or (_33610_, _33609_, _06440_);
  or (_33611_, _33610_, _33608_);
  and (_33612_, _15275_, _07830_);
  or (_33613_, _33510_, _06444_);
  or (_33614_, _33613_, _33612_);
  and (_33615_, _33614_, _01317_);
  and (_33617_, _33615_, _33611_);
  or (_33618_, _33617_, _33509_);
  and (_43744_, _33618_, _43100_);
  and (_33619_, _01321_, \oc8051_golden_model_1.IP [6]);
  and (_33620_, _13300_, \oc8051_golden_model_1.IP [6]);
  and (_33621_, _15300_, _07830_);
  or (_33622_, _33621_, _33620_);
  or (_33623_, _33622_, _06161_);
  and (_33624_, _07830_, \oc8051_golden_model_1.ACC [6]);
  or (_33625_, _33624_, _33620_);
  and (_33627_, _33625_, _07056_);
  and (_33628_, _07057_, \oc8051_golden_model_1.IP [6]);
  or (_33629_, _33628_, _06160_);
  or (_33630_, _33629_, _33627_);
  and (_33631_, _33630_, _06157_);
  and (_33632_, _33631_, _33623_);
  and (_33633_, _13305_, \oc8051_golden_model_1.IP [6]);
  and (_33634_, _15316_, _08415_);
  or (_33635_, _33634_, _33633_);
  and (_33636_, _33635_, _06156_);
  or (_33638_, _33636_, _06217_);
  or (_33639_, _33638_, _33632_);
  and (_33640_, _08012_, _07830_);
  or (_33641_, _33640_, _33620_);
  or (_33642_, _33641_, _07075_);
  and (_33643_, _33642_, _33639_);
  or (_33644_, _33643_, _06220_);
  or (_33645_, _33625_, _06229_);
  and (_33646_, _33645_, _06153_);
  and (_33647_, _33646_, _33644_);
  and (_33649_, _15297_, _08415_);
  or (_33650_, _33649_, _33633_);
  and (_33651_, _33650_, _06152_);
  or (_33652_, _33651_, _06145_);
  or (_33653_, _33652_, _33647_);
  or (_33654_, _33633_, _15331_);
  and (_33655_, _33654_, _33635_);
  or (_33656_, _33655_, _06146_);
  and (_33657_, _33656_, _06140_);
  and (_33658_, _33657_, _33653_);
  and (_33660_, _15348_, _08415_);
  or (_33661_, _33660_, _33633_);
  and (_33662_, _33661_, _06139_);
  or (_33663_, _33662_, _09842_);
  or (_33664_, _33663_, _33658_);
  or (_33665_, _33641_, _06132_);
  and (_33666_, _33665_, _33664_);
  or (_33667_, _33666_, _06116_);
  and (_33668_, _09207_, _07830_);
  or (_33669_, _33620_, _06117_);
  or (_33671_, _33669_, _33668_);
  and (_33672_, _33671_, _06114_);
  and (_33673_, _33672_, _33667_);
  and (_33674_, _15395_, _07830_);
  or (_33675_, _33674_, _33620_);
  and (_33676_, _33675_, _05787_);
  or (_33677_, _33676_, _11136_);
  or (_33678_, _33677_, _33673_);
  and (_33679_, _15413_, _07830_);
  or (_33680_, _33620_, _07127_);
  or (_33682_, _33680_, _33679_);
  and (_33683_, _15402_, _07830_);
  or (_33684_, _33683_, _33620_);
  or (_33685_, _33684_, _06111_);
  and (_33686_, _33685_, _07125_);
  and (_33687_, _33686_, _33682_);
  and (_33688_, _33687_, _33678_);
  and (_33689_, _10295_, _07830_);
  or (_33690_, _33689_, _33620_);
  and (_33691_, _33690_, _06402_);
  or (_33693_, _33691_, _33688_);
  and (_33694_, _33693_, _07132_);
  or (_33695_, _33620_, _08015_);
  and (_33696_, _33684_, _06306_);
  and (_33697_, _33696_, _33695_);
  or (_33698_, _33697_, _33694_);
  and (_33699_, _33698_, _07130_);
  and (_33700_, _33625_, _06411_);
  and (_33701_, _33700_, _33695_);
  or (_33702_, _33701_, _06303_);
  or (_33704_, _33702_, _33699_);
  and (_33705_, _15410_, _07830_);
  or (_33706_, _33620_, _08819_);
  or (_33707_, _33706_, _33705_);
  and (_33708_, _33707_, _08824_);
  and (_33709_, _33708_, _33704_);
  nor (_33710_, _10294_, _13300_);
  or (_33711_, _33710_, _33620_);
  and (_33712_, _33711_, _06396_);
  or (_33713_, _33712_, _06433_);
  or (_33715_, _33713_, _33709_);
  or (_33716_, _33622_, _06829_);
  and (_33717_, _33716_, _05749_);
  and (_33718_, _33717_, _33715_);
  and (_33719_, _33650_, _05748_);
  or (_33720_, _33719_, _06440_);
  or (_33721_, _33720_, _33718_);
  and (_33722_, _15478_, _07830_);
  or (_33723_, _33620_, _06444_);
  or (_33724_, _33723_, _33722_);
  and (_33726_, _33724_, _01317_);
  and (_33727_, _33726_, _33721_);
  or (_33728_, _33727_, _33619_);
  and (_43745_, _33728_, _43100_);
  not (_33729_, \oc8051_golden_model_1.IE [0]);
  nor (_33730_, _01317_, _33729_);
  nand (_33731_, _10276_, _07826_);
  nor (_33732_, _07826_, _33729_);
  nor (_33733_, _33732_, _07130_);
  nand (_33734_, _33733_, _33731_);
  and (_33736_, _07826_, _07049_);
  or (_33737_, _33736_, _33732_);
  or (_33738_, _33737_, _06132_);
  nor (_33739_, _08211_, _13402_);
  or (_33740_, _33739_, _33732_);
  or (_33741_, _33740_, _06161_);
  and (_33742_, _07826_, \oc8051_golden_model_1.ACC [0]);
  or (_33743_, _33742_, _33732_);
  and (_33744_, _33743_, _07056_);
  nor (_33745_, _07056_, _33729_);
  or (_33747_, _33745_, _06160_);
  or (_33748_, _33747_, _33744_);
  and (_33749_, _33748_, _06157_);
  and (_33750_, _33749_, _33741_);
  nor (_33751_, _08418_, _33729_);
  and (_33752_, _14169_, _08418_);
  or (_33753_, _33752_, _33751_);
  and (_33754_, _33753_, _06156_);
  or (_33755_, _33754_, _33750_);
  and (_33756_, _33755_, _07075_);
  and (_33758_, _33737_, _06217_);
  or (_33759_, _33758_, _06220_);
  or (_33760_, _33759_, _33756_);
  or (_33761_, _33743_, _06229_);
  and (_33762_, _33761_, _06153_);
  and (_33763_, _33762_, _33760_);
  and (_33764_, _33732_, _06152_);
  or (_33765_, _33764_, _06145_);
  or (_33766_, _33765_, _33763_);
  or (_33767_, _33740_, _06146_);
  and (_33769_, _33767_, _06140_);
  and (_33770_, _33769_, _33766_);
  or (_33771_, _33751_, _14170_);
  and (_33772_, _33771_, _06139_);
  and (_33773_, _33772_, _33753_);
  or (_33774_, _33773_, _09842_);
  or (_33775_, _33774_, _33770_);
  and (_33776_, _33775_, _33738_);
  or (_33777_, _33776_, _06116_);
  and (_33778_, _09160_, _07826_);
  or (_33780_, _33732_, _06117_);
  or (_33781_, _33780_, _33778_);
  and (_33782_, _33781_, _06114_);
  and (_33783_, _33782_, _33777_);
  and (_33784_, _14260_, _07826_);
  or (_33785_, _33784_, _33732_);
  and (_33786_, _33785_, _05787_);
  or (_33787_, _33786_, _33783_);
  or (_33788_, _33787_, _11136_);
  and (_33789_, _14275_, _07826_);
  or (_33791_, _33732_, _07127_);
  or (_33792_, _33791_, _33789_);
  and (_33793_, _07826_, _08708_);
  or (_33794_, _33793_, _33732_);
  or (_33795_, _33794_, _06111_);
  and (_33796_, _33795_, _07125_);
  and (_33797_, _33796_, _33792_);
  and (_33798_, _33797_, _33788_);
  nor (_33799_, _12321_, _13402_);
  or (_33800_, _33799_, _33732_);
  and (_33802_, _33731_, _06402_);
  and (_33803_, _33802_, _33800_);
  or (_33804_, _33803_, _33798_);
  and (_33805_, _33804_, _07132_);
  nand (_33806_, _33794_, _06306_);
  nor (_33807_, _33806_, _33739_);
  or (_33808_, _33807_, _06411_);
  or (_33809_, _33808_, _33805_);
  and (_33810_, _33809_, _33734_);
  or (_33811_, _33810_, _06303_);
  and (_33813_, _14167_, _07826_);
  or (_33814_, _33732_, _08819_);
  or (_33815_, _33814_, _33813_);
  and (_33816_, _33815_, _08824_);
  and (_33817_, _33816_, _33811_);
  and (_33818_, _33800_, _06396_);
  or (_33819_, _33818_, _06433_);
  or (_33820_, _33819_, _33817_);
  or (_33821_, _33740_, _06829_);
  and (_33822_, _33821_, _33820_);
  or (_33824_, _33822_, _05748_);
  or (_33825_, _33732_, _05749_);
  and (_33826_, _33825_, _33824_);
  or (_33827_, _33826_, _06440_);
  or (_33828_, _33740_, _06444_);
  and (_33829_, _33828_, _01317_);
  and (_33830_, _33829_, _33827_);
  or (_33831_, _33830_, _33730_);
  and (_43747_, _33831_, _43100_);
  not (_33832_, \oc8051_golden_model_1.IE [1]);
  nor (_33834_, _01317_, _33832_);
  nor (_33835_, _07826_, _33832_);
  nor (_33836_, _10277_, _13402_);
  or (_33837_, _33836_, _33835_);
  or (_33838_, _33837_, _08824_);
  and (_33839_, _07826_, _07306_);
  or (_33840_, _33839_, _33835_);
  or (_33841_, _33840_, _07075_);
  or (_33842_, _07826_, \oc8051_golden_model_1.IE [1]);
  and (_33843_, _14363_, _07826_);
  not (_33845_, _33843_);
  and (_33846_, _33845_, _33842_);
  or (_33847_, _33846_, _06161_);
  and (_33848_, _07826_, \oc8051_golden_model_1.ACC [1]);
  or (_33849_, _33848_, _33835_);
  and (_33850_, _33849_, _07056_);
  nor (_33851_, _07056_, _33832_);
  or (_33852_, _33851_, _06160_);
  or (_33853_, _33852_, _33850_);
  and (_33854_, _33853_, _06157_);
  and (_33856_, _33854_, _33847_);
  nor (_33857_, _08418_, _33832_);
  and (_33858_, _14367_, _08418_);
  or (_33859_, _33858_, _33857_);
  and (_33860_, _33859_, _06156_);
  or (_33861_, _33860_, _06217_);
  or (_33862_, _33861_, _33856_);
  and (_33863_, _33862_, _33841_);
  or (_33864_, _33863_, _06220_);
  or (_33865_, _33849_, _06229_);
  and (_33867_, _33865_, _06153_);
  and (_33868_, _33867_, _33864_);
  and (_33869_, _14349_, _08418_);
  or (_33870_, _33869_, _33857_);
  and (_33871_, _33870_, _06152_);
  or (_33872_, _33871_, _06145_);
  or (_33873_, _33872_, _33868_);
  and (_33874_, _33858_, _14382_);
  or (_33875_, _33857_, _06146_);
  or (_33876_, _33875_, _33874_);
  and (_33878_, _33876_, _33873_);
  and (_33879_, _33878_, _06140_);
  and (_33880_, _14351_, _08418_);
  or (_33881_, _33857_, _33880_);
  and (_33882_, _33881_, _06139_);
  or (_33883_, _33882_, _09842_);
  or (_33884_, _33883_, _33879_);
  or (_33885_, _33840_, _06132_);
  and (_33886_, _33885_, _33884_);
  or (_33887_, _33886_, _06116_);
  and (_33889_, _09115_, _07826_);
  or (_33890_, _33835_, _06117_);
  or (_33891_, _33890_, _33889_);
  and (_33892_, _33891_, _06114_);
  and (_33893_, _33892_, _33887_);
  and (_33894_, _14442_, _07826_);
  or (_33895_, _33894_, _33835_);
  and (_33896_, _33895_, _05787_);
  or (_33897_, _33896_, _33893_);
  and (_33898_, _33897_, _06298_);
  or (_33900_, _14346_, _13402_);
  and (_33901_, _33900_, _06297_);
  nand (_33902_, _07826_, _06945_);
  and (_33903_, _33902_, _06110_);
  or (_33904_, _33903_, _33901_);
  and (_33905_, _33904_, _33842_);
  or (_33906_, _33905_, _06402_);
  or (_33907_, _33906_, _33898_);
  nand (_33908_, _10275_, _07826_);
  and (_33909_, _33908_, _33837_);
  or (_33911_, _33909_, _07125_);
  and (_33912_, _33911_, _07132_);
  and (_33913_, _33912_, _33907_);
  or (_33914_, _14344_, _13402_);
  and (_33915_, _33842_, _06306_);
  and (_33916_, _33915_, _33914_);
  or (_33917_, _33916_, _06411_);
  or (_33918_, _33917_, _33913_);
  nor (_33919_, _33835_, _07130_);
  nand (_33920_, _33919_, _33908_);
  and (_33922_, _33920_, _08819_);
  and (_33923_, _33922_, _33918_);
  or (_33924_, _33902_, _08176_);
  and (_33925_, _33842_, _06303_);
  and (_33926_, _33925_, _33924_);
  or (_33927_, _33926_, _06396_);
  or (_33928_, _33927_, _33923_);
  and (_33929_, _33928_, _33838_);
  or (_33930_, _33929_, _06433_);
  or (_33931_, _33846_, _06829_);
  and (_33933_, _33931_, _05749_);
  and (_33934_, _33933_, _33930_);
  and (_33935_, _33870_, _05748_);
  or (_33936_, _33935_, _06440_);
  or (_33937_, _33936_, _33934_);
  or (_33938_, _33835_, _06444_);
  or (_33939_, _33938_, _33843_);
  and (_33940_, _33939_, _01317_);
  and (_33941_, _33940_, _33937_);
  or (_33942_, _33941_, _33834_);
  and (_43748_, _33942_, _43100_);
  and (_33944_, _01321_, \oc8051_golden_model_1.IE [2]);
  and (_33945_, _13402_, \oc8051_golden_model_1.IE [2]);
  and (_33946_, _07826_, _07708_);
  or (_33947_, _33946_, _33945_);
  or (_33948_, _33947_, _06132_);
  or (_33949_, _33947_, _07075_);
  and (_33950_, _14542_, _07826_);
  or (_33951_, _33950_, _33945_);
  or (_33952_, _33951_, _06161_);
  and (_33954_, _07826_, \oc8051_golden_model_1.ACC [2]);
  or (_33955_, _33954_, _33945_);
  and (_33956_, _33955_, _07056_);
  and (_33957_, _07057_, \oc8051_golden_model_1.IE [2]);
  or (_33958_, _33957_, _06160_);
  or (_33959_, _33958_, _33956_);
  and (_33960_, _33959_, _06157_);
  and (_33961_, _33960_, _33952_);
  and (_33962_, _13407_, \oc8051_golden_model_1.IE [2]);
  and (_33963_, _14538_, _08418_);
  or (_33965_, _33963_, _33962_);
  and (_33966_, _33965_, _06156_);
  or (_33967_, _33966_, _06217_);
  or (_33968_, _33967_, _33961_);
  and (_33969_, _33968_, _33949_);
  or (_33970_, _33969_, _06220_);
  or (_33971_, _33955_, _06229_);
  and (_33972_, _33971_, _06153_);
  and (_33973_, _33972_, _33970_);
  and (_33974_, _14536_, _08418_);
  or (_33976_, _33974_, _33962_);
  and (_33977_, _33976_, _06152_);
  or (_33978_, _33977_, _06145_);
  or (_33979_, _33978_, _33973_);
  and (_33980_, _33963_, _14569_);
  or (_33981_, _33962_, _06146_);
  or (_33982_, _33981_, _33980_);
  and (_33983_, _33982_, _06140_);
  and (_33984_, _33983_, _33979_);
  and (_33985_, _14583_, _08418_);
  or (_33987_, _33985_, _33962_);
  and (_33988_, _33987_, _06139_);
  or (_33989_, _33988_, _09842_);
  or (_33990_, _33989_, _33984_);
  and (_33991_, _33990_, _33948_);
  or (_33992_, _33991_, _06116_);
  and (_33993_, _09211_, _07826_);
  or (_33994_, _33945_, _06117_);
  or (_33995_, _33994_, _33993_);
  and (_33996_, _33995_, _06114_);
  and (_33998_, _33996_, _33992_);
  and (_33999_, _14630_, _07826_);
  or (_34000_, _33945_, _33999_);
  and (_34001_, _34000_, _05787_);
  or (_34002_, _34001_, _33998_);
  or (_34003_, _34002_, _11136_);
  and (_34004_, _14646_, _07826_);
  or (_34005_, _33945_, _07127_);
  or (_34006_, _34005_, _34004_);
  and (_34007_, _07826_, _08768_);
  or (_34009_, _34007_, _33945_);
  or (_34010_, _34009_, _06111_);
  and (_34011_, _34010_, _07125_);
  and (_34012_, _34011_, _34006_);
  and (_34013_, _34012_, _34003_);
  and (_34014_, _10282_, _07826_);
  or (_34015_, _34014_, _33945_);
  and (_34016_, _34015_, _06402_);
  or (_34017_, _34016_, _34013_);
  and (_34018_, _34017_, _07132_);
  or (_34020_, _33945_, _08248_);
  and (_34021_, _34009_, _06306_);
  and (_34022_, _34021_, _34020_);
  or (_34023_, _34022_, _34018_);
  and (_34024_, _34023_, _07130_);
  and (_34025_, _33955_, _06411_);
  and (_34026_, _34025_, _34020_);
  or (_34027_, _34026_, _06303_);
  or (_34028_, _34027_, _34024_);
  and (_34029_, _14643_, _07826_);
  or (_34031_, _33945_, _08819_);
  or (_34032_, _34031_, _34029_);
  and (_34033_, _34032_, _08824_);
  and (_34034_, _34033_, _34028_);
  nor (_34035_, _10281_, _13402_);
  or (_34036_, _34035_, _33945_);
  and (_34037_, _34036_, _06396_);
  or (_34038_, _34037_, _06433_);
  or (_34039_, _34038_, _34034_);
  or (_34040_, _33951_, _06829_);
  and (_34042_, _34040_, _05749_);
  and (_34043_, _34042_, _34039_);
  and (_34044_, _33976_, _05748_);
  or (_34045_, _34044_, _06440_);
  or (_34046_, _34045_, _34043_);
  and (_34047_, _14710_, _07826_);
  or (_34048_, _33945_, _06444_);
  or (_34049_, _34048_, _34047_);
  and (_34050_, _34049_, _01317_);
  and (_34051_, _34050_, _34046_);
  or (_34053_, _34051_, _33944_);
  and (_43749_, _34053_, _43100_);
  and (_34054_, _01321_, \oc8051_golden_model_1.IE [3]);
  and (_34055_, _13402_, \oc8051_golden_model_1.IE [3]);
  and (_34056_, _07826_, _07544_);
  or (_34057_, _34056_, _34055_);
  or (_34058_, _34057_, _06132_);
  and (_34059_, _14738_, _07826_);
  or (_34060_, _34059_, _34055_);
  or (_34061_, _34060_, _06161_);
  and (_34063_, _07826_, \oc8051_golden_model_1.ACC [3]);
  or (_34064_, _34063_, _34055_);
  and (_34065_, _34064_, _07056_);
  and (_34066_, _07057_, \oc8051_golden_model_1.IE [3]);
  or (_34067_, _34066_, _06160_);
  or (_34068_, _34067_, _34065_);
  and (_34069_, _34068_, _06157_);
  and (_34070_, _34069_, _34061_);
  and (_34071_, _13407_, \oc8051_golden_model_1.IE [3]);
  and (_34072_, _14735_, _08418_);
  or (_34074_, _34072_, _34071_);
  and (_34075_, _34074_, _06156_);
  or (_34076_, _34075_, _06217_);
  or (_34077_, _34076_, _34070_);
  or (_34078_, _34057_, _07075_);
  and (_34079_, _34078_, _34077_);
  or (_34080_, _34079_, _06220_);
  or (_34081_, _34064_, _06229_);
  and (_34082_, _34081_, _06153_);
  and (_34083_, _34082_, _34080_);
  and (_34085_, _14731_, _08418_);
  or (_34086_, _34085_, _34071_);
  and (_34087_, _34086_, _06152_);
  or (_34088_, _34087_, _06145_);
  or (_34089_, _34088_, _34083_);
  or (_34090_, _34071_, _14764_);
  and (_34091_, _34090_, _34074_);
  or (_34092_, _34091_, _06146_);
  and (_34093_, _34092_, _06140_);
  and (_34094_, _34093_, _34089_);
  and (_34096_, _14732_, _08418_);
  or (_34097_, _34096_, _34071_);
  and (_34098_, _34097_, _06139_);
  or (_34099_, _34098_, _09842_);
  or (_34100_, _34099_, _34094_);
  and (_34101_, _34100_, _34058_);
  or (_34102_, _34101_, _06116_);
  and (_34103_, _09210_, _07826_);
  or (_34104_, _34055_, _06117_);
  or (_34105_, _34104_, _34103_);
  and (_34107_, _34105_, _06114_);
  and (_34108_, _34107_, _34102_);
  and (_34109_, _14825_, _07826_);
  or (_34110_, _34055_, _34109_);
  and (_34111_, _34110_, _05787_);
  or (_34112_, _34111_, _34108_);
  or (_34113_, _34112_, _11136_);
  and (_34114_, _14727_, _07826_);
  or (_34115_, _34055_, _07127_);
  or (_34116_, _34115_, _34114_);
  and (_34118_, _07826_, _08712_);
  or (_34119_, _34118_, _34055_);
  or (_34120_, _34119_, _06111_);
  and (_34121_, _34120_, _07125_);
  and (_34122_, _34121_, _34116_);
  and (_34123_, _34122_, _34113_);
  and (_34124_, _12318_, _07826_);
  or (_34125_, _34124_, _34055_);
  and (_34126_, _34125_, _06402_);
  or (_34127_, _34126_, _34123_);
  and (_34129_, _34127_, _07132_);
  or (_34130_, _34055_, _08140_);
  and (_34131_, _34119_, _06306_);
  and (_34132_, _34131_, _34130_);
  or (_34133_, _34132_, _34129_);
  and (_34134_, _34133_, _07130_);
  and (_34135_, _34064_, _06411_);
  and (_34136_, _34135_, _34130_);
  or (_34137_, _34136_, _06303_);
  or (_34138_, _34137_, _34134_);
  and (_34140_, _14724_, _07826_);
  or (_34141_, _34055_, _08819_);
  or (_34142_, _34141_, _34140_);
  and (_34143_, _34142_, _08824_);
  and (_34144_, _34143_, _34138_);
  nor (_34145_, _10273_, _13402_);
  or (_34146_, _34145_, _34055_);
  and (_34147_, _34146_, _06396_);
  or (_34148_, _34147_, _06433_);
  or (_34149_, _34148_, _34144_);
  or (_34151_, _34060_, _06829_);
  and (_34152_, _34151_, _05749_);
  and (_34153_, _34152_, _34149_);
  and (_34154_, _34086_, _05748_);
  or (_34155_, _34154_, _06440_);
  or (_34156_, _34155_, _34153_);
  and (_34157_, _14897_, _07826_);
  or (_34158_, _34055_, _06444_);
  or (_34159_, _34158_, _34157_);
  and (_34160_, _34159_, _01317_);
  and (_34161_, _34160_, _34156_);
  or (_34162_, _34161_, _34054_);
  and (_43750_, _34162_, _43100_);
  and (_34163_, _01321_, \oc8051_golden_model_1.IE [4]);
  and (_34164_, _13402_, \oc8051_golden_model_1.IE [4]);
  and (_34165_, _08336_, _07826_);
  or (_34166_, _34165_, _34164_);
  or (_34167_, _34166_, _06132_);
  and (_34168_, _13407_, \oc8051_golden_model_1.IE [4]);
  and (_34169_, _14942_, _08418_);
  or (_34171_, _34169_, _34168_);
  and (_34172_, _34171_, _06152_);
  and (_34173_, _14928_, _07826_);
  or (_34174_, _34173_, _34164_);
  or (_34175_, _34174_, _06161_);
  and (_34176_, _07826_, \oc8051_golden_model_1.ACC [4]);
  or (_34177_, _34176_, _34164_);
  and (_34178_, _34177_, _07056_);
  and (_34179_, _07057_, \oc8051_golden_model_1.IE [4]);
  or (_34180_, _34179_, _06160_);
  or (_34182_, _34180_, _34178_);
  and (_34183_, _34182_, _06157_);
  and (_34184_, _34183_, _34175_);
  and (_34185_, _14932_, _08418_);
  or (_34186_, _34185_, _34168_);
  and (_34187_, _34186_, _06156_);
  or (_34188_, _34187_, _06217_);
  or (_34189_, _34188_, _34184_);
  or (_34190_, _34166_, _07075_);
  and (_34191_, _34190_, _34189_);
  or (_34193_, _34191_, _06220_);
  or (_34194_, _34177_, _06229_);
  and (_34195_, _34194_, _06153_);
  and (_34196_, _34195_, _34193_);
  or (_34197_, _34196_, _34172_);
  and (_34198_, _34197_, _06146_);
  and (_34199_, _14950_, _08418_);
  or (_34200_, _34199_, _34168_);
  and (_34201_, _34200_, _06145_);
  or (_34202_, _34201_, _34198_);
  and (_34204_, _34202_, _06140_);
  and (_34205_, _14966_, _08418_);
  or (_34206_, _34205_, _34168_);
  and (_34207_, _34206_, _06139_);
  or (_34208_, _34207_, _09842_);
  or (_34209_, _34208_, _34204_);
  and (_34210_, _34209_, _34167_);
  or (_34211_, _34210_, _06116_);
  and (_34212_, _09209_, _07826_);
  or (_34213_, _34164_, _06117_);
  or (_34215_, _34213_, _34212_);
  and (_34216_, _34215_, _06114_);
  and (_34217_, _34216_, _34211_);
  and (_34218_, _15013_, _07826_);
  or (_34219_, _34218_, _34164_);
  and (_34220_, _34219_, _05787_);
  or (_34221_, _34220_, _11136_);
  or (_34222_, _34221_, _34217_);
  and (_34223_, _15029_, _07826_);
  or (_34224_, _34164_, _07127_);
  or (_34226_, _34224_, _34223_);
  and (_34227_, _08715_, _07826_);
  or (_34228_, _34227_, _34164_);
  or (_34229_, _34228_, _06111_);
  and (_34230_, _34229_, _07125_);
  and (_34231_, _34230_, _34226_);
  and (_34232_, _34231_, _34222_);
  and (_34233_, _10289_, _07826_);
  or (_34234_, _34233_, _34164_);
  and (_34235_, _34234_, _06402_);
  or (_34237_, _34235_, _34232_);
  and (_34238_, _34237_, _07132_);
  or (_34239_, _34164_, _08339_);
  and (_34240_, _34228_, _06306_);
  and (_34241_, _34240_, _34239_);
  or (_34242_, _34241_, _34238_);
  and (_34243_, _34242_, _07130_);
  and (_34244_, _34177_, _06411_);
  and (_34245_, _34244_, _34239_);
  or (_34246_, _34245_, _06303_);
  or (_34248_, _34246_, _34243_);
  and (_34249_, _15026_, _07826_);
  or (_34250_, _34164_, _08819_);
  or (_34251_, _34250_, _34249_);
  and (_34252_, _34251_, _08824_);
  and (_34253_, _34252_, _34248_);
  nor (_34254_, _10288_, _13402_);
  or (_34255_, _34254_, _34164_);
  and (_34256_, _34255_, _06396_);
  or (_34257_, _34256_, _06433_);
  or (_34259_, _34257_, _34253_);
  or (_34260_, _34174_, _06829_);
  and (_34261_, _34260_, _05749_);
  and (_34262_, _34261_, _34259_);
  and (_34263_, _34171_, _05748_);
  or (_34264_, _34263_, _06440_);
  or (_34265_, _34264_, _34262_);
  and (_34266_, _15087_, _07826_);
  or (_34267_, _34164_, _06444_);
  or (_34268_, _34267_, _34266_);
  and (_34270_, _34268_, _01317_);
  and (_34271_, _34270_, _34265_);
  or (_34272_, _34271_, _34163_);
  and (_43751_, _34272_, _43100_);
  and (_34273_, _01321_, \oc8051_golden_model_1.IE [5]);
  and (_34274_, _13402_, \oc8051_golden_model_1.IE [5]);
  and (_34275_, _15119_, _07826_);
  or (_34276_, _34275_, _34274_);
  or (_34278_, _34276_, _06161_);
  and (_34280_, _07826_, \oc8051_golden_model_1.ACC [5]);
  or (_34283_, _34280_, _34274_);
  and (_34285_, _34283_, _07056_);
  and (_34287_, _07057_, \oc8051_golden_model_1.IE [5]);
  or (_34289_, _34287_, _06160_);
  or (_34291_, _34289_, _34285_);
  and (_34293_, _34291_, _06157_);
  and (_34295_, _34293_, _34278_);
  and (_34297_, _13407_, \oc8051_golden_model_1.IE [5]);
  and (_34298_, _15123_, _08418_);
  or (_34299_, _34298_, _34297_);
  and (_34301_, _34299_, _06156_);
  or (_34302_, _34301_, _06217_);
  or (_34303_, _34302_, _34295_);
  and (_34304_, _08101_, _07826_);
  or (_34305_, _34304_, _34274_);
  or (_34306_, _34305_, _07075_);
  and (_34307_, _34306_, _34303_);
  or (_34308_, _34307_, _06220_);
  or (_34309_, _34283_, _06229_);
  and (_34310_, _34309_, _06153_);
  and (_34312_, _34310_, _34308_);
  and (_34313_, _15104_, _08418_);
  or (_34314_, _34313_, _34297_);
  and (_34315_, _34314_, _06152_);
  or (_34316_, _34315_, _06145_);
  or (_34317_, _34316_, _34312_);
  or (_34318_, _34297_, _15138_);
  and (_34319_, _34318_, _34299_);
  or (_34320_, _34319_, _06146_);
  and (_34321_, _34320_, _06140_);
  and (_34323_, _34321_, _34317_);
  and (_34324_, _15155_, _08418_);
  or (_34325_, _34324_, _34297_);
  and (_34326_, _34325_, _06139_);
  or (_34327_, _34326_, _09842_);
  or (_34328_, _34327_, _34323_);
  or (_34329_, _34305_, _06132_);
  and (_34330_, _34329_, _34328_);
  or (_34331_, _34330_, _06116_);
  and (_34332_, _09208_, _07826_);
  or (_34334_, _34274_, _06117_);
  or (_34335_, _34334_, _34332_);
  and (_34336_, _34335_, _06114_);
  and (_34337_, _34336_, _34331_);
  and (_34338_, _15203_, _07826_);
  or (_34339_, _34338_, _34274_);
  and (_34340_, _34339_, _05787_);
  or (_34341_, _34340_, _11136_);
  or (_34342_, _34341_, _34337_);
  and (_34343_, _15219_, _07826_);
  or (_34345_, _34274_, _07127_);
  or (_34346_, _34345_, _34343_);
  and (_34347_, _08736_, _07826_);
  or (_34348_, _34347_, _34274_);
  or (_34349_, _34348_, _06111_);
  and (_34350_, _34349_, _07125_);
  and (_34351_, _34350_, _34346_);
  and (_34352_, _34351_, _34342_);
  and (_34353_, _12325_, _07826_);
  or (_34354_, _34353_, _34274_);
  and (_34356_, _34354_, _06402_);
  or (_34357_, _34356_, _34352_);
  and (_34358_, _34357_, _07132_);
  or (_34359_, _34274_, _08104_);
  and (_34360_, _34348_, _06306_);
  and (_34361_, _34360_, _34359_);
  or (_34362_, _34361_, _34358_);
  and (_34363_, _34362_, _07130_);
  and (_34364_, _34283_, _06411_);
  and (_34365_, _34364_, _34359_);
  or (_34367_, _34365_, _06303_);
  or (_34368_, _34367_, _34363_);
  and (_34369_, _15216_, _07826_);
  or (_34370_, _34274_, _08819_);
  or (_34371_, _34370_, _34369_);
  and (_34372_, _34371_, _08824_);
  and (_34373_, _34372_, _34368_);
  nor (_34374_, _10269_, _13402_);
  or (_34375_, _34374_, _34274_);
  and (_34376_, _34375_, _06396_);
  or (_34378_, _34376_, _06433_);
  or (_34379_, _34378_, _34373_);
  or (_34380_, _34276_, _06829_);
  and (_34381_, _34380_, _05749_);
  and (_34382_, _34381_, _34379_);
  and (_34383_, _34314_, _05748_);
  or (_34384_, _34383_, _06440_);
  or (_34385_, _34384_, _34382_);
  and (_34386_, _15275_, _07826_);
  or (_34387_, _34274_, _06444_);
  or (_34389_, _34387_, _34386_);
  and (_34390_, _34389_, _01317_);
  and (_34391_, _34390_, _34385_);
  or (_34392_, _34391_, _34273_);
  and (_43752_, _34392_, _43100_);
  and (_34393_, _01321_, \oc8051_golden_model_1.IE [6]);
  and (_34394_, _13402_, \oc8051_golden_model_1.IE [6]);
  and (_34395_, _15300_, _07826_);
  or (_34396_, _34395_, _34394_);
  or (_34397_, _34396_, _06161_);
  and (_34399_, _07826_, \oc8051_golden_model_1.ACC [6]);
  or (_34400_, _34399_, _34394_);
  and (_34401_, _34400_, _07056_);
  and (_34402_, _07057_, \oc8051_golden_model_1.IE [6]);
  or (_34403_, _34402_, _06160_);
  or (_34404_, _34403_, _34401_);
  and (_34405_, _34404_, _06157_);
  and (_34406_, _34405_, _34397_);
  and (_34407_, _13407_, \oc8051_golden_model_1.IE [6]);
  and (_34408_, _15316_, _08418_);
  or (_34410_, _34408_, _34407_);
  and (_34411_, _34410_, _06156_);
  or (_34412_, _34411_, _06217_);
  or (_34413_, _34412_, _34406_);
  and (_34414_, _08012_, _07826_);
  or (_34415_, _34414_, _34394_);
  or (_34416_, _34415_, _07075_);
  and (_34417_, _34416_, _34413_);
  or (_34418_, _34417_, _06220_);
  or (_34419_, _34400_, _06229_);
  and (_34421_, _34419_, _06153_);
  and (_34422_, _34421_, _34418_);
  and (_34423_, _15297_, _08418_);
  or (_34424_, _34423_, _34407_);
  and (_34425_, _34424_, _06152_);
  or (_34426_, _34425_, _06145_);
  or (_34427_, _34426_, _34422_);
  or (_34428_, _34407_, _15331_);
  and (_34429_, _34428_, _34410_);
  or (_34430_, _34429_, _06146_);
  and (_34432_, _34430_, _06140_);
  and (_34433_, _34432_, _34427_);
  and (_34434_, _15348_, _08418_);
  or (_34435_, _34434_, _34407_);
  and (_34436_, _34435_, _06139_);
  or (_34437_, _34436_, _09842_);
  or (_34438_, _34437_, _34433_);
  or (_34439_, _34415_, _06132_);
  and (_34440_, _34439_, _34438_);
  or (_34441_, _34440_, _06116_);
  and (_34443_, _09207_, _07826_);
  or (_34444_, _34394_, _06117_);
  or (_34445_, _34444_, _34443_);
  and (_34446_, _34445_, _06114_);
  and (_34447_, _34446_, _34441_);
  and (_34448_, _15395_, _07826_);
  or (_34449_, _34448_, _34394_);
  and (_34450_, _34449_, _05787_);
  or (_34451_, _34450_, _11136_);
  or (_34452_, _34451_, _34447_);
  and (_34454_, _15413_, _07826_);
  or (_34455_, _34394_, _07127_);
  or (_34456_, _34455_, _34454_);
  and (_34457_, _15402_, _07826_);
  or (_34458_, _34457_, _34394_);
  or (_34459_, _34458_, _06111_);
  and (_34460_, _34459_, _07125_);
  and (_34461_, _34460_, _34456_);
  and (_34462_, _34461_, _34452_);
  and (_34463_, _10295_, _07826_);
  or (_34465_, _34463_, _34394_);
  and (_34466_, _34465_, _06402_);
  or (_34467_, _34466_, _34462_);
  and (_34468_, _34467_, _07132_);
  or (_34469_, _34394_, _08015_);
  and (_34470_, _34458_, _06306_);
  and (_34471_, _34470_, _34469_);
  or (_34472_, _34471_, _34468_);
  and (_34473_, _34472_, _07130_);
  and (_34474_, _34400_, _06411_);
  and (_34476_, _34474_, _34469_);
  or (_34477_, _34476_, _06303_);
  or (_34478_, _34477_, _34473_);
  and (_34479_, _15410_, _07826_);
  or (_34480_, _34394_, _08819_);
  or (_34481_, _34480_, _34479_);
  and (_34482_, _34481_, _08824_);
  and (_34483_, _34482_, _34478_);
  nor (_34484_, _10294_, _13402_);
  or (_34485_, _34484_, _34394_);
  and (_34487_, _34485_, _06396_);
  or (_34488_, _34487_, _06433_);
  or (_34489_, _34488_, _34483_);
  or (_34490_, _34396_, _06829_);
  and (_34491_, _34490_, _05749_);
  and (_34492_, _34491_, _34489_);
  and (_34493_, _34424_, _05748_);
  or (_34494_, _34493_, _06440_);
  or (_34495_, _34494_, _34492_);
  and (_34496_, _15478_, _07826_);
  or (_34498_, _34394_, _06444_);
  or (_34499_, _34498_, _34496_);
  and (_34500_, _34499_, _01317_);
  and (_34501_, _34500_, _34495_);
  or (_34502_, _34501_, _34393_);
  and (_43753_, _34502_, _43100_);
  not (_34503_, \oc8051_golden_model_1.SCON [0]);
  nor (_34504_, _01317_, _34503_);
  nor (_34505_, _07778_, _34503_);
  and (_34506_, _07778_, _07049_);
  or (_34508_, _34506_, _34505_);
  or (_34509_, _34508_, _06132_);
  nor (_34510_, _08211_, _13504_);
  or (_34511_, _34510_, _34505_);
  or (_34512_, _34511_, _06161_);
  and (_34513_, _07778_, \oc8051_golden_model_1.ACC [0]);
  or (_34514_, _34513_, _34505_);
  and (_34515_, _34514_, _07056_);
  nor (_34516_, _07056_, _34503_);
  or (_34517_, _34516_, _06160_);
  or (_34519_, _34517_, _34515_);
  and (_34520_, _34519_, _06157_);
  and (_34521_, _34520_, _34512_);
  nor (_34522_, _08413_, _34503_);
  and (_34523_, _14169_, _08413_);
  or (_34524_, _34523_, _34522_);
  and (_34525_, _34524_, _06156_);
  or (_34526_, _34525_, _34521_);
  and (_34527_, _34526_, _07075_);
  and (_34528_, _34508_, _06217_);
  or (_34530_, _34528_, _06220_);
  or (_34531_, _34530_, _34527_);
  or (_34532_, _34514_, _06229_);
  and (_34533_, _34532_, _06153_);
  and (_34534_, _34533_, _34531_);
  and (_34535_, _34505_, _06152_);
  or (_34536_, _34535_, _06145_);
  or (_34537_, _34536_, _34534_);
  or (_34538_, _34511_, _06146_);
  and (_34539_, _34538_, _06140_);
  and (_34541_, _34539_, _34537_);
  or (_34542_, _34522_, _14170_);
  and (_34543_, _34542_, _06139_);
  and (_34544_, _34543_, _34524_);
  or (_34545_, _34544_, _09842_);
  or (_34546_, _34545_, _34541_);
  and (_34547_, _34546_, _34509_);
  or (_34548_, _34547_, _06116_);
  and (_34549_, _09160_, _07778_);
  or (_34550_, _34505_, _06117_);
  or (_34552_, _34550_, _34549_);
  and (_34553_, _34552_, _06114_);
  and (_34554_, _34553_, _34548_);
  and (_34555_, _14260_, _07778_);
  or (_34556_, _34555_, _34505_);
  and (_34557_, _34556_, _05787_);
  or (_34558_, _34557_, _34554_);
  or (_34559_, _34558_, _11136_);
  and (_34560_, _14275_, _07778_);
  or (_34561_, _34505_, _07127_);
  or (_34563_, _34561_, _34560_);
  and (_34564_, _07778_, _08708_);
  or (_34565_, _34564_, _34505_);
  or (_34566_, _34565_, _06111_);
  and (_34567_, _34566_, _07125_);
  and (_34568_, _34567_, _34563_);
  and (_34569_, _34568_, _34559_);
  nor (_34570_, _12321_, _13504_);
  or (_34571_, _34570_, _34505_);
  nand (_34572_, _10276_, _07778_);
  and (_34574_, _34572_, _06402_);
  and (_34575_, _34574_, _34571_);
  or (_34576_, _34575_, _34569_);
  and (_34577_, _34576_, _07132_);
  nand (_34578_, _34565_, _06306_);
  nor (_34579_, _34578_, _34510_);
  or (_34580_, _34579_, _06411_);
  or (_34581_, _34580_, _34577_);
  nor (_34582_, _34505_, _07130_);
  nand (_34583_, _34582_, _34572_);
  and (_34585_, _34583_, _34581_);
  or (_34586_, _34585_, _06303_);
  and (_34587_, _14167_, _07778_);
  or (_34588_, _34505_, _08819_);
  or (_34589_, _34588_, _34587_);
  and (_34590_, _34589_, _08824_);
  and (_34591_, _34590_, _34586_);
  and (_34592_, _34571_, _06396_);
  or (_34593_, _34592_, _06433_);
  or (_34594_, _34593_, _34591_);
  or (_34596_, _34511_, _06829_);
  and (_34597_, _34596_, _34594_);
  or (_34598_, _34597_, _05748_);
  or (_34599_, _34505_, _05749_);
  and (_34600_, _34599_, _34598_);
  or (_34601_, _34600_, _06440_);
  or (_34602_, _34511_, _06444_);
  and (_34603_, _34602_, _01317_);
  and (_34604_, _34603_, _34601_);
  or (_34605_, _34604_, _34504_);
  and (_43755_, _34605_, _43100_);
  not (_34607_, \oc8051_golden_model_1.SCON [1]);
  nor (_34608_, _01317_, _34607_);
  nor (_34609_, _07778_, _34607_);
  and (_34610_, _07778_, _07306_);
  or (_34611_, _34610_, _34609_);
  or (_34612_, _34611_, _07075_);
  or (_34613_, _07778_, \oc8051_golden_model_1.SCON [1]);
  and (_34614_, _14363_, _07778_);
  not (_34615_, _34614_);
  and (_34617_, _34615_, _34613_);
  or (_34618_, _34617_, _06161_);
  and (_34619_, _07778_, \oc8051_golden_model_1.ACC [1]);
  or (_34620_, _34619_, _34609_);
  and (_34621_, _34620_, _07056_);
  nor (_34622_, _07056_, _34607_);
  or (_34623_, _34622_, _06160_);
  or (_34624_, _34623_, _34621_);
  and (_34625_, _34624_, _06157_);
  and (_34626_, _34625_, _34618_);
  nor (_34628_, _08413_, _34607_);
  and (_34629_, _14367_, _08413_);
  or (_34630_, _34629_, _34628_);
  and (_34631_, _34630_, _06156_);
  or (_34632_, _34631_, _06217_);
  or (_34633_, _34632_, _34626_);
  and (_34634_, _34633_, _34612_);
  or (_34635_, _34634_, _06220_);
  or (_34636_, _34620_, _06229_);
  and (_34637_, _34636_, _06153_);
  and (_34639_, _34637_, _34635_);
  and (_34640_, _14349_, _08413_);
  or (_34641_, _34640_, _34628_);
  and (_34642_, _34641_, _06152_);
  or (_34643_, _34642_, _06145_);
  or (_34644_, _34643_, _34639_);
  and (_34645_, _34629_, _14382_);
  or (_34646_, _34628_, _06146_);
  or (_34647_, _34646_, _34645_);
  and (_34648_, _34647_, _34644_);
  and (_34650_, _34648_, _06140_);
  and (_34651_, _14351_, _08413_);
  or (_34652_, _34628_, _34651_);
  and (_34653_, _34652_, _06139_);
  or (_34654_, _34653_, _09842_);
  or (_34655_, _34654_, _34650_);
  or (_34656_, _34611_, _06132_);
  and (_34657_, _34656_, _34655_);
  or (_34658_, _34657_, _06116_);
  and (_34659_, _09115_, _07778_);
  or (_34661_, _34609_, _06117_);
  or (_34662_, _34661_, _34659_);
  and (_34663_, _34662_, _06114_);
  and (_34664_, _34663_, _34658_);
  and (_34665_, _14442_, _07778_);
  or (_34666_, _34665_, _34609_);
  and (_34667_, _34666_, _05787_);
  or (_34668_, _34667_, _34664_);
  and (_34669_, _34668_, _06298_);
  or (_34670_, _14346_, _13504_);
  and (_34672_, _34613_, _06297_);
  and (_34673_, _34672_, _34670_);
  nand (_34674_, _07778_, _06945_);
  and (_34675_, _34674_, _06110_);
  and (_34676_, _34675_, _34613_);
  or (_34677_, _34676_, _06402_);
  or (_34678_, _34677_, _34673_);
  or (_34679_, _34678_, _34669_);
  nor (_34680_, _10277_, _13504_);
  or (_34681_, _34680_, _34609_);
  nand (_34683_, _10275_, _07778_);
  and (_34684_, _34683_, _34681_);
  or (_34685_, _34684_, _07125_);
  and (_34686_, _34685_, _07132_);
  and (_34687_, _34686_, _34679_);
  or (_34688_, _14344_, _13504_);
  and (_34689_, _34613_, _06306_);
  and (_34690_, _34689_, _34688_);
  or (_34691_, _34690_, _06411_);
  or (_34692_, _34691_, _34687_);
  nor (_34694_, _34609_, _07130_);
  nand (_34695_, _34694_, _34683_);
  and (_34696_, _34695_, _08819_);
  and (_34697_, _34696_, _34692_);
  or (_34698_, _34674_, _08176_);
  and (_34699_, _34613_, _06303_);
  and (_34700_, _34699_, _34698_);
  or (_34701_, _34700_, _06396_);
  or (_34702_, _34701_, _34697_);
  or (_34703_, _34681_, _08824_);
  and (_34705_, _34703_, _34702_);
  or (_34706_, _34705_, _06433_);
  or (_34707_, _34617_, _06829_);
  and (_34708_, _34707_, _05749_);
  and (_34709_, _34708_, _34706_);
  and (_34710_, _34641_, _05748_);
  or (_34711_, _34710_, _06440_);
  or (_34712_, _34711_, _34709_);
  or (_34713_, _34609_, _06444_);
  or (_34714_, _34713_, _34614_);
  and (_34716_, _34714_, _01317_);
  and (_34717_, _34716_, _34712_);
  or (_34718_, _34717_, _34608_);
  and (_43756_, _34718_, _43100_);
  and (_34719_, _01321_, \oc8051_golden_model_1.SCON [2]);
  and (_34720_, _13504_, \oc8051_golden_model_1.SCON [2]);
  and (_34721_, _07778_, _07708_);
  or (_34722_, _34721_, _34720_);
  or (_34723_, _34722_, _06132_);
  or (_34724_, _34722_, _07075_);
  and (_34726_, _14542_, _07778_);
  or (_34727_, _34726_, _34720_);
  or (_34728_, _34727_, _06161_);
  and (_34729_, _07778_, \oc8051_golden_model_1.ACC [2]);
  or (_34730_, _34729_, _34720_);
  and (_34731_, _34730_, _07056_);
  and (_34732_, _07057_, \oc8051_golden_model_1.SCON [2]);
  or (_34733_, _34732_, _06160_);
  or (_34734_, _34733_, _34731_);
  and (_34735_, _34734_, _06157_);
  and (_34737_, _34735_, _34728_);
  and (_34738_, _13509_, \oc8051_golden_model_1.SCON [2]);
  and (_34739_, _14538_, _08413_);
  or (_34740_, _34739_, _34738_);
  and (_34741_, _34740_, _06156_);
  or (_34742_, _34741_, _06217_);
  or (_34743_, _34742_, _34737_);
  and (_34744_, _34743_, _34724_);
  or (_34745_, _34744_, _06220_);
  or (_34746_, _34730_, _06229_);
  and (_34748_, _34746_, _06153_);
  and (_34749_, _34748_, _34745_);
  and (_34750_, _14536_, _08413_);
  or (_34751_, _34750_, _34738_);
  and (_34752_, _34751_, _06152_);
  or (_34753_, _34752_, _06145_);
  or (_34754_, _34753_, _34749_);
  and (_34755_, _34739_, _14569_);
  or (_34756_, _34738_, _06146_);
  or (_34757_, _34756_, _34755_);
  and (_34759_, _34757_, _06140_);
  and (_34760_, _34759_, _34754_);
  and (_34761_, _14583_, _08413_);
  or (_34762_, _34761_, _34738_);
  and (_34763_, _34762_, _06139_);
  or (_34764_, _34763_, _09842_);
  or (_34765_, _34764_, _34760_);
  and (_34766_, _34765_, _34723_);
  or (_34767_, _34766_, _06116_);
  and (_34768_, _09211_, _07778_);
  or (_34770_, _34720_, _06117_);
  or (_34771_, _34770_, _34768_);
  and (_34772_, _34771_, _06114_);
  and (_34773_, _34772_, _34767_);
  and (_34774_, _14630_, _07778_);
  or (_34775_, _34720_, _34774_);
  and (_34776_, _34775_, _05787_);
  or (_34777_, _34776_, _34773_);
  or (_34778_, _34777_, _11136_);
  and (_34779_, _14646_, _07778_);
  or (_34781_, _34720_, _07127_);
  or (_34782_, _34781_, _34779_);
  and (_34783_, _07778_, _08768_);
  or (_34784_, _34783_, _34720_);
  or (_34785_, _34784_, _06111_);
  and (_34786_, _34785_, _07125_);
  and (_34787_, _34786_, _34782_);
  and (_34788_, _34787_, _34778_);
  and (_34789_, _10282_, _07778_);
  or (_34790_, _34789_, _34720_);
  and (_34792_, _34790_, _06402_);
  or (_34793_, _34792_, _34788_);
  and (_34794_, _34793_, _07132_);
  or (_34795_, _34720_, _08248_);
  and (_34796_, _34784_, _06306_);
  and (_34797_, _34796_, _34795_);
  or (_34798_, _34797_, _34794_);
  and (_34799_, _34798_, _07130_);
  and (_34800_, _34730_, _06411_);
  and (_34801_, _34800_, _34795_);
  or (_34803_, _34801_, _06303_);
  or (_34804_, _34803_, _34799_);
  and (_34805_, _14643_, _07778_);
  or (_34806_, _34720_, _08819_);
  or (_34807_, _34806_, _34805_);
  and (_34808_, _34807_, _08824_);
  and (_34809_, _34808_, _34804_);
  nor (_34810_, _10281_, _13504_);
  or (_34811_, _34810_, _34720_);
  and (_34812_, _34811_, _06396_);
  or (_34814_, _34812_, _06433_);
  or (_34815_, _34814_, _34809_);
  or (_34816_, _34727_, _06829_);
  and (_34817_, _34816_, _05749_);
  and (_34818_, _34817_, _34815_);
  and (_34819_, _34751_, _05748_);
  or (_34820_, _34819_, _06440_);
  or (_34821_, _34820_, _34818_);
  and (_34822_, _14710_, _07778_);
  or (_34823_, _34720_, _06444_);
  or (_34825_, _34823_, _34822_);
  and (_34826_, _34825_, _01317_);
  and (_34827_, _34826_, _34821_);
  or (_34828_, _34827_, _34719_);
  and (_43757_, _34828_, _43100_);
  and (_34829_, _01321_, \oc8051_golden_model_1.SCON [3]);
  and (_34830_, _13504_, \oc8051_golden_model_1.SCON [3]);
  and (_34831_, _07778_, _07544_);
  or (_34832_, _34831_, _34830_);
  or (_34833_, _34832_, _06132_);
  and (_34835_, _14738_, _07778_);
  or (_34836_, _34835_, _34830_);
  or (_34837_, _34836_, _06161_);
  and (_34838_, _07778_, \oc8051_golden_model_1.ACC [3]);
  or (_34839_, _34838_, _34830_);
  and (_34840_, _34839_, _07056_);
  and (_34841_, _07057_, \oc8051_golden_model_1.SCON [3]);
  or (_34842_, _34841_, _06160_);
  or (_34843_, _34842_, _34840_);
  and (_34844_, _34843_, _06157_);
  and (_34846_, _34844_, _34837_);
  and (_34847_, _13509_, \oc8051_golden_model_1.SCON [3]);
  and (_34848_, _14735_, _08413_);
  or (_34849_, _34848_, _34847_);
  and (_34850_, _34849_, _06156_);
  or (_34851_, _34850_, _06217_);
  or (_34852_, _34851_, _34846_);
  or (_34853_, _34832_, _07075_);
  and (_34854_, _34853_, _34852_);
  or (_34855_, _34854_, _06220_);
  or (_34857_, _34839_, _06229_);
  and (_34858_, _34857_, _06153_);
  and (_34859_, _34858_, _34855_);
  and (_34860_, _14731_, _08413_);
  or (_34861_, _34860_, _34847_);
  and (_34862_, _34861_, _06152_);
  or (_34863_, _34862_, _06145_);
  or (_34864_, _34863_, _34859_);
  or (_34865_, _34847_, _14764_);
  and (_34866_, _34865_, _34849_);
  or (_34868_, _34866_, _06146_);
  and (_34869_, _34868_, _06140_);
  and (_34870_, _34869_, _34864_);
  and (_34871_, _14732_, _08413_);
  or (_34872_, _34871_, _34847_);
  and (_34873_, _34872_, _06139_);
  or (_34874_, _34873_, _09842_);
  or (_34875_, _34874_, _34870_);
  and (_34876_, _34875_, _34833_);
  or (_34877_, _34876_, _06116_);
  and (_34879_, _09210_, _07778_);
  or (_34880_, _34830_, _06117_);
  or (_34881_, _34880_, _34879_);
  and (_34882_, _34881_, _06114_);
  and (_34883_, _34882_, _34877_);
  and (_34884_, _14825_, _07778_);
  or (_34885_, _34830_, _34884_);
  and (_34886_, _34885_, _05787_);
  or (_34887_, _34886_, _34883_);
  or (_34888_, _34887_, _11136_);
  and (_34890_, _14727_, _07778_);
  or (_34891_, _34830_, _07127_);
  or (_34892_, _34891_, _34890_);
  and (_34893_, _07778_, _08712_);
  or (_34894_, _34893_, _34830_);
  or (_34895_, _34894_, _06111_);
  and (_34896_, _34895_, _07125_);
  and (_34897_, _34896_, _34892_);
  and (_34898_, _34897_, _34888_);
  and (_34899_, _12318_, _07778_);
  or (_34901_, _34899_, _34830_);
  and (_34902_, _34901_, _06402_);
  or (_34903_, _34902_, _34898_);
  and (_34904_, _34903_, _07132_);
  or (_34905_, _34830_, _08140_);
  and (_34906_, _34894_, _06306_);
  and (_34907_, _34906_, _34905_);
  or (_34908_, _34907_, _34904_);
  and (_34909_, _34908_, _07130_);
  and (_34910_, _34839_, _06411_);
  and (_34912_, _34910_, _34905_);
  or (_34913_, _34912_, _06303_);
  or (_34914_, _34913_, _34909_);
  and (_34915_, _14724_, _07778_);
  or (_34916_, _34830_, _08819_);
  or (_34917_, _34916_, _34915_);
  and (_34918_, _34917_, _08824_);
  and (_34919_, _34918_, _34914_);
  nor (_34920_, _10273_, _13504_);
  or (_34921_, _34920_, _34830_);
  and (_34923_, _34921_, _06396_);
  or (_34924_, _34923_, _06433_);
  or (_34925_, _34924_, _34919_);
  or (_34926_, _34836_, _06829_);
  and (_34927_, _34926_, _05749_);
  and (_34928_, _34927_, _34925_);
  and (_34929_, _34861_, _05748_);
  or (_34930_, _34929_, _06440_);
  or (_34931_, _34930_, _34928_);
  and (_34932_, _14897_, _07778_);
  or (_34933_, _34830_, _06444_);
  or (_34934_, _34933_, _34932_);
  and (_34935_, _34934_, _01317_);
  and (_34936_, _34935_, _34931_);
  or (_34937_, _34936_, _34829_);
  and (_43758_, _34937_, _43100_);
  and (_34938_, _01321_, \oc8051_golden_model_1.SCON [4]);
  and (_34939_, _13504_, \oc8051_golden_model_1.SCON [4]);
  and (_34940_, _08336_, _07778_);
  or (_34941_, _34940_, _34939_);
  or (_34943_, _34941_, _06132_);
  and (_34944_, _13509_, \oc8051_golden_model_1.SCON [4]);
  and (_34945_, _14942_, _08413_);
  or (_34946_, _34945_, _34944_);
  and (_34947_, _34946_, _06152_);
  and (_34948_, _14928_, _07778_);
  or (_34949_, _34948_, _34939_);
  or (_34950_, _34949_, _06161_);
  and (_34951_, _07778_, \oc8051_golden_model_1.ACC [4]);
  or (_34952_, _34951_, _34939_);
  and (_34954_, _34952_, _07056_);
  and (_34955_, _07057_, \oc8051_golden_model_1.SCON [4]);
  or (_34956_, _34955_, _06160_);
  or (_34957_, _34956_, _34954_);
  and (_34958_, _34957_, _06157_);
  and (_34959_, _34958_, _34950_);
  and (_34960_, _14932_, _08413_);
  or (_34961_, _34960_, _34944_);
  and (_34962_, _34961_, _06156_);
  or (_34963_, _34962_, _06217_);
  or (_34965_, _34963_, _34959_);
  or (_34966_, _34941_, _07075_);
  and (_34967_, _34966_, _34965_);
  or (_34968_, _34967_, _06220_);
  or (_34969_, _34952_, _06229_);
  and (_34970_, _34969_, _06153_);
  and (_34971_, _34970_, _34968_);
  or (_34972_, _34971_, _34947_);
  and (_34973_, _34972_, _06146_);
  and (_34974_, _14950_, _08413_);
  or (_34976_, _34974_, _34944_);
  and (_34977_, _34976_, _06145_);
  or (_34978_, _34977_, _34973_);
  and (_34979_, _34978_, _06140_);
  and (_34980_, _14966_, _08413_);
  or (_34981_, _34980_, _34944_);
  and (_34982_, _34981_, _06139_);
  or (_34983_, _34982_, _09842_);
  or (_34984_, _34983_, _34979_);
  and (_34985_, _34984_, _34943_);
  or (_34987_, _34985_, _06116_);
  and (_34988_, _09209_, _07778_);
  or (_34989_, _34939_, _06117_);
  or (_34990_, _34989_, _34988_);
  and (_34991_, _34990_, _06114_);
  and (_34992_, _34991_, _34987_);
  and (_34993_, _15013_, _07778_);
  or (_34994_, _34993_, _34939_);
  and (_34995_, _34994_, _05787_);
  or (_34996_, _34995_, _11136_);
  or (_34998_, _34996_, _34992_);
  and (_34999_, _15029_, _07778_);
  or (_35000_, _34939_, _07127_);
  or (_35001_, _35000_, _34999_);
  and (_35002_, _08715_, _07778_);
  or (_35003_, _35002_, _34939_);
  or (_35004_, _35003_, _06111_);
  and (_35005_, _35004_, _07125_);
  and (_35006_, _35005_, _35001_);
  and (_35007_, _35006_, _34998_);
  and (_35009_, _10289_, _07778_);
  or (_35010_, _35009_, _34939_);
  and (_35011_, _35010_, _06402_);
  or (_35012_, _35011_, _35007_);
  and (_35013_, _35012_, _07132_);
  or (_35014_, _34939_, _08339_);
  and (_35015_, _35003_, _06306_);
  and (_35016_, _35015_, _35014_);
  or (_35017_, _35016_, _35013_);
  and (_35018_, _35017_, _07130_);
  and (_35020_, _34952_, _06411_);
  and (_35021_, _35020_, _35014_);
  or (_35022_, _35021_, _06303_);
  or (_35023_, _35022_, _35018_);
  and (_35024_, _15026_, _07778_);
  or (_35025_, _34939_, _08819_);
  or (_35026_, _35025_, _35024_);
  and (_35027_, _35026_, _08824_);
  and (_35028_, _35027_, _35023_);
  nor (_35029_, _10288_, _13504_);
  or (_35031_, _35029_, _34939_);
  and (_35032_, _35031_, _06396_);
  or (_35033_, _35032_, _06433_);
  or (_35034_, _35033_, _35028_);
  or (_35035_, _34949_, _06829_);
  and (_35036_, _35035_, _05749_);
  and (_35037_, _35036_, _35034_);
  and (_35038_, _34946_, _05748_);
  or (_35039_, _35038_, _06440_);
  or (_35040_, _35039_, _35037_);
  and (_35042_, _15087_, _07778_);
  or (_35043_, _34939_, _06444_);
  or (_35044_, _35043_, _35042_);
  and (_35045_, _35044_, _01317_);
  and (_35046_, _35045_, _35040_);
  or (_35047_, _35046_, _34938_);
  and (_43759_, _35047_, _43100_);
  and (_35048_, _01321_, \oc8051_golden_model_1.SCON [5]);
  and (_35049_, _13504_, \oc8051_golden_model_1.SCON [5]);
  and (_35050_, _15119_, _07778_);
  or (_35052_, _35050_, _35049_);
  or (_35053_, _35052_, _06161_);
  and (_35054_, _07778_, \oc8051_golden_model_1.ACC [5]);
  or (_35055_, _35054_, _35049_);
  and (_35056_, _35055_, _07056_);
  and (_35057_, _07057_, \oc8051_golden_model_1.SCON [5]);
  or (_35058_, _35057_, _06160_);
  or (_35059_, _35058_, _35056_);
  and (_35060_, _35059_, _06157_);
  and (_35061_, _35060_, _35053_);
  and (_35063_, _13509_, \oc8051_golden_model_1.SCON [5]);
  and (_35064_, _15123_, _08413_);
  or (_35065_, _35064_, _35063_);
  and (_35066_, _35065_, _06156_);
  or (_35067_, _35066_, _06217_);
  or (_35068_, _35067_, _35061_);
  and (_35069_, _08101_, _07778_);
  or (_35070_, _35069_, _35049_);
  or (_35071_, _35070_, _07075_);
  and (_35072_, _35071_, _35068_);
  or (_35074_, _35072_, _06220_);
  or (_35075_, _35055_, _06229_);
  and (_35076_, _35075_, _06153_);
  and (_35077_, _35076_, _35074_);
  and (_35078_, _15104_, _08413_);
  or (_35079_, _35078_, _35063_);
  and (_35080_, _35079_, _06152_);
  or (_35081_, _35080_, _06145_);
  or (_35082_, _35081_, _35077_);
  or (_35083_, _35063_, _15138_);
  and (_35085_, _35083_, _35065_);
  or (_35086_, _35085_, _06146_);
  and (_35087_, _35086_, _06140_);
  and (_35088_, _35087_, _35082_);
  and (_35089_, _15155_, _08413_);
  or (_35090_, _35089_, _35063_);
  and (_35091_, _35090_, _06139_);
  or (_35092_, _35091_, _09842_);
  or (_35093_, _35092_, _35088_);
  or (_35094_, _35070_, _06132_);
  and (_35096_, _35094_, _35093_);
  or (_35097_, _35096_, _06116_);
  and (_35098_, _09208_, _07778_);
  or (_35099_, _35049_, _06117_);
  or (_35100_, _35099_, _35098_);
  and (_35101_, _35100_, _06114_);
  and (_35102_, _35101_, _35097_);
  and (_35103_, _15203_, _07778_);
  or (_35104_, _35103_, _35049_);
  and (_35105_, _35104_, _05787_);
  or (_35107_, _35105_, _11136_);
  or (_35108_, _35107_, _35102_);
  and (_35109_, _15219_, _07778_);
  or (_35110_, _35049_, _07127_);
  or (_35111_, _35110_, _35109_);
  and (_35112_, _08736_, _07778_);
  or (_35113_, _35112_, _35049_);
  or (_35114_, _35113_, _06111_);
  and (_35115_, _35114_, _07125_);
  and (_35116_, _35115_, _35111_);
  and (_35118_, _35116_, _35108_);
  and (_35119_, _12325_, _07778_);
  or (_35120_, _35119_, _35049_);
  and (_35121_, _35120_, _06402_);
  or (_35122_, _35121_, _35118_);
  and (_35123_, _35122_, _07132_);
  or (_35124_, _35049_, _08104_);
  and (_35125_, _35113_, _06306_);
  and (_35126_, _35125_, _35124_);
  or (_35127_, _35126_, _35123_);
  and (_35129_, _35127_, _07130_);
  and (_35130_, _35055_, _06411_);
  and (_35131_, _35130_, _35124_);
  or (_35132_, _35131_, _06303_);
  or (_35133_, _35132_, _35129_);
  and (_35134_, _15216_, _07778_);
  or (_35135_, _35049_, _08819_);
  or (_35136_, _35135_, _35134_);
  and (_35137_, _35136_, _08824_);
  and (_35138_, _35137_, _35133_);
  nor (_35140_, _10269_, _13504_);
  or (_35141_, _35140_, _35049_);
  and (_35142_, _35141_, _06396_);
  or (_35143_, _35142_, _06433_);
  or (_35144_, _35143_, _35138_);
  or (_35145_, _35052_, _06829_);
  and (_35146_, _35145_, _05749_);
  and (_35147_, _35146_, _35144_);
  and (_35148_, _35079_, _05748_);
  or (_35149_, _35148_, _06440_);
  or (_35151_, _35149_, _35147_);
  and (_35152_, _15275_, _07778_);
  or (_35153_, _35049_, _06444_);
  or (_35154_, _35153_, _35152_);
  and (_35155_, _35154_, _01317_);
  and (_35156_, _35155_, _35151_);
  or (_35157_, _35156_, _35048_);
  and (_43761_, _35157_, _43100_);
  and (_35158_, _01321_, \oc8051_golden_model_1.SCON [6]);
  and (_35159_, _13504_, \oc8051_golden_model_1.SCON [6]);
  and (_35161_, _15300_, _07778_);
  or (_35162_, _35161_, _35159_);
  or (_35163_, _35162_, _06161_);
  and (_35164_, _07778_, \oc8051_golden_model_1.ACC [6]);
  or (_35165_, _35164_, _35159_);
  and (_35166_, _35165_, _07056_);
  and (_35167_, _07057_, \oc8051_golden_model_1.SCON [6]);
  or (_35168_, _35167_, _06160_);
  or (_35169_, _35168_, _35166_);
  and (_35170_, _35169_, _06157_);
  and (_35172_, _35170_, _35163_);
  and (_35173_, _13509_, \oc8051_golden_model_1.SCON [6]);
  and (_35174_, _15316_, _08413_);
  or (_35175_, _35174_, _35173_);
  and (_35176_, _35175_, _06156_);
  or (_35177_, _35176_, _06217_);
  or (_35178_, _35177_, _35172_);
  and (_35179_, _08012_, _07778_);
  or (_35180_, _35179_, _35159_);
  or (_35181_, _35180_, _07075_);
  and (_35183_, _35181_, _35178_);
  or (_35184_, _35183_, _06220_);
  or (_35185_, _35165_, _06229_);
  and (_35186_, _35185_, _06153_);
  and (_35187_, _35186_, _35184_);
  and (_35188_, _15297_, _08413_);
  or (_35189_, _35188_, _35173_);
  and (_35190_, _35189_, _06152_);
  or (_35191_, _35190_, _06145_);
  or (_35192_, _35191_, _35187_);
  or (_35194_, _35173_, _15331_);
  and (_35195_, _35194_, _35175_);
  or (_35196_, _35195_, _06146_);
  and (_35197_, _35196_, _06140_);
  and (_35198_, _35197_, _35192_);
  and (_35199_, _15348_, _08413_);
  or (_35200_, _35199_, _35173_);
  and (_35201_, _35200_, _06139_);
  or (_35202_, _35201_, _09842_);
  or (_35203_, _35202_, _35198_);
  or (_35205_, _35180_, _06132_);
  and (_35206_, _35205_, _35203_);
  or (_35207_, _35206_, _06116_);
  and (_35208_, _09207_, _07778_);
  or (_35209_, _35159_, _06117_);
  or (_35210_, _35209_, _35208_);
  and (_35211_, _35210_, _06114_);
  and (_35212_, _35211_, _35207_);
  and (_35213_, _15395_, _07778_);
  or (_35214_, _35213_, _35159_);
  and (_35216_, _35214_, _05787_);
  or (_35217_, _35216_, _11136_);
  or (_35218_, _35217_, _35212_);
  and (_35219_, _15413_, _07778_);
  or (_35220_, _35159_, _07127_);
  or (_35221_, _35220_, _35219_);
  and (_35222_, _15402_, _07778_);
  or (_35223_, _35222_, _35159_);
  or (_35224_, _35223_, _06111_);
  and (_35225_, _35224_, _07125_);
  and (_35227_, _35225_, _35221_);
  and (_35228_, _35227_, _35218_);
  and (_35229_, _10295_, _07778_);
  or (_35230_, _35229_, _35159_);
  and (_35231_, _35230_, _06402_);
  or (_35232_, _35231_, _35228_);
  and (_35233_, _35232_, _07132_);
  or (_35234_, _35159_, _08015_);
  and (_35235_, _35223_, _06306_);
  and (_35236_, _35235_, _35234_);
  or (_35238_, _35236_, _35233_);
  and (_35239_, _35238_, _07130_);
  and (_35240_, _35165_, _06411_);
  and (_35241_, _35240_, _35234_);
  or (_35242_, _35241_, _06303_);
  or (_35243_, _35242_, _35239_);
  and (_35244_, _15410_, _07778_);
  or (_35245_, _35159_, _08819_);
  or (_35246_, _35245_, _35244_);
  and (_35247_, _35246_, _08824_);
  and (_35249_, _35247_, _35243_);
  nor (_35250_, _10294_, _13504_);
  or (_35251_, _35250_, _35159_);
  and (_35252_, _35251_, _06396_);
  or (_35253_, _35252_, _06433_);
  or (_35254_, _35253_, _35249_);
  or (_35255_, _35162_, _06829_);
  and (_35256_, _35255_, _05749_);
  and (_35257_, _35256_, _35254_);
  and (_35258_, _35189_, _05748_);
  or (_35260_, _35258_, _06440_);
  or (_35261_, _35260_, _35257_);
  and (_35262_, _15478_, _07778_);
  or (_35263_, _35159_, _06444_);
  or (_35264_, _35263_, _35262_);
  and (_35265_, _35264_, _01317_);
  and (_35266_, _35265_, _35261_);
  or (_35267_, _35266_, _35158_);
  and (_43762_, _35267_, _43100_);
  nor (_35268_, _01317_, _06142_);
  nor (_35270_, _13615_, _06142_);
  and (_35271_, _13615_, \oc8051_golden_model_1.ACC [0]);
  and (_35272_, _35271_, _08211_);
  or (_35273_, _35272_, _35270_);
  or (_35274_, _35273_, _07130_);
  nor (_35275_, _08211_, _13718_);
  or (_35276_, _35275_, _35270_);
  or (_35277_, _35276_, _06161_);
  or (_35278_, _35271_, _35270_);
  and (_35279_, _35278_, _07056_);
  nor (_35281_, _07056_, _06142_);
  or (_35282_, _35281_, _06160_);
  or (_35283_, _35282_, _35279_);
  and (_35284_, _35283_, _07075_);
  and (_35285_, _35284_, _35277_);
  or (_35286_, _35285_, _06671_);
  or (_35287_, _35278_, _06229_);
  and (_35288_, _35287_, _07191_);
  and (_35289_, _35288_, _35286_);
  nand (_35290_, _06132_, _07093_);
  or (_35292_, _35290_, _35289_);
  and (_35293_, _07858_, _07049_);
  or (_35294_, _35270_, _06132_);
  or (_35295_, _35294_, _35293_);
  and (_35296_, _35295_, _35292_);
  or (_35297_, _35296_, _06116_);
  or (_35298_, _35270_, _06117_);
  and (_35299_, _09160_, _13615_);
  or (_35300_, _35299_, _35298_);
  and (_35301_, _35300_, _35297_);
  or (_35303_, _35301_, _05787_);
  and (_35304_, _14260_, _07858_);
  or (_35305_, _35270_, _06114_);
  or (_35306_, _35305_, _35304_);
  and (_35307_, _35306_, _06111_);
  and (_35308_, _35307_, _35303_);
  and (_35309_, _13615_, _08708_);
  or (_35310_, _35309_, _35270_);
  and (_35311_, _35310_, _06110_);
  or (_35312_, _35311_, _06297_);
  or (_35314_, _35312_, _35308_);
  and (_35315_, _14275_, _13615_);
  or (_35316_, _35315_, _35270_);
  or (_35317_, _35316_, _07127_);
  and (_35318_, _35317_, _07125_);
  and (_35319_, _35318_, _35314_);
  nor (_35320_, _12321_, _13718_);
  or (_35321_, _35320_, _35270_);
  nor (_35322_, _35272_, _07125_);
  and (_35323_, _35322_, _35321_);
  or (_35325_, _35323_, _35319_);
  and (_35326_, _35325_, _07132_);
  nand (_35327_, _35310_, _06306_);
  nor (_35328_, _35327_, _35275_);
  or (_35329_, _35328_, _06411_);
  or (_35330_, _35329_, _35326_);
  and (_35331_, _35330_, _35274_);
  or (_35332_, _35331_, _06303_);
  and (_35333_, _14167_, _07858_);
  or (_35334_, _35270_, _08819_);
  or (_35336_, _35334_, _35333_);
  and (_35337_, _35336_, _08824_);
  and (_35338_, _35337_, _35332_);
  and (_35339_, _35321_, _06396_);
  or (_35340_, _35339_, _19287_);
  or (_35341_, _35340_, _35338_);
  or (_35342_, _35276_, _06630_);
  and (_35343_, _35342_, _01317_);
  and (_35344_, _35343_, _35341_);
  or (_35345_, _35344_, _35268_);
  and (_43763_, _35345_, _43100_);
  nand (_35347_, _06417_, \oc8051_golden_model_1.SP [1]);
  nand (_35348_, _07858_, _06945_);
  or (_35349_, _35348_, _08176_);
  or (_35350_, _13615_, \oc8051_golden_model_1.SP [1]);
  and (_35351_, _35350_, _06303_);
  and (_35352_, _35351_, _35349_);
  and (_35353_, _35350_, _05787_);
  or (_35354_, _14442_, _13718_);
  and (_35355_, _35354_, _35353_);
  and (_35357_, _14363_, _07858_);
  not (_35358_, _35357_);
  and (_35359_, _35358_, _35350_);
  or (_35360_, _35359_, _06161_);
  nor (_35361_, _13615_, _06979_);
  and (_35362_, _13615_, \oc8051_golden_model_1.ACC [1]);
  or (_35363_, _35362_, _35361_);
  or (_35364_, _35363_, _07057_);
  or (_35365_, _07056_, \oc8051_golden_model_1.SP [1]);
  and (_35366_, _35365_, _06582_);
  and (_35368_, _35366_, _35364_);
  and (_35369_, _06581_, _06979_);
  or (_35370_, _35369_, _06160_);
  or (_35371_, _35370_, _35368_);
  and (_35372_, _35371_, _05764_);
  and (_35373_, _35372_, _35360_);
  nor (_35374_, _05764_, \oc8051_golden_model_1.SP [1]);
  or (_35375_, _35374_, _06217_);
  or (_35376_, _35375_, _35373_);
  nand (_35377_, _07189_, _06217_);
  and (_35379_, _35377_, _35376_);
  or (_35380_, _35379_, _06220_);
  or (_35381_, _35363_, _06229_);
  and (_35382_, _35381_, _07191_);
  and (_35383_, _35382_, _35380_);
  not (_35384_, _07389_);
  or (_35385_, _35384_, _07190_);
  or (_35386_, _35385_, _35383_);
  or (_35387_, _07389_, _06979_);
  and (_35388_, _35387_, _06132_);
  and (_35390_, _35388_, _35386_);
  or (_35391_, _13718_, _07306_);
  and (_35392_, _35350_, _09842_);
  and (_35393_, _35392_, _35391_);
  or (_35394_, _35393_, _06116_);
  or (_35395_, _35394_, _35390_);
  or (_35396_, _35361_, _06117_);
  and (_35397_, _09115_, _13615_);
  or (_35398_, _35397_, _35396_);
  and (_35399_, _35398_, _06114_);
  and (_35401_, _35399_, _35395_);
  or (_35402_, _35401_, _35355_);
  and (_35403_, _35402_, _06111_);
  and (_35404_, _35350_, _06110_);
  and (_35405_, _35404_, _35348_);
  or (_35406_, _35405_, _06076_);
  or (_35407_, _35406_, _35403_);
  or (_35408_, _05836_, _06979_);
  and (_35409_, _35408_, _07127_);
  and (_35410_, _35409_, _35407_);
  or (_35412_, _14346_, _13718_);
  and (_35413_, _35350_, _06297_);
  and (_35414_, _35413_, _35412_);
  or (_35415_, _35414_, _06402_);
  or (_35416_, _35415_, _35410_);
  and (_35417_, _10278_, _13615_);
  or (_35418_, _35417_, _35361_);
  or (_35419_, _35418_, _07125_);
  and (_35420_, _35419_, _07132_);
  and (_35421_, _35420_, _35416_);
  or (_35423_, _14344_, _13718_);
  and (_35424_, _35350_, _06306_);
  and (_35425_, _35424_, _35423_);
  or (_35426_, _35425_, _06411_);
  or (_35427_, _35426_, _35421_);
  and (_35428_, _35362_, _08176_);
  or (_35429_, _35428_, _35361_);
  or (_35430_, _35429_, _07130_);
  and (_35431_, _35430_, _35427_);
  or (_35432_, _35431_, _07124_);
  nor (_35434_, _05848_, _06979_);
  nor (_35435_, _35434_, _06303_);
  and (_35436_, _35435_, _35432_);
  or (_35437_, _35436_, _35352_);
  and (_35438_, _35437_, _08824_);
  nor (_35439_, _10277_, _13718_);
  or (_35440_, _35439_, _35361_);
  and (_35441_, _35440_, _06396_);
  or (_35442_, _35441_, _06417_);
  or (_35443_, _35442_, _35438_);
  nand (_35445_, _35443_, _35347_);
  nor (_35446_, _06167_, _07142_);
  nand (_35447_, _35446_, _35445_);
  or (_35448_, _35446_, _06979_);
  and (_35449_, _35448_, _06829_);
  and (_35450_, _35449_, _35447_);
  and (_35451_, _35359_, _06433_);
  or (_35452_, _35451_, _07577_);
  or (_35453_, _35452_, _35450_);
  or (_35454_, _07160_, _06979_);
  and (_35456_, _35454_, _06444_);
  and (_35457_, _35456_, _35453_);
  or (_35458_, _35357_, _35361_);
  and (_35459_, _35458_, _06440_);
  or (_35460_, _35459_, _01321_);
  or (_35461_, _35460_, _35457_);
  or (_35462_, _01317_, \oc8051_golden_model_1.SP [1]);
  and (_35463_, _35462_, _43100_);
  and (_43765_, _35463_, _35461_);
  nor (_35464_, _01317_, _06566_);
  or (_35466_, _07755_, _05836_);
  and (_35467_, _07858_, _07708_);
  nor (_35468_, _13615_, _06566_);
  or (_35469_, _35468_, _06132_);
  or (_35470_, _35469_, _35467_);
  and (_35471_, _14542_, _07858_);
  or (_35472_, _35471_, _35468_);
  or (_35473_, _35472_, _06161_);
  and (_35474_, _13615_, \oc8051_golden_model_1.ACC [2]);
  or (_35475_, _35474_, _35468_);
  or (_35477_, _35475_, _07057_);
  or (_35478_, _07056_, \oc8051_golden_model_1.SP [2]);
  and (_35479_, _35478_, _06582_);
  and (_35480_, _35479_, _35477_);
  and (_35481_, _07755_, _06581_);
  or (_35482_, _35481_, _06160_);
  or (_35483_, _35482_, _35480_);
  and (_35484_, _35483_, _05764_);
  and (_35485_, _35484_, _35473_);
  nor (_35486_, _15819_, _05764_);
  or (_35488_, _35486_, _06217_);
  or (_35489_, _35488_, _35485_);
  nand (_35490_, _08465_, _06217_);
  and (_35491_, _35490_, _35489_);
  or (_35492_, _35491_, _06220_);
  or (_35493_, _35475_, _06229_);
  and (_35494_, _35493_, _07191_);
  and (_35495_, _35494_, _35492_);
  or (_35496_, _07601_, _07388_);
  or (_35497_, _35496_, _35495_);
  nor (_35499_, _07755_, _05760_);
  nor (_35500_, _35499_, _05791_);
  and (_35501_, _35500_, _35497_);
  nand (_35502_, _07755_, _05791_);
  nand (_35503_, _35502_, _06132_);
  or (_35504_, _35503_, _35501_);
  and (_35505_, _35504_, _35470_);
  or (_35506_, _35505_, _06116_);
  or (_35507_, _35468_, _06117_);
  and (_35508_, _09211_, _13615_);
  or (_35510_, _35508_, _35507_);
  and (_35511_, _35510_, _06114_);
  and (_35512_, _35511_, _35506_);
  and (_35513_, _14630_, _13615_);
  or (_35514_, _35513_, _35468_);
  and (_35515_, _35514_, _05787_);
  or (_35516_, _35515_, _06110_);
  or (_35517_, _35516_, _35512_);
  and (_35518_, _13615_, _08768_);
  or (_35519_, _35518_, _35468_);
  or (_35521_, _35519_, _06111_);
  and (_35522_, _35521_, _35517_);
  or (_35523_, _35522_, _06076_);
  and (_35524_, _35523_, _35466_);
  or (_35525_, _35524_, _06297_);
  and (_35526_, _14646_, _13615_);
  or (_35527_, _35526_, _35468_);
  or (_35528_, _35527_, _07127_);
  and (_35529_, _35528_, _07125_);
  and (_35530_, _35529_, _35525_);
  and (_35532_, _10282_, _13615_);
  or (_35533_, _35532_, _35468_);
  and (_35534_, _35533_, _06402_);
  or (_35535_, _35534_, _35530_);
  and (_35536_, _35535_, _07132_);
  or (_35537_, _35468_, _08248_);
  and (_35538_, _35519_, _06306_);
  and (_35539_, _35538_, _35537_);
  or (_35540_, _35539_, _35536_);
  and (_35541_, _35540_, _12514_);
  and (_35543_, _35475_, _06411_);
  and (_35544_, _35543_, _35537_);
  nor (_35545_, _15819_, _05848_);
  or (_35546_, _35545_, _06303_);
  or (_35547_, _35546_, _35544_);
  or (_35548_, _35547_, _35541_);
  and (_35549_, _14643_, _07858_);
  or (_35550_, _35468_, _08819_);
  or (_35551_, _35550_, _35549_);
  and (_35552_, _35551_, _35548_);
  or (_35554_, _35552_, _06396_);
  nor (_35555_, _10281_, _13718_);
  or (_35556_, _35555_, _35468_);
  or (_35557_, _35556_, _08824_);
  and (_35558_, _35557_, _12558_);
  and (_35559_, _35558_, _35554_);
  and (_35560_, _15819_, _06417_);
  or (_35561_, _35560_, _07142_);
  or (_35562_, _35561_, _35559_);
  or (_35563_, _07755_, _05846_);
  and (_35565_, _35563_, _06168_);
  and (_35566_, _35565_, _35562_);
  and (_35567_, _15819_, _06167_);
  or (_35568_, _35567_, _06433_);
  or (_35569_, _35568_, _35566_);
  or (_35570_, _35472_, _06829_);
  and (_35571_, _35570_, _07160_);
  and (_35572_, _35571_, _35569_);
  nor (_35573_, _15819_, _07160_);
  or (_35574_, _35573_, _06440_);
  or (_35576_, _35574_, _35572_);
  and (_35577_, _14710_, _07858_);
  or (_35578_, _35468_, _06444_);
  or (_35579_, _35578_, _35577_);
  and (_35580_, _35579_, _01317_);
  and (_35581_, _35580_, _35576_);
  or (_35582_, _35581_, _35464_);
  and (_43766_, _35582_, _43100_);
  nor (_35583_, _01317_, _06216_);
  or (_35584_, _07759_, _07160_);
  or (_35586_, _07759_, _05836_);
  and (_35587_, _07858_, _07544_);
  nor (_35588_, _13615_, _06216_);
  or (_35589_, _35588_, _06116_);
  or (_35590_, _35589_, _35587_);
  and (_35591_, _35590_, _13620_);
  and (_35592_, _14738_, _07858_);
  or (_35593_, _35592_, _35588_);
  or (_35594_, _35593_, _06161_);
  and (_35595_, _13615_, \oc8051_golden_model_1.ACC [3]);
  or (_35597_, _35595_, _35588_);
  or (_35598_, _35597_, _07057_);
  or (_35599_, _07056_, \oc8051_golden_model_1.SP [3]);
  and (_35600_, _35599_, _06582_);
  and (_35601_, _35600_, _35598_);
  and (_35602_, _07759_, _06581_);
  or (_35603_, _35602_, _06160_);
  or (_35604_, _35603_, _35601_);
  and (_35605_, _35604_, _05764_);
  and (_35606_, _35605_, _35594_);
  nor (_35608_, _15639_, _05764_);
  or (_35609_, _35608_, _06217_);
  or (_35610_, _35609_, _35606_);
  nand (_35611_, _08455_, _06217_);
  and (_35612_, _35611_, _35610_);
  or (_35613_, _35612_, _06220_);
  or (_35614_, _35597_, _06229_);
  and (_35615_, _35614_, _07191_);
  and (_35616_, _35615_, _35613_);
  or (_35617_, _07525_, _35384_);
  or (_35619_, _35617_, _35616_);
  or (_35620_, _07759_, _07389_);
  and (_35621_, _35620_, _06132_);
  and (_35622_, _35621_, _35619_);
  or (_35623_, _35622_, _35591_);
  or (_35624_, _35588_, _06117_);
  and (_35625_, _09210_, _13615_);
  or (_35626_, _35625_, _35624_);
  and (_35627_, _35626_, _06114_);
  and (_35628_, _35627_, _35623_);
  and (_35630_, _14825_, _13615_);
  or (_35631_, _35630_, _35588_);
  and (_35632_, _35631_, _05787_);
  or (_35633_, _35632_, _06110_);
  or (_35634_, _35633_, _35628_);
  and (_35635_, _13615_, _08712_);
  or (_35636_, _35635_, _35588_);
  or (_35637_, _35636_, _06111_);
  and (_35638_, _35637_, _35634_);
  or (_35639_, _35638_, _06076_);
  and (_35641_, _35639_, _35586_);
  or (_35642_, _35641_, _06297_);
  and (_35643_, _14727_, _13615_);
  or (_35644_, _35643_, _35588_);
  or (_35645_, _35644_, _07127_);
  and (_35646_, _35645_, _07125_);
  and (_35647_, _35646_, _35642_);
  and (_35648_, _12318_, _13615_);
  or (_35649_, _35648_, _35588_);
  and (_35650_, _35649_, _06402_);
  or (_35652_, _35650_, _35647_);
  and (_35653_, _35652_, _07132_);
  or (_35654_, _35588_, _08140_);
  and (_35655_, _35636_, _06306_);
  and (_35656_, _35655_, _35654_);
  or (_35657_, _35656_, _35653_);
  and (_35658_, _35657_, _12514_);
  and (_35659_, _35597_, _06411_);
  and (_35660_, _35659_, _35654_);
  nor (_35661_, _15639_, _05848_);
  or (_35663_, _35661_, _06303_);
  or (_35664_, _35663_, _35660_);
  or (_35665_, _35664_, _35658_);
  and (_35666_, _14724_, _07858_);
  or (_35667_, _35588_, _08819_);
  or (_35668_, _35667_, _35666_);
  and (_35669_, _35668_, _35665_);
  or (_35670_, _35669_, _06396_);
  nor (_35671_, _10273_, _13718_);
  or (_35672_, _35671_, _35588_);
  or (_35674_, _35672_, _08824_);
  and (_35675_, _35674_, _12558_);
  and (_35676_, _35675_, _35670_);
  nor (_35677_, _08452_, _06216_);
  or (_35678_, _35677_, _08453_);
  and (_35679_, _35678_, _06417_);
  or (_35680_, _35679_, _07142_);
  or (_35681_, _35680_, _35676_);
  or (_35682_, _07759_, _05846_);
  and (_35683_, _35682_, _35681_);
  or (_35685_, _35683_, _06167_);
  or (_35686_, _35678_, _06168_);
  and (_35687_, _35686_, _06829_);
  and (_35688_, _35687_, _35685_);
  and (_35689_, _35593_, _06433_);
  or (_35690_, _35689_, _07577_);
  or (_35691_, _35690_, _35688_);
  and (_35692_, _35691_, _35584_);
  or (_35693_, _35692_, _06440_);
  and (_35694_, _14897_, _07858_);
  or (_35695_, _35588_, _06444_);
  or (_35696_, _35695_, _35694_);
  and (_35697_, _35696_, _01317_);
  and (_35698_, _35697_, _35693_);
  or (_35699_, _35698_, _35583_);
  and (_43767_, _35699_, _43100_);
  nor (_35700_, _01317_, _13644_);
  nor (_35701_, _07756_, \oc8051_golden_model_1.SP [4]);
  nor (_35702_, _35701_, _13607_);
  or (_35703_, _35702_, _07160_);
  or (_35705_, _35702_, _05846_);
  and (_35706_, _08336_, _07858_);
  nor (_35707_, _13615_, _13644_);
  or (_35708_, _35707_, _06116_);
  or (_35709_, _35708_, _35706_);
  and (_35710_, _35709_, _13620_);
  and (_35711_, _14928_, _07858_);
  or (_35712_, _35711_, _35707_);
  or (_35713_, _35712_, _06161_);
  and (_35714_, _13615_, \oc8051_golden_model_1.ACC [4]);
  or (_35716_, _35714_, _35707_);
  or (_35717_, _35716_, _07057_);
  or (_35718_, _07056_, \oc8051_golden_model_1.SP [4]);
  and (_35719_, _35718_, _06582_);
  and (_35720_, _35719_, _35717_);
  and (_35721_, _35702_, _06581_);
  or (_35722_, _35721_, _06160_);
  or (_35723_, _35722_, _35720_);
  and (_35724_, _35723_, _05764_);
  and (_35725_, _35724_, _35713_);
  and (_35727_, _35702_, _07485_);
  or (_35728_, _35727_, _06217_);
  or (_35729_, _35728_, _35725_);
  and (_35730_, _13645_, _06142_);
  nor (_35731_, _08454_, _13644_);
  nor (_35732_, _35731_, _35730_);
  nand (_35733_, _35732_, _06217_);
  and (_35734_, _35733_, _35729_);
  or (_35735_, _35734_, _06220_);
  or (_35736_, _35716_, _06229_);
  and (_35738_, _35736_, _07191_);
  and (_35739_, _35738_, _35735_);
  and (_35740_, _07479_, \oc8051_golden_model_1.SP [4]);
  nor (_35741_, _07479_, \oc8051_golden_model_1.SP [4]);
  nor (_35742_, _35741_, _35740_);
  nand (_35743_, _35742_, _06151_);
  nand (_35744_, _35743_, _07389_);
  or (_35745_, _35744_, _35739_);
  or (_35746_, _35702_, _07389_);
  and (_35747_, _35746_, _06132_);
  and (_35749_, _35747_, _35745_);
  or (_35750_, _35749_, _35710_);
  or (_35751_, _35707_, _06117_);
  and (_35752_, _09209_, _13615_);
  or (_35753_, _35752_, _35751_);
  and (_35754_, _35753_, _06114_);
  and (_35755_, _35754_, _35750_);
  and (_35756_, _15013_, _13615_);
  or (_35757_, _35756_, _35707_);
  and (_35758_, _35757_, _05787_);
  or (_35760_, _35758_, _06110_);
  or (_35761_, _35760_, _35755_);
  and (_35762_, _08715_, _13615_);
  or (_35763_, _35762_, _35707_);
  or (_35764_, _35763_, _06111_);
  and (_35765_, _35764_, _35761_);
  or (_35766_, _35765_, _06076_);
  or (_35767_, _35702_, _05836_);
  and (_35768_, _35767_, _35766_);
  or (_35769_, _35768_, _06297_);
  and (_35771_, _15029_, _07858_);
  or (_35772_, _35707_, _07127_);
  or (_35773_, _35772_, _35771_);
  and (_35774_, _35773_, _07125_);
  and (_35775_, _35774_, _35769_);
  and (_35776_, _10289_, _13615_);
  or (_35777_, _35776_, _35707_);
  and (_35778_, _35777_, _06402_);
  or (_35779_, _35778_, _35775_);
  and (_35780_, _35779_, _07132_);
  or (_35782_, _35707_, _08339_);
  and (_35783_, _35763_, _06306_);
  and (_35784_, _35783_, _35782_);
  or (_35785_, _35784_, _35780_);
  and (_35786_, _35785_, _12514_);
  and (_35787_, _35716_, _06411_);
  and (_35788_, _35787_, _35782_);
  and (_35789_, _35702_, _07124_);
  or (_35790_, _35789_, _06303_);
  or (_35791_, _35790_, _35788_);
  or (_35793_, _35791_, _35786_);
  and (_35794_, _15026_, _07858_);
  or (_35795_, _35707_, _08819_);
  or (_35796_, _35795_, _35794_);
  and (_35797_, _35796_, _35793_);
  or (_35798_, _35797_, _06396_);
  nor (_35799_, _10288_, _13718_);
  or (_35800_, _35799_, _35707_);
  or (_35801_, _35800_, _08824_);
  and (_35802_, _35801_, _12558_);
  and (_35804_, _35802_, _35798_);
  nor (_35805_, _08453_, _13644_);
  or (_35806_, _35805_, _13645_);
  and (_35807_, _35806_, _06417_);
  or (_35808_, _35807_, _07142_);
  or (_35809_, _35808_, _35804_);
  and (_35810_, _35809_, _35705_);
  or (_35811_, _35810_, _06167_);
  or (_35812_, _35806_, _06168_);
  and (_35813_, _35812_, _06829_);
  and (_35815_, _35813_, _35811_);
  and (_35816_, _35712_, _06433_);
  or (_35817_, _35816_, _07577_);
  or (_35818_, _35817_, _35815_);
  and (_35819_, _35818_, _35703_);
  or (_35820_, _35819_, _06440_);
  and (_35821_, _15087_, _07858_);
  or (_35822_, _35707_, _06444_);
  or (_35823_, _35822_, _35821_);
  and (_35824_, _35823_, _01317_);
  and (_35826_, _35824_, _35820_);
  or (_35827_, _35826_, _35700_);
  and (_43768_, _35827_, _43100_);
  nor (_35828_, _01317_, _13643_);
  nor (_35829_, _13607_, \oc8051_golden_model_1.SP [5]);
  nor (_35830_, _35829_, _13608_);
  or (_35831_, _35830_, _07160_);
  and (_35832_, _08101_, _07858_);
  nor (_35833_, _13615_, _13643_);
  or (_35834_, _35833_, _06116_);
  or (_35836_, _35834_, _35832_);
  and (_35837_, _35836_, _13620_);
  and (_35838_, _15119_, _07858_);
  or (_35839_, _35838_, _35833_);
  or (_35840_, _35839_, _06161_);
  and (_35841_, _13615_, \oc8051_golden_model_1.ACC [5]);
  or (_35842_, _35841_, _35833_);
  or (_35843_, _35842_, _07057_);
  or (_35844_, _07056_, \oc8051_golden_model_1.SP [5]);
  and (_35845_, _35844_, _06582_);
  and (_35847_, _35845_, _35843_);
  and (_35848_, _35830_, _06581_);
  or (_35849_, _35848_, _06160_);
  or (_35850_, _35849_, _35847_);
  and (_35851_, _35850_, _05764_);
  and (_35852_, _35851_, _35840_);
  and (_35853_, _35830_, _07485_);
  or (_35854_, _35853_, _06217_);
  or (_35855_, _35854_, _35852_);
  and (_35856_, _13646_, _06142_);
  nor (_35858_, _35730_, _13643_);
  nor (_35859_, _35858_, _35856_);
  nand (_35860_, _35859_, _06217_);
  and (_35861_, _35860_, _35855_);
  or (_35862_, _35861_, _06220_);
  or (_35863_, _35842_, _06229_);
  and (_35864_, _35863_, _07191_);
  and (_35865_, _35864_, _35862_);
  nor (_35866_, _35740_, \oc8051_golden_model_1.SP [5]);
  nor (_35867_, _35866_, _13659_);
  nand (_35869_, _35867_, _06151_);
  nand (_35870_, _35869_, _07389_);
  or (_35871_, _35870_, _35865_);
  or (_35872_, _35830_, _07389_);
  and (_35873_, _35872_, _06132_);
  and (_35874_, _35873_, _35871_);
  or (_35875_, _35874_, _35837_);
  or (_35876_, _35833_, _06117_);
  and (_35877_, _09208_, _13615_);
  or (_35878_, _35877_, _35876_);
  and (_35880_, _35878_, _06114_);
  and (_35881_, _35880_, _35875_);
  and (_35882_, _15203_, _13615_);
  or (_35883_, _35882_, _35833_);
  and (_35884_, _35883_, _05787_);
  or (_35885_, _35884_, _06110_);
  or (_35886_, _35885_, _35881_);
  and (_35887_, _08736_, _13615_);
  or (_35888_, _35887_, _35833_);
  or (_35889_, _35888_, _06111_);
  and (_35891_, _35889_, _35886_);
  or (_35892_, _35891_, _06076_);
  or (_35893_, _35830_, _05836_);
  and (_35894_, _35893_, _35892_);
  or (_35895_, _35894_, _06297_);
  and (_35896_, _15219_, _07858_);
  or (_35897_, _35833_, _07127_);
  or (_35898_, _35897_, _35896_);
  and (_35899_, _35898_, _07125_);
  and (_35900_, _35899_, _35895_);
  and (_35902_, _12325_, _13615_);
  or (_35903_, _35902_, _35833_);
  and (_35904_, _35903_, _06402_);
  or (_35905_, _35904_, _35900_);
  and (_35906_, _35905_, _07132_);
  or (_35907_, _35833_, _08104_);
  and (_35908_, _35888_, _06306_);
  and (_35909_, _35908_, _35907_);
  or (_35910_, _35909_, _35906_);
  and (_35911_, _35910_, _12514_);
  and (_35913_, _35842_, _06411_);
  and (_35914_, _35913_, _35907_);
  and (_35915_, _35830_, _07124_);
  or (_35916_, _35915_, _06303_);
  or (_35917_, _35916_, _35914_);
  or (_35918_, _35917_, _35911_);
  and (_35919_, _15216_, _07858_);
  or (_35920_, _35833_, _08819_);
  or (_35921_, _35920_, _35919_);
  and (_35922_, _35921_, _35918_);
  or (_35924_, _35922_, _06396_);
  nor (_35925_, _10269_, _13718_);
  or (_35926_, _35925_, _35833_);
  or (_35927_, _35926_, _08824_);
  and (_35928_, _35927_, _12558_);
  and (_35929_, _35928_, _35924_);
  nor (_35930_, _13645_, _13643_);
  or (_35931_, _35930_, _13646_);
  and (_35932_, _35931_, _06417_);
  or (_35933_, _35932_, _07142_);
  or (_35935_, _35933_, _35929_);
  or (_35936_, _35830_, _05846_);
  and (_35937_, _35936_, _35935_);
  or (_35938_, _35937_, _06167_);
  or (_35939_, _35931_, _06168_);
  and (_35940_, _35939_, _06829_);
  and (_35941_, _35940_, _35938_);
  and (_35942_, _35839_, _06433_);
  or (_35943_, _35942_, _07577_);
  or (_35944_, _35943_, _35941_);
  and (_35946_, _35944_, _35831_);
  or (_35947_, _35946_, _06440_);
  and (_35948_, _15275_, _07858_);
  or (_35949_, _35833_, _06444_);
  or (_35950_, _35949_, _35948_);
  and (_35951_, _35950_, _01317_);
  and (_35952_, _35951_, _35947_);
  or (_35953_, _35952_, _35828_);
  and (_43769_, _35953_, _43100_);
  nor (_35954_, _01317_, _13642_);
  nor (_35956_, _13615_, _13642_);
  and (_35957_, _15300_, _07858_);
  or (_35958_, _35957_, _35956_);
  or (_35959_, _35958_, _06161_);
  and (_35960_, _13615_, \oc8051_golden_model_1.ACC [6]);
  or (_35961_, _35960_, _35956_);
  or (_35962_, _35961_, _07057_);
  or (_35963_, _07056_, \oc8051_golden_model_1.SP [6]);
  and (_35964_, _35963_, _06582_);
  and (_35965_, _35964_, _35962_);
  nor (_35967_, _13608_, \oc8051_golden_model_1.SP [6]);
  nor (_35968_, _35967_, _13609_);
  and (_35969_, _35968_, _06581_);
  or (_35970_, _35969_, _06160_);
  or (_35971_, _35970_, _35965_);
  and (_35972_, _35971_, _05764_);
  and (_35973_, _35972_, _35959_);
  and (_35974_, _35968_, _07485_);
  or (_35975_, _35974_, _06217_);
  or (_35976_, _35975_, _35973_);
  nor (_35978_, _35856_, _13642_);
  nor (_35979_, _35978_, _13648_);
  nand (_35980_, _35979_, _06217_);
  and (_35981_, _35980_, _35976_);
  or (_35982_, _35981_, _06220_);
  or (_35983_, _35961_, _06229_);
  and (_35984_, _35983_, _07191_);
  and (_35985_, _35984_, _35982_);
  nor (_35986_, _13659_, \oc8051_golden_model_1.SP [6]);
  nor (_35987_, _35986_, _13661_);
  and (_35989_, _35987_, _06151_);
  or (_35990_, _35989_, _35985_);
  and (_35991_, _35990_, _07389_);
  nand (_35992_, _35968_, _35384_);
  nand (_35993_, _35992_, _06132_);
  or (_35994_, _35993_, _35991_);
  and (_35995_, _08012_, _07858_);
  or (_35996_, _35956_, _06132_);
  or (_35997_, _35996_, _35995_);
  and (_35998_, _35997_, _35994_);
  or (_36000_, _35998_, _06116_);
  and (_36001_, _09207_, _13615_);
  or (_36002_, _35956_, _06117_);
  or (_36003_, _36002_, _36001_);
  and (_36004_, _36003_, _06114_);
  and (_36005_, _36004_, _36000_);
  and (_36006_, _15395_, _07858_);
  or (_36007_, _36006_, _35956_);
  and (_36008_, _36007_, _05787_);
  or (_36009_, _36008_, _06110_);
  or (_36011_, _36009_, _36005_);
  and (_36012_, _15402_, _13615_);
  or (_36013_, _36012_, _35956_);
  or (_36014_, _36013_, _06111_);
  and (_36015_, _36014_, _36011_);
  or (_36016_, _36015_, _06076_);
  or (_36017_, _35968_, _05836_);
  and (_36018_, _36017_, _36016_);
  or (_36019_, _36018_, _06297_);
  and (_36020_, _15413_, _07858_);
  or (_36022_, _35956_, _07127_);
  or (_36023_, _36022_, _36020_);
  and (_36024_, _36023_, _07125_);
  and (_36025_, _36024_, _36019_);
  and (_36026_, _10295_, _13615_);
  or (_36027_, _36026_, _35956_);
  and (_36028_, _36027_, _06402_);
  or (_36029_, _36028_, _36025_);
  and (_36030_, _36029_, _07132_);
  or (_36031_, _35956_, _08015_);
  and (_36033_, _36013_, _06306_);
  and (_36034_, _36033_, _36031_);
  or (_36035_, _36034_, _36030_);
  and (_36036_, _36035_, _12514_);
  and (_36037_, _35961_, _06411_);
  and (_36038_, _36037_, _36031_);
  and (_36039_, _35968_, _07124_);
  or (_36040_, _36039_, _06303_);
  or (_36041_, _36040_, _36038_);
  or (_36042_, _36041_, _36036_);
  and (_36044_, _15410_, _07858_);
  or (_36045_, _35956_, _08819_);
  or (_36046_, _36045_, _36044_);
  and (_36047_, _36046_, _36042_);
  or (_36048_, _36047_, _06396_);
  nor (_36049_, _10294_, _13718_);
  or (_36050_, _36049_, _35956_);
  or (_36051_, _36050_, _08824_);
  and (_36052_, _36051_, _12558_);
  and (_36053_, _36052_, _36048_);
  nor (_36055_, _13646_, _13642_);
  or (_36056_, _36055_, _13647_);
  and (_36057_, _36056_, _06417_);
  or (_36058_, _36057_, _07142_);
  or (_36059_, _36058_, _36053_);
  or (_36060_, _35968_, _05846_);
  and (_36061_, _36060_, _06168_);
  and (_36062_, _36061_, _36059_);
  and (_36063_, _36056_, _06167_);
  or (_36064_, _36063_, _06433_);
  or (_36066_, _36064_, _36062_);
  or (_36067_, _35958_, _06829_);
  and (_36068_, _36067_, _07160_);
  and (_36069_, _36068_, _36066_);
  and (_36070_, _35968_, _07577_);
  or (_36071_, _36070_, _06440_);
  or (_36072_, _36071_, _36069_);
  and (_36073_, _15478_, _07858_);
  or (_36074_, _35956_, _06444_);
  or (_36075_, _36074_, _36073_);
  and (_36077_, _36075_, _01317_);
  and (_36078_, _36077_, _36072_);
  or (_36079_, _36078_, _35954_);
  and (_43770_, _36079_, _43100_);
  not (_36080_, \oc8051_golden_model_1.SBUF [0]);
  nor (_36081_, _01317_, _36080_);
  nor (_36082_, _07783_, _36080_);
  nor (_36083_, _08211_, _13750_);
  or (_36084_, _36083_, _36082_);
  or (_36085_, _36084_, _06161_);
  and (_36087_, _07783_, \oc8051_golden_model_1.ACC [0]);
  or (_36088_, _36087_, _36082_);
  and (_36089_, _36088_, _07056_);
  nor (_36090_, _07056_, _36080_);
  or (_36091_, _36090_, _06160_);
  or (_36092_, _36091_, _36089_);
  and (_36093_, _36092_, _07075_);
  and (_36094_, _36093_, _36085_);
  and (_36095_, _07783_, _07049_);
  or (_36096_, _36095_, _36082_);
  and (_36098_, _36096_, _06217_);
  or (_36099_, _36098_, _36094_);
  and (_36100_, _36099_, _06229_);
  and (_36101_, _36088_, _06220_);
  or (_36102_, _36101_, _09842_);
  or (_36103_, _36102_, _36100_);
  or (_36104_, _36096_, _06132_);
  and (_36105_, _36104_, _36103_);
  or (_36106_, _36105_, _06116_);
  and (_36107_, _09160_, _07783_);
  or (_36109_, _36082_, _06117_);
  or (_36110_, _36109_, _36107_);
  and (_36111_, _36110_, _36106_);
  or (_36112_, _36111_, _05787_);
  and (_36113_, _14260_, _07783_);
  or (_36114_, _36082_, _06114_);
  or (_36115_, _36114_, _36113_);
  and (_36116_, _36115_, _06111_);
  and (_36117_, _36116_, _36112_);
  and (_36118_, _07783_, _08708_);
  or (_36120_, _36118_, _36082_);
  and (_36121_, _36120_, _06110_);
  or (_36122_, _36121_, _06297_);
  or (_36123_, _36122_, _36117_);
  and (_36124_, _14275_, _07783_);
  or (_36125_, _36082_, _07127_);
  or (_36126_, _36125_, _36124_);
  and (_36127_, _36126_, _07125_);
  and (_36128_, _36127_, _36123_);
  nor (_36129_, _12321_, _13750_);
  or (_36131_, _36129_, _36082_);
  nand (_36132_, _10276_, _07783_);
  and (_36133_, _36132_, _06402_);
  and (_36134_, _36133_, _36131_);
  or (_36135_, _36134_, _36128_);
  and (_36136_, _36135_, _07132_);
  nand (_36137_, _36120_, _06306_);
  nor (_36138_, _36137_, _36083_);
  or (_36139_, _36138_, _06411_);
  or (_36140_, _36139_, _36136_);
  nor (_36142_, _36082_, _07130_);
  nand (_36143_, _36142_, _36132_);
  and (_36144_, _36143_, _36140_);
  or (_36145_, _36144_, _06303_);
  and (_36146_, _14167_, _07783_);
  or (_36147_, _36082_, _08819_);
  or (_36148_, _36147_, _36146_);
  and (_36149_, _36148_, _08824_);
  and (_36150_, _36149_, _36145_);
  and (_36151_, _36131_, _06396_);
  or (_36153_, _36151_, _19287_);
  or (_36154_, _36153_, _36150_);
  or (_36155_, _36084_, _06630_);
  and (_36156_, _36155_, _01317_);
  and (_36157_, _36156_, _36154_);
  or (_36158_, _36157_, _36081_);
  and (_43772_, _36158_, _43100_);
  not (_36159_, \oc8051_golden_model_1.SBUF [1]);
  nor (_36160_, _01317_, _36159_);
  or (_36161_, _14442_, _13750_);
  or (_36163_, _07783_, \oc8051_golden_model_1.SBUF [1]);
  and (_36164_, _36163_, _05787_);
  and (_36165_, _36164_, _36161_);
  and (_36166_, _09115_, _07783_);
  nor (_36167_, _07783_, _36159_);
  or (_36168_, _36167_, _06117_);
  or (_36169_, _36168_, _36166_);
  and (_36170_, _14363_, _07783_);
  not (_36171_, _36170_);
  and (_36172_, _36171_, _36163_);
  or (_36174_, _36172_, _06161_);
  and (_36175_, _07783_, \oc8051_golden_model_1.ACC [1]);
  or (_36176_, _36175_, _36167_);
  and (_36177_, _36176_, _07056_);
  nor (_36178_, _07056_, _36159_);
  or (_36179_, _36178_, _06160_);
  or (_36180_, _36179_, _36177_);
  and (_36181_, _36180_, _07075_);
  and (_36182_, _36181_, _36174_);
  and (_36183_, _07783_, _07306_);
  or (_36185_, _36183_, _36167_);
  and (_36186_, _36185_, _06217_);
  or (_36187_, _36186_, _36182_);
  and (_36188_, _36187_, _06229_);
  and (_36189_, _36176_, _06220_);
  or (_36190_, _36189_, _09842_);
  or (_36191_, _36190_, _36188_);
  or (_36192_, _36185_, _06132_);
  and (_36193_, _36192_, _36191_);
  or (_36194_, _36193_, _06116_);
  and (_36196_, _36194_, _06114_);
  and (_36197_, _36196_, _36169_);
  or (_36198_, _36197_, _36165_);
  and (_36199_, _36198_, _06298_);
  or (_36200_, _14346_, _13750_);
  and (_36201_, _36163_, _06297_);
  and (_36202_, _36201_, _36200_);
  nand (_36203_, _07783_, _06945_);
  and (_36204_, _36163_, _06110_);
  and (_36205_, _36204_, _36203_);
  or (_36207_, _36205_, _06402_);
  or (_36208_, _36207_, _36202_);
  or (_36209_, _36208_, _36199_);
  nor (_36210_, _10277_, _13750_);
  or (_36211_, _36210_, _36167_);
  nand (_36212_, _10275_, _07783_);
  and (_36213_, _36212_, _36211_);
  or (_36214_, _36213_, _07125_);
  and (_36215_, _36214_, _07132_);
  and (_36216_, _36215_, _36209_);
  or (_36218_, _14344_, _13750_);
  and (_36219_, _36163_, _06306_);
  and (_36220_, _36219_, _36218_);
  or (_36221_, _36220_, _06411_);
  or (_36222_, _36221_, _36216_);
  nor (_36223_, _36167_, _07130_);
  nand (_36224_, _36223_, _36212_);
  and (_36225_, _36224_, _08819_);
  and (_36226_, _36225_, _36222_);
  or (_36227_, _36203_, _08176_);
  and (_36229_, _36163_, _06303_);
  and (_36230_, _36229_, _36227_);
  or (_36231_, _36230_, _06396_);
  or (_36232_, _36231_, _36226_);
  or (_36233_, _36211_, _08824_);
  and (_36234_, _36233_, _36232_);
  and (_36235_, _36234_, _06829_);
  and (_36236_, _36172_, _06433_);
  or (_36237_, _36236_, _06440_);
  or (_36238_, _36237_, _36235_);
  or (_36240_, _36167_, _06444_);
  or (_36241_, _36240_, _36170_);
  and (_36242_, _36241_, _01317_);
  and (_36243_, _36242_, _36238_);
  or (_36244_, _36243_, _36160_);
  and (_43773_, _36244_, _43100_);
  and (_36245_, _01321_, \oc8051_golden_model_1.SBUF [2]);
  and (_36246_, _13750_, \oc8051_golden_model_1.SBUF [2]);
  or (_36247_, _36246_, _08248_);
  and (_36248_, _07783_, _08768_);
  or (_36250_, _36248_, _36246_);
  and (_36251_, _36250_, _06306_);
  and (_36252_, _36251_, _36247_);
  and (_36253_, _09211_, _07783_);
  or (_36254_, _36253_, _36246_);
  and (_36255_, _36254_, _06116_);
  and (_36256_, _14542_, _07783_);
  or (_36257_, _36256_, _36246_);
  or (_36258_, _36257_, _06161_);
  and (_36259_, _07783_, \oc8051_golden_model_1.ACC [2]);
  or (_36261_, _36259_, _36246_);
  and (_36262_, _36261_, _07056_);
  and (_36263_, _07057_, \oc8051_golden_model_1.SBUF [2]);
  or (_36264_, _36263_, _06160_);
  or (_36265_, _36264_, _36262_);
  and (_36266_, _36265_, _07075_);
  and (_36267_, _36266_, _36258_);
  and (_36268_, _07783_, _07708_);
  or (_36269_, _36268_, _36246_);
  and (_36270_, _36269_, _06217_);
  or (_36272_, _36270_, _36267_);
  and (_36273_, _36272_, _06229_);
  and (_36274_, _36261_, _06220_);
  or (_36275_, _36274_, _09842_);
  or (_36276_, _36275_, _36273_);
  or (_36277_, _36269_, _06132_);
  and (_36278_, _36277_, _06117_);
  and (_36279_, _36278_, _36276_);
  or (_36280_, _36279_, _05787_);
  or (_36281_, _36280_, _36255_);
  and (_36283_, _14630_, _07783_);
  or (_36284_, _36283_, _36246_);
  or (_36285_, _36284_, _06114_);
  and (_36286_, _36285_, _06111_);
  and (_36287_, _36286_, _36281_);
  and (_36288_, _36250_, _06110_);
  or (_36289_, _36288_, _06297_);
  or (_36290_, _36289_, _36287_);
  and (_36291_, _14646_, _07783_);
  or (_36292_, _36246_, _07127_);
  or (_36294_, _36292_, _36291_);
  and (_36295_, _36294_, _07125_);
  and (_36296_, _36295_, _36290_);
  and (_36297_, _10282_, _07783_);
  or (_36298_, _36297_, _36246_);
  and (_36299_, _36298_, _06402_);
  or (_36300_, _36299_, _36296_);
  and (_36301_, _36300_, _07132_);
  or (_36302_, _36301_, _36252_);
  and (_36303_, _36302_, _07130_);
  and (_36305_, _36261_, _06411_);
  and (_36306_, _36305_, _36247_);
  or (_36307_, _36306_, _06303_);
  or (_36308_, _36307_, _36303_);
  and (_36309_, _14643_, _07783_);
  or (_36310_, _36246_, _08819_);
  or (_36311_, _36310_, _36309_);
  and (_36312_, _36311_, _08824_);
  and (_36313_, _36312_, _36308_);
  nor (_36314_, _10281_, _13750_);
  or (_36316_, _36314_, _36246_);
  and (_36317_, _36316_, _06396_);
  or (_36318_, _36317_, _36313_);
  and (_36319_, _36318_, _06829_);
  and (_36320_, _36257_, _06433_);
  or (_36321_, _36320_, _06440_);
  or (_36322_, _36321_, _36319_);
  and (_36323_, _14710_, _07783_);
  or (_36324_, _36246_, _06444_);
  or (_36325_, _36324_, _36323_);
  and (_36327_, _36325_, _01317_);
  and (_36328_, _36327_, _36322_);
  or (_36329_, _36328_, _36245_);
  and (_43774_, _36329_, _43100_);
  and (_36330_, _13750_, \oc8051_golden_model_1.SBUF [3]);
  or (_36331_, _36330_, _08140_);
  and (_36332_, _07783_, _08712_);
  or (_36333_, _36332_, _36330_);
  and (_36334_, _36333_, _06306_);
  and (_36335_, _36334_, _36331_);
  and (_36337_, _14738_, _07783_);
  or (_36338_, _36337_, _36330_);
  or (_36339_, _36338_, _06161_);
  and (_36340_, _07783_, \oc8051_golden_model_1.ACC [3]);
  or (_36341_, _36340_, _36330_);
  and (_36342_, _36341_, _07056_);
  and (_36343_, _07057_, \oc8051_golden_model_1.SBUF [3]);
  or (_36344_, _36343_, _06160_);
  or (_36345_, _36344_, _36342_);
  and (_36346_, _36345_, _07075_);
  and (_36348_, _36346_, _36339_);
  and (_36349_, _07783_, _07544_);
  or (_36350_, _36349_, _36330_);
  and (_36351_, _36350_, _06217_);
  or (_36352_, _36351_, _36348_);
  and (_36353_, _36352_, _06229_);
  and (_36354_, _36341_, _06220_);
  or (_36355_, _36354_, _09842_);
  or (_36356_, _36355_, _36353_);
  and (_36357_, _36350_, _06117_);
  or (_36359_, _36357_, _06133_);
  and (_36360_, _36359_, _36356_);
  and (_36361_, _09210_, _07783_);
  or (_36362_, _36361_, _36330_);
  and (_36363_, _36362_, _06116_);
  or (_36364_, _36363_, _05787_);
  or (_36365_, _36364_, _36360_);
  and (_36366_, _14825_, _07783_);
  or (_36367_, _36330_, _06114_);
  or (_36368_, _36367_, _36366_);
  and (_36370_, _36368_, _06111_);
  and (_36371_, _36370_, _36365_);
  and (_36372_, _36333_, _06110_);
  or (_36373_, _36372_, _06297_);
  or (_36374_, _36373_, _36371_);
  and (_36375_, _14727_, _07783_);
  or (_36376_, _36330_, _07127_);
  or (_36377_, _36376_, _36375_);
  and (_36378_, _36377_, _07125_);
  and (_36379_, _36378_, _36374_);
  and (_36381_, _12318_, _07783_);
  or (_36382_, _36381_, _36330_);
  and (_36383_, _36382_, _06402_);
  or (_36384_, _36383_, _36379_);
  and (_36385_, _36384_, _07132_);
  or (_36386_, _36385_, _36335_);
  and (_36387_, _36386_, _07130_);
  and (_36388_, _36341_, _06411_);
  and (_36389_, _36388_, _36331_);
  or (_36390_, _36389_, _06303_);
  or (_36392_, _36390_, _36387_);
  and (_36393_, _14724_, _07783_);
  or (_36394_, _36330_, _08819_);
  or (_36395_, _36394_, _36393_);
  and (_36396_, _36395_, _08824_);
  and (_36397_, _36396_, _36392_);
  nor (_36398_, _10273_, _13750_);
  or (_36399_, _36398_, _36330_);
  and (_36400_, _36399_, _06396_);
  or (_36401_, _36400_, _06433_);
  or (_36403_, _36401_, _36397_);
  or (_36404_, _36338_, _06829_);
  and (_36405_, _36404_, _06444_);
  and (_36406_, _36405_, _36403_);
  and (_36407_, _14897_, _07783_);
  or (_36408_, _36407_, _36330_);
  and (_36409_, _36408_, _06440_);
  or (_36410_, _36409_, _01321_);
  or (_36411_, _36410_, _36406_);
  or (_36412_, _01317_, \oc8051_golden_model_1.SBUF [3]);
  and (_36414_, _36412_, _43100_);
  and (_43775_, _36414_, _36411_);
  and (_36415_, _13750_, \oc8051_golden_model_1.SBUF [4]);
  and (_36416_, _14928_, _07783_);
  or (_36417_, _36416_, _36415_);
  or (_36418_, _36417_, _06161_);
  and (_36419_, _07783_, \oc8051_golden_model_1.ACC [4]);
  or (_36420_, _36419_, _36415_);
  and (_36421_, _36420_, _07056_);
  and (_36422_, _07057_, \oc8051_golden_model_1.SBUF [4]);
  or (_36423_, _36422_, _06160_);
  or (_36424_, _36423_, _36421_);
  and (_36425_, _36424_, _07075_);
  and (_36426_, _36425_, _36418_);
  and (_36427_, _08336_, _07783_);
  or (_36428_, _36427_, _36415_);
  and (_36429_, _36428_, _06217_);
  or (_36430_, _36429_, _36426_);
  and (_36431_, _36430_, _06229_);
  and (_36432_, _36420_, _06220_);
  or (_36434_, _36432_, _09842_);
  or (_36435_, _36434_, _36431_);
  or (_36436_, _36428_, _06132_);
  and (_36437_, _36436_, _36435_);
  or (_36438_, _36437_, _06116_);
  and (_36439_, _09209_, _07783_);
  or (_36440_, _36415_, _06117_);
  or (_36441_, _36440_, _36439_);
  and (_36442_, _36441_, _06114_);
  and (_36443_, _36442_, _36438_);
  and (_36445_, _15013_, _07783_);
  or (_36446_, _36445_, _36415_);
  and (_36447_, _36446_, _05787_);
  or (_36448_, _36447_, _36443_);
  or (_36449_, _36448_, _11136_);
  and (_36450_, _15029_, _07783_);
  or (_36451_, _36415_, _07127_);
  or (_36452_, _36451_, _36450_);
  and (_36453_, _08715_, _07783_);
  or (_36454_, _36453_, _36415_);
  or (_36456_, _36454_, _06111_);
  and (_36457_, _36456_, _07125_);
  and (_36458_, _36457_, _36452_);
  and (_36459_, _36458_, _36449_);
  and (_36460_, _10289_, _07783_);
  or (_36461_, _36460_, _36415_);
  and (_36462_, _36461_, _06402_);
  or (_36463_, _36462_, _36459_);
  and (_36464_, _36463_, _07132_);
  or (_36465_, _36415_, _08339_);
  and (_36467_, _36454_, _06306_);
  and (_36468_, _36467_, _36465_);
  or (_36469_, _36468_, _36464_);
  and (_36470_, _36469_, _07130_);
  and (_36471_, _36420_, _06411_);
  and (_36472_, _36471_, _36465_);
  or (_36473_, _36472_, _06303_);
  or (_36474_, _36473_, _36470_);
  and (_36475_, _15026_, _07783_);
  or (_36476_, _36415_, _08819_);
  or (_36478_, _36476_, _36475_);
  and (_36479_, _36478_, _08824_);
  and (_36480_, _36479_, _36474_);
  nor (_36481_, _10288_, _13750_);
  or (_36482_, _36481_, _36415_);
  and (_36483_, _36482_, _06396_);
  or (_36484_, _36483_, _06433_);
  or (_36485_, _36484_, _36480_);
  or (_36486_, _36417_, _06829_);
  and (_36487_, _36486_, _06444_);
  and (_36489_, _36487_, _36485_);
  and (_36490_, _15087_, _07783_);
  or (_36491_, _36490_, _36415_);
  and (_36492_, _36491_, _06440_);
  or (_36493_, _36492_, _01321_);
  or (_36494_, _36493_, _36489_);
  or (_36495_, _01317_, \oc8051_golden_model_1.SBUF [4]);
  and (_36496_, _36495_, _43100_);
  and (_43776_, _36496_, _36494_);
  and (_36497_, _13750_, \oc8051_golden_model_1.SBUF [5]);
  or (_36499_, _36497_, _08104_);
  and (_36500_, _08736_, _07783_);
  or (_36501_, _36500_, _36497_);
  and (_36502_, _36501_, _06306_);
  and (_36503_, _36502_, _36499_);
  and (_36504_, _15119_, _07783_);
  or (_36505_, _36504_, _36497_);
  or (_36506_, _36505_, _06161_);
  and (_36507_, _07783_, \oc8051_golden_model_1.ACC [5]);
  or (_36508_, _36507_, _36497_);
  and (_36510_, _36508_, _07056_);
  and (_36511_, _07057_, \oc8051_golden_model_1.SBUF [5]);
  or (_36512_, _36511_, _06160_);
  or (_36513_, _36512_, _36510_);
  and (_36514_, _36513_, _07075_);
  and (_36515_, _36514_, _36506_);
  and (_36516_, _08101_, _07783_);
  or (_36517_, _36516_, _36497_);
  and (_36518_, _36517_, _06217_);
  or (_36519_, _36518_, _36515_);
  and (_36521_, _36519_, _06229_);
  and (_36522_, _36508_, _06220_);
  or (_36523_, _36522_, _09842_);
  or (_36524_, _36523_, _36521_);
  or (_36525_, _36517_, _06132_);
  and (_36526_, _36525_, _36524_);
  or (_36527_, _36526_, _06116_);
  and (_36528_, _09208_, _07783_);
  or (_36529_, _36497_, _06117_);
  or (_36530_, _36529_, _36528_);
  and (_36532_, _36530_, _06114_);
  and (_36533_, _36532_, _36527_);
  and (_36534_, _15203_, _07783_);
  or (_36535_, _36534_, _36497_);
  and (_36536_, _36535_, _05787_);
  or (_36537_, _36536_, _11136_);
  or (_36538_, _36537_, _36533_);
  and (_36539_, _15219_, _07783_);
  or (_36540_, _36497_, _07127_);
  or (_36541_, _36540_, _36539_);
  or (_36543_, _36501_, _06111_);
  and (_36544_, _36543_, _07125_);
  and (_36545_, _36544_, _36541_);
  and (_36546_, _36545_, _36538_);
  and (_36547_, _12325_, _07783_);
  or (_36548_, _36547_, _36497_);
  and (_36549_, _36548_, _06402_);
  or (_36550_, _36549_, _36546_);
  and (_36551_, _36550_, _07132_);
  or (_36552_, _36551_, _36503_);
  and (_36554_, _36552_, _07130_);
  and (_36555_, _36508_, _06411_);
  and (_36556_, _36555_, _36499_);
  or (_36557_, _36556_, _06303_);
  or (_36558_, _36557_, _36554_);
  and (_36559_, _15216_, _07783_);
  or (_36560_, _36497_, _08819_);
  or (_36561_, _36560_, _36559_);
  and (_36562_, _36561_, _08824_);
  and (_36563_, _36562_, _36558_);
  nor (_36565_, _10269_, _13750_);
  or (_36566_, _36565_, _36497_);
  and (_36567_, _36566_, _06396_);
  or (_36568_, _36567_, _06433_);
  or (_36569_, _36568_, _36563_);
  or (_36570_, _36505_, _06829_);
  and (_36571_, _36570_, _06444_);
  and (_36572_, _36571_, _36569_);
  and (_36573_, _15275_, _07783_);
  or (_36574_, _36573_, _36497_);
  and (_36576_, _36574_, _06440_);
  or (_36577_, _36576_, _01321_);
  or (_36578_, _36577_, _36572_);
  or (_36579_, _01317_, \oc8051_golden_model_1.SBUF [5]);
  and (_36580_, _36579_, _43100_);
  and (_43777_, _36580_, _36578_);
  and (_36581_, _13750_, \oc8051_golden_model_1.SBUF [6]);
  and (_36582_, _15300_, _07783_);
  or (_36583_, _36582_, _36581_);
  or (_36584_, _36583_, _06161_);
  and (_36586_, _07783_, \oc8051_golden_model_1.ACC [6]);
  or (_36587_, _36586_, _36581_);
  and (_36588_, _36587_, _07056_);
  and (_36589_, _07057_, \oc8051_golden_model_1.SBUF [6]);
  or (_36590_, _36589_, _06160_);
  or (_36591_, _36590_, _36588_);
  and (_36592_, _36591_, _07075_);
  and (_36593_, _36592_, _36584_);
  and (_36594_, _08012_, _07783_);
  or (_36595_, _36594_, _36581_);
  and (_36597_, _36595_, _06217_);
  or (_36598_, _36597_, _36593_);
  and (_36599_, _36598_, _06229_);
  and (_36600_, _36587_, _06220_);
  or (_36601_, _36600_, _09842_);
  or (_36602_, _36601_, _36599_);
  or (_36603_, _36595_, _06132_);
  and (_36604_, _36603_, _36602_);
  or (_36605_, _36604_, _06116_);
  and (_36606_, _09207_, _07783_);
  or (_36608_, _36581_, _06117_);
  or (_36609_, _36608_, _36606_);
  and (_36610_, _36609_, _06114_);
  and (_36611_, _36610_, _36605_);
  and (_36612_, _15395_, _07783_);
  or (_36613_, _36612_, _36581_);
  and (_36614_, _36613_, _05787_);
  or (_36615_, _36614_, _11136_);
  or (_36616_, _36615_, _36611_);
  and (_36617_, _15413_, _07783_);
  or (_36619_, _36581_, _07127_);
  or (_36620_, _36619_, _36617_);
  and (_36621_, _15402_, _07783_);
  or (_36622_, _36621_, _36581_);
  or (_36623_, _36622_, _06111_);
  and (_36624_, _36623_, _07125_);
  and (_36625_, _36624_, _36620_);
  and (_36626_, _36625_, _36616_);
  and (_36627_, _10295_, _07783_);
  or (_36628_, _36627_, _36581_);
  and (_36630_, _36628_, _06402_);
  or (_36631_, _36630_, _36626_);
  and (_36632_, _36631_, _07132_);
  or (_36633_, _36581_, _08015_);
  and (_36634_, _36622_, _06306_);
  and (_36635_, _36634_, _36633_);
  or (_36636_, _36635_, _36632_);
  and (_36637_, _36636_, _07130_);
  and (_36638_, _36587_, _06411_);
  and (_36639_, _36638_, _36633_);
  or (_36641_, _36639_, _06303_);
  or (_36642_, _36641_, _36637_);
  and (_36643_, _15410_, _07783_);
  or (_36644_, _36581_, _08819_);
  or (_36645_, _36644_, _36643_);
  and (_36646_, _36645_, _08824_);
  and (_36647_, _36646_, _36642_);
  nor (_36648_, _10294_, _13750_);
  or (_36649_, _36648_, _36581_);
  and (_36650_, _36649_, _06396_);
  or (_36652_, _36650_, _06433_);
  or (_36653_, _36652_, _36647_);
  or (_36654_, _36583_, _06829_);
  and (_36655_, _36654_, _06444_);
  and (_36656_, _36655_, _36653_);
  and (_36657_, _15478_, _07783_);
  or (_36658_, _36657_, _36581_);
  and (_36659_, _36658_, _06440_);
  or (_36660_, _36659_, _01321_);
  or (_36661_, _36660_, _36656_);
  or (_36663_, _01317_, \oc8051_golden_model_1.SBUF [6]);
  and (_36664_, _36663_, _43100_);
  and (_43778_, _36664_, _36661_);
  not (_36665_, \oc8051_golden_model_1.PSW [0]);
  nor (_36666_, _01317_, _36665_);
  nand (_36667_, _10276_, _07794_);
  nor (_36668_, _07794_, _36665_);
  nor (_36669_, _36668_, _07130_);
  nand (_36670_, _36669_, _36667_);
  nor (_36671_, _08404_, _36665_);
  and (_36673_, _14169_, _08404_);
  or (_36674_, _36673_, _36671_);
  or (_36675_, _36674_, _06157_);
  nor (_36676_, _08211_, _14076_);
  or (_36677_, _36676_, _36668_);
  and (_36678_, _36677_, _06160_);
  nor (_36679_, _07056_, _36665_);
  and (_36680_, _07794_, \oc8051_golden_model_1.ACC [0]);
  or (_36681_, _36680_, _36668_);
  and (_36682_, _36681_, _07056_);
  or (_36684_, _36682_, _36679_);
  and (_36685_, _36684_, _06161_);
  or (_36686_, _36685_, _06156_);
  or (_36687_, _36686_, _36678_);
  and (_36688_, _36687_, _36675_);
  and (_36689_, _36688_, _07075_);
  and (_36690_, _07794_, _07049_);
  or (_36691_, _36690_, _36668_);
  and (_36692_, _36691_, _06217_);
  or (_36693_, _36692_, _06220_);
  or (_36695_, _36693_, _36689_);
  or (_36696_, _36681_, _06229_);
  and (_36697_, _36696_, _06153_);
  and (_36698_, _36697_, _36695_);
  and (_36699_, _36668_, _06152_);
  or (_36700_, _36699_, _06145_);
  or (_36701_, _36700_, _36698_);
  or (_36702_, _36677_, _06146_);
  and (_36703_, _36702_, _06140_);
  and (_36704_, _36703_, _36701_);
  or (_36706_, _36671_, _14170_);
  and (_36707_, _36706_, _06139_);
  and (_36708_, _36707_, _36674_);
  or (_36709_, _36708_, _09842_);
  or (_36710_, _36709_, _36704_);
  or (_36711_, _36691_, _06132_);
  and (_36712_, _36711_, _36710_);
  or (_36713_, _36712_, _06116_);
  and (_36714_, _09160_, _07794_);
  or (_36715_, _36668_, _06117_);
  or (_36717_, _36715_, _36714_);
  and (_36718_, _36717_, _06114_);
  and (_36719_, _36718_, _36713_);
  and (_36720_, _14260_, _07794_);
  or (_36721_, _36720_, _36668_);
  and (_36722_, _36721_, _05787_);
  or (_36723_, _36722_, _36719_);
  or (_36724_, _36723_, _11136_);
  and (_36725_, _14275_, _07794_);
  or (_36726_, _36668_, _07127_);
  or (_36728_, _36726_, _36725_);
  and (_36729_, _07794_, _08708_);
  or (_36730_, _36729_, _36668_);
  or (_36731_, _36730_, _06111_);
  and (_36732_, _36731_, _07125_);
  and (_36733_, _36732_, _36728_);
  and (_36734_, _36733_, _36724_);
  nor (_36735_, _12321_, _14076_);
  or (_36736_, _36735_, _36668_);
  and (_36737_, _36667_, _06402_);
  and (_36739_, _36737_, _36736_);
  or (_36740_, _36739_, _36734_);
  and (_36741_, _36740_, _07132_);
  nand (_36742_, _36730_, _06306_);
  nor (_36743_, _36742_, _36676_);
  or (_36744_, _36743_, _06411_);
  or (_36745_, _36744_, _36741_);
  and (_36746_, _36745_, _36670_);
  or (_36747_, _36746_, _06303_);
  and (_36748_, _14167_, _07794_);
  or (_36750_, _36668_, _08819_);
  or (_36751_, _36750_, _36748_);
  and (_36752_, _36751_, _08824_);
  and (_36753_, _36752_, _36747_);
  and (_36754_, _36736_, _06396_);
  or (_36755_, _36754_, _06433_);
  or (_36756_, _36755_, _36753_);
  or (_36757_, _36677_, _06829_);
  and (_36758_, _36757_, _36756_);
  or (_36759_, _36758_, _05748_);
  or (_36761_, _36668_, _05749_);
  and (_36762_, _36761_, _36759_);
  or (_36763_, _36762_, _06440_);
  or (_36764_, _36677_, _06444_);
  and (_36765_, _36764_, _01317_);
  and (_36766_, _36765_, _36763_);
  or (_36767_, _36766_, _36666_);
  and (_43779_, _36767_, _43100_);
  not (_36768_, \oc8051_golden_model_1.PSW [1]);
  nor (_36769_, _01317_, _36768_);
  or (_36771_, _14442_, _14076_);
  or (_36772_, _07794_, \oc8051_golden_model_1.PSW [1]);
  and (_36773_, _36772_, _05787_);
  and (_36774_, _36773_, _36771_);
  nor (_36775_, _07794_, _36768_);
  and (_36776_, _07794_, _07306_);
  or (_36777_, _36776_, _36775_);
  or (_36778_, _36777_, _07075_);
  and (_36779_, _14363_, _07794_);
  not (_36780_, _36779_);
  and (_36782_, _36780_, _36772_);
  or (_36783_, _36782_, _06161_);
  and (_36784_, _07794_, \oc8051_golden_model_1.ACC [1]);
  or (_36785_, _36784_, _36775_);
  and (_36786_, _36785_, _07056_);
  nor (_36787_, _07056_, _36768_);
  or (_36788_, _36787_, _06160_);
  or (_36789_, _36788_, _36786_);
  and (_36790_, _36789_, _06157_);
  and (_36791_, _36790_, _36783_);
  nor (_36793_, _08404_, _36768_);
  and (_36794_, _14367_, _08404_);
  or (_36795_, _36794_, _36793_);
  and (_36796_, _36795_, _06156_);
  or (_36797_, _36796_, _06217_);
  or (_36798_, _36797_, _36791_);
  and (_36799_, _36798_, _36778_);
  or (_36800_, _36799_, _06220_);
  or (_36801_, _36785_, _06229_);
  and (_36802_, _36801_, _06153_);
  and (_36804_, _36802_, _36800_);
  and (_36805_, _14349_, _08404_);
  or (_36806_, _36805_, _36793_);
  and (_36807_, _36806_, _06152_);
  or (_36808_, _36807_, _06145_);
  or (_36809_, _36808_, _36804_);
  and (_36810_, _36794_, _14382_);
  or (_36811_, _36793_, _06146_);
  or (_36812_, _36811_, _36810_);
  and (_36813_, _36812_, _36809_);
  and (_36815_, _36813_, _06140_);
  and (_36816_, _14351_, _08404_);
  or (_36817_, _36793_, _36816_);
  and (_36818_, _36817_, _06139_);
  or (_36819_, _36818_, _09842_);
  or (_36820_, _36819_, _36815_);
  or (_36821_, _36777_, _06132_);
  and (_36822_, _36821_, _36820_);
  or (_36823_, _36822_, _06116_);
  and (_36824_, _09115_, _07794_);
  or (_36826_, _36775_, _06117_);
  or (_36827_, _36826_, _36824_);
  and (_36828_, _36827_, _06114_);
  and (_36829_, _36828_, _36823_);
  or (_36830_, _36829_, _36774_);
  and (_36831_, _36830_, _06298_);
  or (_36832_, _14346_, _14076_);
  and (_36833_, _36772_, _06297_);
  and (_36834_, _36833_, _36832_);
  nand (_36835_, _07794_, _06945_);
  and (_36837_, _36835_, _06110_);
  and (_36838_, _36837_, _36772_);
  or (_36839_, _36838_, _06402_);
  or (_36840_, _36839_, _36834_);
  or (_36841_, _36840_, _36831_);
  nor (_36842_, _10277_, _14076_);
  or (_36843_, _36842_, _36775_);
  nand (_36844_, _10275_, _07794_);
  and (_36845_, _36844_, _36843_);
  or (_36846_, _36845_, _07125_);
  and (_36848_, _36846_, _07132_);
  and (_36849_, _36848_, _36841_);
  or (_36850_, _14344_, _14076_);
  and (_36851_, _36772_, _06306_);
  and (_36852_, _36851_, _36850_);
  or (_36853_, _36852_, _06411_);
  or (_36854_, _36853_, _36849_);
  nor (_36855_, _36775_, _07130_);
  nand (_36856_, _36855_, _36844_);
  and (_36857_, _36856_, _08819_);
  and (_36859_, _36857_, _36854_);
  or (_36860_, _36835_, _08176_);
  and (_36861_, _36772_, _06303_);
  and (_36862_, _36861_, _36860_);
  or (_36863_, _36862_, _06396_);
  or (_36864_, _36863_, _36859_);
  or (_36865_, _36843_, _08824_);
  and (_36866_, _36865_, _36864_);
  or (_36867_, _36866_, _06433_);
  or (_36868_, _36782_, _06829_);
  and (_36870_, _36868_, _05749_);
  and (_36871_, _36870_, _36867_);
  and (_36872_, _36806_, _05748_);
  or (_36873_, _36872_, _06440_);
  or (_36874_, _36873_, _36871_);
  or (_36875_, _36775_, _06444_);
  or (_36876_, _36875_, _36779_);
  and (_36877_, _36876_, _01317_);
  and (_36878_, _36877_, _36874_);
  or (_36879_, _36878_, _36769_);
  and (_43780_, _36879_, _43100_);
  and (_36881_, _01321_, \oc8051_golden_model_1.PSW [2]);
  or (_36882_, _14118_, _11038_);
  or (_36883_, _11039_, _10781_);
  and (_36884_, _36883_, _36882_);
  and (_36885_, _36884_, _17199_);
  nor (_36886_, _10657_, _06172_);
  or (_36887_, _36886_, \oc8051_golden_model_1.ACC [7]);
  nor (_36888_, _10657_, _14131_);
  not (_36889_, _36888_);
  and (_36891_, _36889_, _36887_);
  not (_36892_, _36891_);
  or (_36893_, _36892_, _14100_);
  and (_36894_, _36889_, _10951_);
  and (_36895_, _36894_, _36893_);
  and (_36896_, _36888_, _10948_);
  or (_36897_, _36896_, _36895_);
  and (_36898_, _36897_, _10895_);
  and (_36899_, _06122_, _06300_);
  not (_36900_, _36899_);
  not (_36902_, _10765_);
  nor (_36903_, _36902_, _10302_);
  nor (_36904_, _10303_, \oc8051_golden_model_1.ACC [7]);
  nor (_36905_, _36903_, _36904_);
  not (_36906_, _36905_);
  nor (_36907_, _36906_, _14087_);
  nor (_36908_, _36907_, _36903_);
  and (_36909_, _36908_, _10370_);
  and (_36910_, _36903_, _10367_);
  or (_36911_, _36910_, _36909_);
  or (_36913_, _36911_, _36900_);
  and (_36914_, _14076_, \oc8051_golden_model_1.PSW [2]);
  and (_36915_, _14630_, _07794_);
  or (_36916_, _36915_, _36914_);
  and (_36917_, _36916_, _05787_);
  and (_36918_, _07794_, _07708_);
  or (_36919_, _36918_, _36914_);
  or (_36920_, _36919_, _06132_);
  and (_36921_, _10584_, \oc8051_golden_model_1.ACC [7]);
  nor (_36922_, _10584_, \oc8051_golden_model_1.ACC [7]);
  or (_36924_, _36922_, _36921_);
  and (_36925_, _36924_, _14007_);
  nor (_36926_, _36924_, _14007_);
  nor (_36927_, _36926_, _36925_);
  not (_36928_, _36927_);
  nor (_36929_, _36928_, _10646_);
  and (_36930_, _36928_, _10646_);
  or (_36931_, _36930_, _12380_);
  or (_36932_, _36931_, _36929_);
  or (_36933_, _36906_, _13995_);
  nand (_36935_, _36906_, _13995_);
  and (_36936_, _36935_, _36933_);
  and (_36937_, _36936_, _10577_);
  nor (_36938_, _36936_, _10577_);
  or (_36939_, _36938_, _36937_);
  and (_36940_, _36939_, _10557_);
  not (_36941_, _08404_);
  and (_36942_, _36941_, \oc8051_golden_model_1.PSW [2]);
  and (_36943_, _14536_, _08404_);
  or (_36944_, _36943_, _36942_);
  and (_36946_, _36944_, _06152_);
  or (_36947_, _36919_, _07075_);
  and (_36948_, _14542_, _07794_);
  or (_36949_, _36948_, _36914_);
  or (_36950_, _36949_, _06161_);
  and (_36951_, _07794_, \oc8051_golden_model_1.ACC [2]);
  or (_36952_, _36951_, _36914_);
  and (_36953_, _36952_, _07056_);
  and (_36954_, _07057_, \oc8051_golden_model_1.PSW [2]);
  or (_36955_, _36954_, _06160_);
  or (_36957_, _36955_, _36953_);
  and (_36958_, _36957_, _06157_);
  and (_36959_, _36958_, _36950_);
  and (_36960_, _14538_, _08404_);
  or (_36961_, _36960_, _36942_);
  and (_36962_, _36961_, _06156_);
  or (_36963_, _36962_, _06217_);
  or (_36964_, _36963_, _36959_);
  and (_36965_, _36964_, _36947_);
  or (_36966_, _36965_, _06220_);
  or (_36968_, _36952_, _06229_);
  and (_36969_, _36968_, _06153_);
  and (_36970_, _36969_, _36966_);
  or (_36971_, _36970_, _36946_);
  and (_36972_, _36971_, _06146_);
  and (_36973_, _36960_, _14569_);
  or (_36974_, _36973_, _36942_);
  and (_36975_, _36974_, _06145_);
  or (_36976_, _36975_, _09295_);
  or (_36977_, _36976_, _36972_);
  or (_36979_, _16326_, _16210_);
  or (_36980_, _36979_, _16438_);
  or (_36981_, _36980_, _16556_);
  or (_36982_, _36981_, _16673_);
  or (_36983_, _36982_, _16790_);
  or (_36984_, _36983_, _09838_);
  or (_36985_, _36984_, _16908_);
  and (_36986_, _36985_, _10554_);
  and (_36987_, _36986_, _36977_);
  or (_36988_, _36987_, _12379_);
  or (_36990_, _36988_, _36940_);
  and (_36991_, _36990_, _06265_);
  and (_36992_, _36991_, _36932_);
  nor (_36993_, _10396_, \oc8051_golden_model_1.ACC [7]);
  nor (_36994_, _10395_, _14125_);
  nor (_36995_, _36994_, _36993_);
  nor (_36996_, _36995_, _10401_);
  nor (_36997_, _14017_, _10397_);
  or (_36998_, _36997_, _36996_);
  or (_36999_, _36998_, _10450_);
  nand (_37001_, _36998_, _10450_);
  and (_37002_, _37001_, _06260_);
  and (_37003_, _37002_, _36999_);
  or (_37004_, _37003_, _10387_);
  or (_37005_, _37004_, _36992_);
  and (_37006_, _36891_, _14027_);
  nor (_37007_, _36891_, _14027_);
  nor (_37008_, _37007_, _37006_);
  and (_37009_, _37008_, _10719_);
  nor (_37010_, _37008_, _10719_);
  or (_37012_, _37010_, _37009_);
  or (_37013_, _37012_, _10388_);
  and (_37014_, _37013_, _06140_);
  and (_37015_, _37014_, _37005_);
  and (_37016_, _14583_, _08404_);
  or (_37017_, _37016_, _36942_);
  and (_37018_, _37017_, _06139_);
  or (_37019_, _37018_, _09842_);
  or (_37020_, _37019_, _37015_);
  and (_37021_, _37020_, _36920_);
  or (_37023_, _37021_, _06116_);
  and (_37024_, _09211_, _07794_);
  or (_37025_, _36914_, _06117_);
  or (_37026_, _37025_, _37024_);
  and (_37027_, _37026_, _06114_);
  and (_37028_, _37027_, _37023_);
  or (_37029_, _37028_, _36917_);
  and (_37030_, _37029_, _09861_);
  nor (_37031_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and (_37032_, _37031_, _09882_);
  nand (_37034_, _37032_, _09855_);
  nand (_37035_, _37034_, _06298_);
  or (_37036_, _37035_, _37030_);
  and (_37037_, _14646_, _07794_);
  or (_37038_, _36914_, _07127_);
  or (_37039_, _37038_, _37037_);
  and (_37040_, _07794_, _08768_);
  or (_37041_, _37040_, _36914_);
  or (_37042_, _37041_, _06111_);
  and (_37043_, _37042_, _07125_);
  and (_37045_, _37043_, _37039_);
  and (_37046_, _37045_, _37036_);
  and (_37047_, _10282_, _07794_);
  or (_37048_, _37047_, _36914_);
  and (_37049_, _37048_, _06402_);
  or (_37050_, _37049_, _37046_);
  and (_37051_, _37050_, _07132_);
  or (_37052_, _36914_, _08248_);
  and (_37053_, _37041_, _06306_);
  and (_37054_, _37053_, _37052_);
  or (_37056_, _37054_, _37051_);
  and (_37057_, _37056_, _07130_);
  and (_37058_, _36952_, _06411_);
  and (_37059_, _37058_, _37052_);
  or (_37060_, _37059_, _06303_);
  or (_37061_, _37060_, _37057_);
  and (_37062_, _14643_, _07794_);
  or (_37063_, _36914_, _08819_);
  or (_37064_, _37063_, _37062_);
  and (_37065_, _37064_, _08824_);
  and (_37067_, _37065_, _37061_);
  nor (_37068_, _10281_, _14076_);
  or (_37069_, _37068_, _36914_);
  and (_37070_, _37069_, _06396_);
  or (_37071_, _37070_, _36899_);
  or (_37072_, _37071_, _37067_);
  nand (_37073_, _37072_, _36913_);
  and (_37074_, _06288_, _06300_);
  nor (_37075_, _37074_, _06976_);
  nand (_37076_, _37075_, _37073_);
  or (_37078_, _37075_, _36911_);
  and (_37079_, _37078_, _06791_);
  and (_37080_, _37079_, _37076_);
  and (_37081_, _36911_, _06790_);
  or (_37082_, _37081_, _10865_);
  or (_37083_, _37082_, _37080_);
  nor (_37084_, _36924_, _14083_);
  nor (_37085_, _37084_, _36921_);
  and (_37086_, _37085_, _10891_);
  and (_37087_, _36921_, _10888_);
  or (_37089_, _37087_, _10867_);
  or (_37090_, _37089_, _37086_);
  and (_37091_, _37090_, _37083_);
  or (_37092_, _37091_, _06406_);
  nor (_37093_, _36993_, _14094_);
  nor (_37094_, _37093_, _36994_);
  and (_37095_, _37094_, _10921_);
  and (_37096_, _36994_, _10918_);
  or (_37097_, _37096_, _06407_);
  or (_37098_, _37097_, _37095_);
  and (_37100_, _37098_, _10927_);
  and (_37101_, _37100_, _37092_);
  or (_37102_, _37101_, _36898_);
  and (_37103_, _37102_, _10963_);
  nand (_37104_, _10997_, _36902_);
  nand (_37105_, _37104_, _18454_);
  nor (_37106_, _37105_, _14108_);
  or (_37107_, _37106_, _17195_);
  or (_37108_, _37107_, _37103_);
  and (_37109_, _36884_, _06276_);
  or (_37111_, _37109_, _11041_);
  and (_37112_, _37111_, _37108_);
  or (_37113_, _37112_, _36885_);
  and (_37114_, _37113_, _12690_);
  or (_37115_, _10297_, _08809_);
  and (_37116_, _14127_, _37115_);
  nand (_37117_, _11080_, _14131_);
  and (_37118_, _37117_, _14133_);
  or (_37119_, _37118_, _06433_);
  or (_37120_, _37119_, _37116_);
  or (_37122_, _37120_, _37114_);
  or (_37123_, _36949_, _06829_);
  and (_37124_, _37123_, _05749_);
  and (_37125_, _37124_, _37122_);
  and (_37126_, _36944_, _05748_);
  or (_37127_, _37126_, _06440_);
  or (_37128_, _37127_, _37125_);
  and (_37129_, _14710_, _07794_);
  or (_37130_, _36914_, _06444_);
  or (_37131_, _37130_, _37129_);
  and (_37133_, _37131_, _01317_);
  and (_37134_, _37133_, _37128_);
  or (_37135_, _37134_, _36881_);
  and (_43781_, _37135_, _43100_);
  and (_37136_, _01321_, \oc8051_golden_model_1.PSW [3]);
  and (_37137_, _14076_, \oc8051_golden_model_1.PSW [3]);
  and (_37138_, _07794_, _07544_);
  or (_37139_, _37138_, _37137_);
  or (_37140_, _37139_, _06132_);
  and (_37141_, _14738_, _07794_);
  or (_37143_, _37141_, _37137_);
  or (_37144_, _37143_, _06161_);
  and (_37145_, _07794_, \oc8051_golden_model_1.ACC [3]);
  or (_37146_, _37145_, _37137_);
  and (_37147_, _37146_, _07056_);
  and (_37148_, _07057_, \oc8051_golden_model_1.PSW [3]);
  or (_37149_, _37148_, _06160_);
  or (_37150_, _37149_, _37147_);
  and (_37151_, _37150_, _06157_);
  and (_37152_, _37151_, _37144_);
  and (_37154_, _36941_, \oc8051_golden_model_1.PSW [3]);
  and (_37155_, _14735_, _08404_);
  or (_37156_, _37155_, _37154_);
  and (_37157_, _37156_, _06156_);
  or (_37158_, _37157_, _06217_);
  or (_37159_, _37158_, _37152_);
  or (_37160_, _37139_, _07075_);
  and (_37161_, _37160_, _37159_);
  or (_37162_, _37161_, _06220_);
  or (_37163_, _37146_, _06229_);
  and (_37165_, _37163_, _06153_);
  and (_37166_, _37165_, _37162_);
  and (_37167_, _14731_, _08404_);
  or (_37168_, _37167_, _37154_);
  and (_37169_, _37168_, _06152_);
  or (_37170_, _37169_, _06145_);
  or (_37171_, _37170_, _37166_);
  or (_37172_, _37154_, _14764_);
  and (_37173_, _37172_, _37156_);
  or (_37174_, _37173_, _06146_);
  and (_37176_, _37174_, _06140_);
  and (_37177_, _37176_, _37171_);
  and (_37178_, _14732_, _08404_);
  or (_37179_, _37178_, _37154_);
  and (_37180_, _37179_, _06139_);
  or (_37181_, _37180_, _09842_);
  or (_37182_, _37181_, _37177_);
  and (_37183_, _37182_, _37140_);
  or (_37184_, _37183_, _06116_);
  and (_37185_, _09210_, _07794_);
  or (_37187_, _37137_, _06117_);
  or (_37188_, _37187_, _37185_);
  and (_37189_, _37188_, _06114_);
  and (_37190_, _37189_, _37184_);
  and (_37191_, _14825_, _07794_);
  or (_37192_, _37137_, _37191_);
  and (_37193_, _37192_, _05787_);
  or (_37194_, _37193_, _37190_);
  or (_37195_, _37194_, _11136_);
  and (_37196_, _14727_, _07794_);
  or (_37198_, _37137_, _07127_);
  or (_37199_, _37198_, _37196_);
  and (_37200_, _07794_, _08712_);
  or (_37201_, _37200_, _37137_);
  or (_37202_, _37201_, _06111_);
  and (_37203_, _37202_, _07125_);
  and (_37204_, _37203_, _37199_);
  and (_37205_, _37204_, _37195_);
  and (_37206_, _12318_, _07794_);
  or (_37207_, _37206_, _37137_);
  and (_37209_, _37207_, _06402_);
  or (_37210_, _37209_, _37205_);
  and (_37211_, _37210_, _07132_);
  or (_37212_, _37137_, _08140_);
  and (_37213_, _37201_, _06306_);
  and (_37214_, _37213_, _37212_);
  or (_37215_, _37214_, _37211_);
  and (_37216_, _37215_, _07130_);
  and (_37217_, _37146_, _06411_);
  and (_37218_, _37217_, _37212_);
  or (_37220_, _37218_, _06303_);
  or (_37221_, _37220_, _37216_);
  and (_37222_, _14724_, _07794_);
  or (_37223_, _37137_, _08819_);
  or (_37224_, _37223_, _37222_);
  and (_37225_, _37224_, _08824_);
  and (_37226_, _37225_, _37221_);
  nor (_37227_, _10273_, _14076_);
  or (_37228_, _37227_, _37137_);
  and (_37229_, _37228_, _06396_);
  or (_37231_, _37229_, _06433_);
  or (_37232_, _37231_, _37226_);
  or (_37233_, _37143_, _06829_);
  and (_37234_, _37233_, _05749_);
  and (_37235_, _37234_, _37232_);
  and (_37236_, _37168_, _05748_);
  or (_37237_, _37236_, _06440_);
  or (_37238_, _37237_, _37235_);
  and (_37239_, _14897_, _07794_);
  or (_37240_, _37137_, _06444_);
  or (_37242_, _37240_, _37239_);
  and (_37243_, _37242_, _01317_);
  and (_37244_, _37243_, _37238_);
  or (_37245_, _37244_, _37136_);
  and (_43783_, _37245_, _43100_);
  and (_37246_, _01321_, \oc8051_golden_model_1.PSW [4]);
  and (_37247_, _06284_, _05781_);
  and (_37248_, _14076_, \oc8051_golden_model_1.PSW [4]);
  and (_37249_, _08336_, _07794_);
  or (_37250_, _37249_, _37248_);
  or (_37252_, _37250_, _06132_);
  and (_37253_, _14928_, _07794_);
  or (_37254_, _37253_, _37248_);
  or (_37255_, _37254_, _06161_);
  and (_37256_, _07794_, \oc8051_golden_model_1.ACC [4]);
  or (_37257_, _37256_, _37248_);
  and (_37258_, _37257_, _07056_);
  and (_37259_, _07057_, \oc8051_golden_model_1.PSW [4]);
  or (_37260_, _37259_, _06160_);
  or (_37261_, _37260_, _37258_);
  and (_37263_, _37261_, _06157_);
  and (_37264_, _37263_, _37255_);
  and (_37265_, _36941_, \oc8051_golden_model_1.PSW [4]);
  and (_37266_, _14932_, _08404_);
  or (_37267_, _37266_, _37265_);
  and (_37268_, _37267_, _06156_);
  or (_37269_, _37268_, _06217_);
  or (_37270_, _37269_, _37264_);
  or (_37271_, _37250_, _07075_);
  and (_37272_, _37271_, _37270_);
  or (_37274_, _37272_, _06220_);
  or (_37275_, _37257_, _06229_);
  and (_37276_, _37275_, _06153_);
  and (_37277_, _37276_, _37274_);
  and (_37278_, _14942_, _08404_);
  or (_37279_, _37278_, _37265_);
  and (_37280_, _37279_, _06152_);
  or (_37281_, _37280_, _06145_);
  or (_37282_, _37281_, _37277_);
  or (_37283_, _37265_, _14949_);
  and (_37285_, _37283_, _37267_);
  or (_37286_, _37285_, _06146_);
  and (_37287_, _37286_, _06140_);
  and (_37288_, _37287_, _37282_);
  and (_37289_, _14966_, _08404_);
  or (_37290_, _37289_, _37265_);
  and (_37291_, _37290_, _06139_);
  or (_37292_, _37291_, _09842_);
  or (_37293_, _37292_, _37288_);
  and (_37294_, _37293_, _37252_);
  or (_37296_, _37294_, _37247_);
  and (_37297_, _09209_, _07794_);
  or (_37298_, _37297_, _37248_);
  and (_37299_, _37298_, _06276_);
  or (_37300_, _37299_, _06117_);
  and (_37301_, _37300_, _37296_);
  and (_37302_, _06281_, _05781_);
  and (_37303_, _37298_, _37302_);
  or (_37304_, _37303_, _05787_);
  or (_37305_, _37304_, _37301_);
  and (_37307_, _15013_, _07794_);
  or (_37308_, _37248_, _06114_);
  or (_37309_, _37308_, _37307_);
  and (_37310_, _37309_, _06111_);
  and (_37311_, _37310_, _37305_);
  and (_37312_, _08715_, _07794_);
  or (_37313_, _37312_, _37248_);
  and (_37314_, _37313_, _06110_);
  or (_37315_, _37314_, _06297_);
  or (_37316_, _37315_, _37311_);
  and (_37318_, _15029_, _07794_);
  or (_37319_, _37248_, _07127_);
  or (_37320_, _37319_, _37318_);
  and (_37321_, _37320_, _07125_);
  and (_37322_, _37321_, _37316_);
  and (_37323_, _10289_, _07794_);
  or (_37324_, _37323_, _37248_);
  and (_37325_, _37324_, _06402_);
  or (_37326_, _37325_, _37322_);
  and (_37327_, _37326_, _07132_);
  or (_37329_, _37248_, _08339_);
  and (_37330_, _37313_, _06306_);
  and (_37331_, _37330_, _37329_);
  or (_37332_, _37331_, _37327_);
  and (_37333_, _37332_, _07130_);
  and (_37334_, _37257_, _06411_);
  and (_37335_, _37334_, _37329_);
  or (_37336_, _37335_, _06303_);
  or (_37337_, _37336_, _37333_);
  and (_37338_, _15026_, _07794_);
  or (_37340_, _37248_, _08819_);
  or (_37341_, _37340_, _37338_);
  and (_37342_, _37341_, _08824_);
  and (_37343_, _37342_, _37337_);
  nor (_37344_, _10288_, _14076_);
  or (_37345_, _37344_, _37248_);
  and (_37346_, _37345_, _06396_);
  or (_37347_, _37346_, _06433_);
  or (_37348_, _37347_, _37343_);
  or (_37349_, _37254_, _06829_);
  and (_37351_, _37349_, _05749_);
  and (_37352_, _37351_, _37348_);
  and (_37353_, _37279_, _05748_);
  or (_37354_, _37353_, _06440_);
  or (_37355_, _37354_, _37352_);
  and (_37356_, _15087_, _07794_);
  or (_37357_, _37248_, _06444_);
  or (_37358_, _37357_, _37356_);
  and (_37359_, _37358_, _01317_);
  and (_37360_, _37359_, _37355_);
  or (_37362_, _37360_, _37246_);
  and (_43784_, _37362_, _43100_);
  and (_37363_, _01321_, \oc8051_golden_model_1.PSW [5]);
  and (_37364_, _14076_, \oc8051_golden_model_1.PSW [5]);
  and (_37365_, _15119_, _07794_);
  or (_37366_, _37365_, _37364_);
  or (_37367_, _37366_, _06161_);
  and (_37368_, _07794_, \oc8051_golden_model_1.ACC [5]);
  or (_37369_, _37368_, _37364_);
  and (_37370_, _37369_, _07056_);
  and (_37372_, _07057_, \oc8051_golden_model_1.PSW [5]);
  or (_37373_, _37372_, _06160_);
  or (_37374_, _37373_, _37370_);
  and (_37375_, _37374_, _06157_);
  and (_37376_, _37375_, _37367_);
  and (_37377_, _36941_, \oc8051_golden_model_1.PSW [5]);
  and (_37378_, _15123_, _08404_);
  or (_37379_, _37378_, _37377_);
  and (_37380_, _37379_, _06156_);
  or (_37381_, _37380_, _06217_);
  or (_37383_, _37381_, _37376_);
  and (_37384_, _08101_, _07794_);
  or (_37385_, _37384_, _37364_);
  or (_37386_, _37385_, _07075_);
  and (_37387_, _37386_, _37383_);
  or (_37388_, _37387_, _06220_);
  or (_37389_, _37369_, _06229_);
  and (_37390_, _37389_, _06153_);
  and (_37391_, _37390_, _37388_);
  and (_37392_, _15104_, _08404_);
  or (_37394_, _37392_, _37377_);
  and (_37395_, _37394_, _06152_);
  or (_37396_, _37395_, _06145_);
  or (_37397_, _37396_, _37391_);
  or (_37398_, _37377_, _15138_);
  and (_37399_, _37398_, _37379_);
  or (_37400_, _37399_, _06146_);
  and (_37401_, _37400_, _06140_);
  and (_37402_, _37401_, _37397_);
  and (_37403_, _15155_, _08404_);
  or (_37405_, _37403_, _37377_);
  and (_37406_, _37405_, _06139_);
  or (_37407_, _37406_, _09842_);
  or (_37408_, _37407_, _37402_);
  or (_37409_, _37385_, _06132_);
  and (_37410_, _37409_, _37408_);
  or (_37411_, _37410_, _06116_);
  and (_37412_, _09208_, _07794_);
  or (_37413_, _37364_, _06117_);
  or (_37414_, _37413_, _37412_);
  and (_37416_, _37414_, _06114_);
  and (_37417_, _37416_, _37411_);
  and (_37418_, _15203_, _07794_);
  or (_37419_, _37418_, _37364_);
  and (_37420_, _37419_, _05787_);
  or (_37421_, _37420_, _11136_);
  or (_37422_, _37421_, _37417_);
  and (_37423_, _15219_, _07794_);
  or (_37424_, _37364_, _07127_);
  or (_37425_, _37424_, _37423_);
  and (_37427_, _08736_, _07794_);
  or (_37428_, _37427_, _37364_);
  or (_37429_, _37428_, _06111_);
  and (_37430_, _37429_, _07125_);
  and (_37431_, _37430_, _37425_);
  and (_37432_, _37431_, _37422_);
  and (_37433_, _12325_, _07794_);
  or (_37434_, _37433_, _37364_);
  and (_37435_, _37434_, _06402_);
  or (_37436_, _37435_, _37432_);
  and (_37438_, _37436_, _07132_);
  or (_37439_, _37364_, _08104_);
  and (_37440_, _37428_, _06306_);
  and (_37441_, _37440_, _37439_);
  or (_37442_, _37441_, _37438_);
  and (_37443_, _37442_, _07130_);
  and (_37444_, _37369_, _06411_);
  and (_37445_, _37444_, _37439_);
  or (_37446_, _37445_, _06303_);
  or (_37447_, _37446_, _37443_);
  and (_37449_, _15216_, _07794_);
  or (_37450_, _37364_, _08819_);
  or (_37451_, _37450_, _37449_);
  and (_37452_, _37451_, _08824_);
  and (_37453_, _37452_, _37447_);
  nor (_37454_, _10269_, _14076_);
  or (_37455_, _37454_, _37364_);
  and (_37456_, _37455_, _06396_);
  or (_37457_, _37456_, _06433_);
  or (_37458_, _37457_, _37453_);
  or (_37460_, _37366_, _06829_);
  and (_37461_, _37460_, _05749_);
  and (_37462_, _37461_, _37458_);
  and (_37463_, _37394_, _05748_);
  or (_37464_, _37463_, _06440_);
  or (_37465_, _37464_, _37462_);
  and (_37466_, _15275_, _07794_);
  or (_37467_, _37364_, _06444_);
  or (_37468_, _37467_, _37466_);
  and (_37469_, _37468_, _01317_);
  and (_37471_, _37469_, _37465_);
  or (_37472_, _37471_, _37363_);
  and (_43785_, _37472_, _43100_);
  nor (_37473_, _01317_, _17884_);
  or (_37474_, _10942_, _10654_);
  and (_37475_, _37474_, _10895_);
  nor (_37476_, _10882_, _10601_);
  nand (_37477_, _37476_, _17240_);
  not (_37478_, _10372_);
  or (_37479_, _10361_, _10324_);
  and (_37481_, _37479_, _37478_);
  and (_37482_, _15410_, _07794_);
  nor (_37483_, _07794_, _17884_);
  or (_37484_, _37483_, _08819_);
  or (_37485_, _37484_, _37482_);
  and (_37486_, _08012_, _07794_);
  or (_37487_, _37486_, _37483_);
  or (_37488_, _37487_, _06132_);
  or (_37489_, _10634_, _10601_);
  or (_37490_, _37489_, _12380_);
  nor (_37492_, _08404_, _17884_);
  and (_37493_, _15297_, _08404_);
  or (_37494_, _37493_, _37492_);
  and (_37495_, _37494_, _06152_);
  and (_37496_, _15300_, _07794_);
  or (_37497_, _37496_, _37483_);
  or (_37498_, _37497_, _06161_);
  and (_37499_, _07794_, \oc8051_golden_model_1.ACC [6]);
  or (_37500_, _37499_, _37483_);
  and (_37501_, _37500_, _07056_);
  nor (_37503_, _07056_, _17884_);
  or (_37504_, _37503_, _06160_);
  or (_37505_, _37504_, _37501_);
  and (_37506_, _37505_, _06157_);
  and (_37507_, _37506_, _37498_);
  and (_37508_, _15316_, _08404_);
  or (_37509_, _37508_, _37492_);
  and (_37510_, _37509_, _06156_);
  or (_37511_, _37510_, _06217_);
  or (_37512_, _37511_, _37507_);
  or (_37514_, _37487_, _07075_);
  and (_37515_, _37514_, _37512_);
  or (_37516_, _37515_, _06220_);
  or (_37517_, _37500_, _06229_);
  and (_37518_, _37517_, _06153_);
  and (_37519_, _37518_, _37516_);
  or (_37520_, _37519_, _37495_);
  and (_37521_, _37520_, _06146_);
  or (_37522_, _37492_, _15331_);
  and (_37523_, _37522_, _06145_);
  and (_37525_, _37523_, _37509_);
  or (_37526_, _37525_, _10557_);
  or (_37527_, _37526_, _37521_);
  or (_37528_, _10554_, _10324_);
  or (_37529_, _37528_, _10568_);
  and (_37530_, _37529_, _37527_);
  or (_37531_, _37530_, _12379_);
  and (_37532_, _37531_, _37490_);
  and (_37533_, _37532_, _06265_);
  or (_37534_, _10441_, _10392_);
  and (_37536_, _37534_, _06260_);
  or (_37537_, _37536_, _10387_);
  or (_37538_, _37537_, _37533_);
  or (_37539_, _10654_, _10388_);
  or (_37540_, _37539_, _10708_);
  and (_37541_, _37540_, _06140_);
  and (_37542_, _37541_, _37538_);
  and (_37543_, _15348_, _08404_);
  or (_37544_, _37543_, _37492_);
  and (_37545_, _37544_, _06139_);
  or (_37547_, _37545_, _09842_);
  or (_37548_, _37547_, _37542_);
  and (_37549_, _37548_, _37488_);
  or (_37550_, _37549_, _06116_);
  and (_37551_, _09207_, _07794_);
  or (_37552_, _37483_, _06117_);
  or (_37553_, _37552_, _37551_);
  and (_37554_, _37553_, _06114_);
  and (_37555_, _37554_, _37550_);
  and (_37556_, _15395_, _07794_);
  or (_37558_, _37556_, _37483_);
  and (_37559_, _37558_, _05787_);
  or (_37560_, _37559_, _11136_);
  or (_37561_, _37560_, _37555_);
  and (_37562_, _15413_, _07794_);
  or (_37563_, _37483_, _07127_);
  or (_37564_, _37563_, _37562_);
  and (_37565_, _15402_, _07794_);
  or (_37566_, _37565_, _37483_);
  or (_37567_, _37566_, _06111_);
  and (_37569_, _37567_, _07125_);
  and (_37570_, _37569_, _37564_);
  and (_37571_, _37570_, _37561_);
  and (_37572_, _10295_, _07794_);
  or (_37573_, _37572_, _37483_);
  and (_37574_, _37573_, _06402_);
  or (_37575_, _37574_, _37571_);
  and (_37576_, _37575_, _07132_);
  or (_37577_, _37483_, _08015_);
  and (_37578_, _37566_, _06306_);
  and (_37580_, _37578_, _37577_);
  or (_37581_, _37580_, _37576_);
  and (_37582_, _37581_, _07130_);
  and (_37583_, _37500_, _06411_);
  and (_37584_, _37583_, _37577_);
  or (_37585_, _37584_, _06303_);
  or (_37586_, _37585_, _37582_);
  and (_37587_, _37586_, _37485_);
  or (_37588_, _37587_, _06396_);
  nor (_37589_, _10294_, _14076_);
  or (_37591_, _37589_, _37483_);
  or (_37592_, _37591_, _08824_);
  and (_37593_, _37592_, _10372_);
  and (_37594_, _37593_, _37588_);
  or (_37595_, _37594_, _37481_);
  and (_37596_, _37595_, _10375_);
  and (_37597_, _37479_, _06794_);
  nor (_37598_, _37597_, _37596_);
  nor (_37599_, _37598_, _10376_);
  and (_37600_, _37479_, _10376_);
  or (_37602_, _37600_, _06795_);
  or (_37603_, _37602_, _37599_);
  not (_37604_, _06795_);
  or (_37605_, _37479_, _37604_);
  and (_37606_, _37605_, _10374_);
  and (_37607_, _37606_, _37603_);
  and (_37608_, _37479_, _10373_);
  or (_37609_, _37608_, _37607_);
  or (_37610_, _37609_, _17240_);
  and (_37611_, _37610_, _37477_);
  or (_37613_, _37611_, _06792_);
  nand (_37614_, _37476_, _06792_);
  and (_37615_, _37614_, _37613_);
  or (_37616_, _37615_, _06406_);
  nor (_37617_, _10901_, _10392_);
  nand (_37618_, _37617_, _18090_);
  and (_37619_, _37618_, _10927_);
  and (_37620_, _37619_, _37616_);
  or (_37621_, _37620_, _37475_);
  and (_37622_, _37621_, _10963_);
  and (_37624_, _10991_, _18454_);
  or (_37625_, _37624_, _11003_);
  or (_37626_, _37625_, _37622_);
  or (_37627_, _11033_, _11041_);
  and (_37628_, _37627_, _06171_);
  and (_37629_, _37628_, _37626_);
  and (_37630_, _10287_, _06169_);
  or (_37631_, _37630_, _10264_);
  or (_37632_, _37631_, _37629_);
  or (_37633_, _11074_, _10265_);
  and (_37635_, _37633_, _37632_);
  or (_37636_, _37635_, _06433_);
  or (_37637_, _37497_, _06829_);
  and (_37638_, _37637_, _05749_);
  and (_37639_, _37638_, _37636_);
  and (_37640_, _37494_, _05748_);
  or (_37641_, _37640_, _06440_);
  or (_37642_, _37641_, _37639_);
  and (_37643_, _15478_, _07794_);
  or (_37644_, _37483_, _06444_);
  or (_37646_, _37644_, _37643_);
  and (_37647_, _37646_, _01317_);
  and (_37648_, _37647_, _37642_);
  or (_37649_, _37648_, _37473_);
  and (_43786_, _37649_, _43100_);
  and (_37650_, _05820_, op0_cnst);
  or (_00001_, _37650_, rst);
  and (_37651_, inst_finished_r, op0_cnst);
  not (_37652_, word_in[1]);
  and (_37653_, _37652_, word_in[0]);
  and (_37655_, _37653_, \oc8051_golden_model_1.IRAM[1] [3]);
  nor (_37656_, _37652_, word_in[0]);
  and (_37657_, _37656_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor (_37658_, _37657_, _37655_);
  nor (_37659_, word_in[1], word_in[0]);
  and (_37660_, _37659_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_37661_, word_in[1], word_in[0]);
  and (_37662_, _37661_, \oc8051_golden_model_1.IRAM[3] [3]);
  nor (_37663_, _37662_, _37660_);
  and (_37664_, _37663_, _37658_);
  nor (_37666_, word_in[3], word_in[2]);
  not (_37667_, _37666_);
  nor (_37668_, _37667_, _37664_);
  and (_37669_, _37653_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_37670_, _37656_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor (_37671_, _37670_, _37669_);
  and (_37672_, _37659_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_37673_, _37661_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor (_37674_, _37673_, _37672_);
  and (_37675_, _37674_, _37671_);
  and (_37677_, word_in[3], word_in[2]);
  not (_37678_, _37677_);
  nor (_37679_, _37678_, _37675_);
  nor (_37680_, _37679_, _37668_);
  and (_37681_, _37653_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_37682_, _37656_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor (_37683_, _37682_, _37681_);
  and (_37684_, _37659_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_37685_, _37661_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor (_37686_, _37685_, _37684_);
  and (_37688_, _37686_, _37683_);
  not (_37689_, word_in[3]);
  and (_37690_, _37689_, word_in[2]);
  not (_37691_, _37690_);
  nor (_37692_, _37691_, _37688_);
  and (_37693_, _37653_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_37694_, _37656_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor (_37695_, _37694_, _37693_);
  and (_37696_, _37659_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_37697_, _37661_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor (_37699_, _37697_, _37696_);
  and (_37700_, _37699_, _37695_);
  nor (_37701_, _37689_, word_in[2]);
  not (_37702_, _37701_);
  nor (_37703_, _37702_, _37700_);
  nor (_37704_, _37703_, _37692_);
  and (_37705_, _37704_, _37680_);
  and (_37706_, _37690_, _37661_);
  and (_37707_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_37708_, _37666_, _37661_);
  and (_37710_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_37711_, _37710_, _37707_);
  and (_37712_, _37677_, _37656_);
  and (_37713_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_37714_, _37677_, _37659_);
  and (_37715_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_37716_, _37715_, _37713_);
  and (_37717_, _37716_, _37711_);
  and (_37718_, _37666_, _37656_);
  and (_37719_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_37721_, _37666_, _37653_);
  and (_37722_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_37723_, _37722_, _37719_);
  and (_37724_, _37690_, _37653_);
  and (_37725_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_37726_, _37690_, _37659_);
  and (_37727_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_37728_, _37727_, _37725_);
  and (_37729_, _37728_, _37723_);
  and (_37730_, _37729_, _37717_);
  and (_37732_, _37701_, _37656_);
  and (_37733_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_37734_, _37701_, _37659_);
  and (_37735_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_37736_, _37735_, _37733_);
  and (_37737_, _37677_, _37661_);
  and (_37738_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_37739_, _37677_, _37653_);
  and (_37740_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_37741_, _37740_, _37738_);
  and (_37743_, _37741_, _37736_);
  and (_37744_, _37690_, _37656_);
  and (_37745_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_37746_, _37666_, _37659_);
  and (_37747_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_37748_, _37747_, _37745_);
  and (_37749_, _37701_, _37661_);
  and (_37750_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_37751_, _37701_, _37653_);
  and (_37752_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_37754_, _37752_, _37750_);
  and (_37755_, _37754_, _37748_);
  and (_37756_, _37755_, _37743_);
  and (_37757_, _37756_, _37730_);
  nand (_37758_, _37757_, _37705_);
  or (_37759_, _37757_, _37705_);
  and (_37760_, _37759_, _37758_);
  and (_37761_, _37653_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_37762_, _37656_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor (_37763_, _37762_, _37761_);
  and (_37765_, _37659_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_37766_, _37661_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor (_37767_, _37766_, _37765_);
  and (_37768_, _37767_, _37763_);
  nor (_37769_, _37768_, _37667_);
  and (_37770_, _37653_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_37771_, _37656_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor (_37772_, _37771_, _37770_);
  and (_37773_, _37659_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_37774_, _37661_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor (_37776_, _37774_, _37773_);
  and (_37777_, _37776_, _37772_);
  nor (_37778_, _37777_, _37678_);
  nor (_37779_, _37778_, _37769_);
  and (_37780_, _37653_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_37781_, _37656_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor (_37782_, _37781_, _37780_);
  and (_37783_, _37659_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_37784_, _37661_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor (_37785_, _37784_, _37783_);
  and (_37787_, _37785_, _37782_);
  nor (_37788_, _37787_, _37691_);
  and (_37789_, _37653_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_37790_, _37656_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor (_37791_, _37790_, _37789_);
  and (_37792_, _37659_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_37793_, _37661_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor (_37794_, _37793_, _37792_);
  and (_37795_, _37794_, _37791_);
  nor (_37796_, _37795_, _37702_);
  nor (_37798_, _37796_, _37788_);
  and (_37799_, _37798_, _37779_);
  and (_37800_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_37801_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_37802_, _37801_, _37800_);
  and (_37803_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_37804_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_37805_, _37804_, _37803_);
  and (_37806_, _37805_, _37802_);
  and (_37807_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_37809_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_37810_, _37809_, _37807_);
  and (_37811_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_37812_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_37813_, _37812_, _37811_);
  and (_37814_, _37813_, _37810_);
  and (_37815_, _37814_, _37806_);
  and (_37816_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_37817_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_37818_, _37817_, _37816_);
  and (_37820_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_37821_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_37822_, _37821_, _37820_);
  and (_37823_, _37822_, _37818_);
  and (_37824_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_37825_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_37826_, _37825_, _37824_);
  and (_37827_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_37828_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_37829_, _37828_, _37827_);
  and (_37831_, _37829_, _37826_);
  and (_37832_, _37831_, _37823_);
  and (_37833_, _37832_, _37815_);
  nand (_37834_, _37833_, _37799_);
  or (_37835_, _37833_, _37799_);
  and (_37836_, _37835_, _37834_);
  or (_37837_, _37836_, _37760_);
  and (_37838_, _37653_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_37839_, _37656_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor (_37840_, _37839_, _37838_);
  and (_37842_, _37659_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_37843_, _37661_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor (_37844_, _37843_, _37842_);
  and (_37845_, _37844_, _37840_);
  nor (_37846_, _37845_, _37691_);
  and (_37847_, _37653_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_37848_, _37656_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor (_37849_, _37848_, _37847_);
  and (_37850_, _37659_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_37851_, _37661_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor (_37853_, _37851_, _37850_);
  and (_37854_, _37853_, _37849_);
  nor (_37855_, _37854_, _37678_);
  nor (_37856_, _37855_, _37846_);
  and (_37857_, _37653_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_37858_, _37656_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor (_37859_, _37858_, _37857_);
  and (_37860_, _37659_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_37861_, _37661_, \oc8051_golden_model_1.IRAM[3] [1]);
  nor (_37862_, _37861_, _37860_);
  and (_37864_, _37862_, _37859_);
  nor (_37865_, _37864_, _37667_);
  and (_37866_, _37653_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_37867_, _37656_, \oc8051_golden_model_1.IRAM[10] [1]);
  nor (_37868_, _37867_, _37866_);
  and (_37869_, _37659_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_37870_, _37661_, \oc8051_golden_model_1.IRAM[11] [1]);
  nor (_37871_, _37870_, _37869_);
  and (_37872_, _37871_, _37868_);
  nor (_37873_, _37872_, _37702_);
  nor (_37875_, _37873_, _37865_);
  and (_37876_, _37875_, _37856_);
  and (_37877_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_37878_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_37879_, _37878_, _37877_);
  and (_37880_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_37881_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_37882_, _37881_, _37880_);
  and (_37883_, _37882_, _37879_);
  and (_37884_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_37886_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_37887_, _37886_, _37884_);
  and (_37888_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_37889_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_37890_, _37889_, _37888_);
  and (_37891_, _37890_, _37887_);
  and (_37892_, _37891_, _37883_);
  and (_37893_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_37894_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_37895_, _37894_, _37893_);
  and (_37897_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_37898_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_37899_, _37898_, _37897_);
  and (_37900_, _37899_, _37895_);
  and (_37901_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_37902_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_37903_, _37902_, _37901_);
  and (_37904_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_37905_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_37906_, _37905_, _37904_);
  and (_37908_, _37906_, _37903_);
  and (_37909_, _37908_, _37900_);
  and (_37910_, _37909_, _37892_);
  nand (_37911_, _37910_, _37876_);
  or (_37912_, _37910_, _37876_);
  and (_37913_, _37912_, _37911_);
  and (_37914_, _37653_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_37915_, _37656_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor (_37916_, _37915_, _37914_);
  and (_37917_, _37659_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_37919_, _37661_, \oc8051_golden_model_1.IRAM[3] [0]);
  nor (_37920_, _37919_, _37917_);
  and (_37921_, _37920_, _37916_);
  nor (_37922_, _37921_, _37667_);
  and (_37923_, _37653_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_37924_, _37656_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor (_37925_, _37924_, _37923_);
  and (_37926_, _37659_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_37927_, _37661_, \oc8051_golden_model_1.IRAM[11] [0]);
  nor (_37928_, _37927_, _37926_);
  and (_37930_, _37928_, _37925_);
  nor (_37931_, _37930_, _37702_);
  nor (_37932_, _37931_, _37922_);
  and (_37933_, _37653_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_37934_, _37656_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor (_37935_, _37934_, _37933_);
  and (_37936_, _37659_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_37937_, _37661_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor (_37938_, _37937_, _37936_);
  and (_37939_, _37938_, _37935_);
  nor (_37941_, _37939_, _37691_);
  and (_37942_, _37653_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_37943_, _37656_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor (_37944_, _37943_, _37942_);
  and (_37945_, _37659_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_37946_, _37661_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor (_37947_, _37946_, _37945_);
  and (_37948_, _37947_, _37944_);
  nor (_37949_, _37948_, _37678_);
  nor (_37950_, _37949_, _37941_);
  and (_37952_, _37950_, _37932_);
  and (_37953_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_37954_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_37955_, _37954_, _37953_);
  and (_37956_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_37957_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_37958_, _37957_, _37956_);
  and (_37959_, _37958_, _37955_);
  and (_37960_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_37961_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_37963_, _37961_, _37960_);
  and (_37964_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_37965_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_37966_, _37965_, _37964_);
  and (_37967_, _37966_, _37963_);
  and (_37968_, _37967_, _37959_);
  and (_37969_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_37970_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_37971_, _37970_, _37969_);
  and (_37972_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_37974_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_37975_, _37974_, _37972_);
  and (_37976_, _37975_, _37971_);
  and (_37977_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_37978_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_37979_, _37978_, _37977_);
  and (_37980_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_37981_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_37982_, _37981_, _37980_);
  and (_37983_, _37982_, _37979_);
  and (_37985_, _37983_, _37976_);
  and (_37986_, _37985_, _37968_);
  nand (_37987_, _37986_, _37952_);
  or (_37988_, _37986_, _37952_);
  and (_37989_, _37988_, _37987_);
  or (_37990_, _37989_, _37913_);
  or (_37991_, _37990_, _37837_);
  and (_37992_, _37653_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_37993_, _37656_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor (_37994_, _37993_, _37992_);
  and (_37996_, _37659_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_37997_, _37661_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor (_37998_, _37997_, _37996_);
  and (_37999_, _37998_, _37994_);
  nor (_38000_, _37999_, _37691_);
  and (_38001_, _37653_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_38002_, _37656_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor (_38003_, _38002_, _38001_);
  and (_38004_, _37659_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_38005_, _37661_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor (_38007_, _38005_, _38004_);
  and (_38008_, _38007_, _38003_);
  nor (_38009_, _38008_, _37678_);
  nor (_38010_, _38009_, _38000_);
  and (_38011_, _37653_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_38012_, _37656_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor (_38013_, _38012_, _38011_);
  and (_38014_, _37659_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_38015_, _37661_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor (_38016_, _38015_, _38014_);
  and (_38018_, _38016_, _38013_);
  nor (_38019_, _38018_, _37667_);
  and (_38020_, _37653_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_38021_, _37656_, \oc8051_golden_model_1.IRAM[10] [4]);
  nor (_38022_, _38021_, _38020_);
  and (_38023_, _37659_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_38024_, _37661_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor (_38025_, _38024_, _38023_);
  and (_38026_, _38025_, _38022_);
  nor (_38027_, _38026_, _37702_);
  nor (_38029_, _38027_, _38019_);
  and (_38030_, _38029_, _38010_);
  and (_38031_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_38032_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_38033_, _38032_, _38031_);
  and (_38034_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_38035_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_38036_, _38035_, _38034_);
  and (_38037_, _38036_, _38033_);
  and (_38038_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_38040_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_38041_, _38040_, _38038_);
  and (_38042_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_38043_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_38044_, _38043_, _38042_);
  and (_38045_, _38044_, _38041_);
  and (_38046_, _38045_, _38037_);
  and (_38047_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_38048_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_38049_, _38048_, _38047_);
  and (_38051_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_38052_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_38053_, _38052_, _38051_);
  and (_38054_, _38053_, _38049_);
  and (_38055_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_38056_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_38057_, _38056_, _38055_);
  and (_38058_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_38059_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_38060_, _38059_, _38058_);
  and (_38062_, _38060_, _38057_);
  and (_38063_, _38062_, _38054_);
  and (_38064_, _38063_, _38046_);
  nand (_38065_, _38064_, _38030_);
  or (_38066_, _38064_, _38030_);
  and (_38067_, _38066_, _38065_);
  and (_38068_, _37653_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_38069_, _37656_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor (_38070_, _38069_, _38068_);
  and (_38071_, _37659_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_38073_, _37661_, \oc8051_golden_model_1.IRAM[3] [5]);
  nor (_38074_, _38073_, _38071_);
  and (_38075_, _38074_, _38070_);
  nor (_38076_, _38075_, _37667_);
  and (_38077_, _37653_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_38078_, _37656_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor (_38079_, _38078_, _38077_);
  and (_38080_, _37659_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_38081_, _37661_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor (_38082_, _38081_, _38080_);
  and (_38084_, _38082_, _38079_);
  nor (_38085_, _38084_, _37678_);
  nor (_38086_, _38085_, _38076_);
  and (_38087_, _37653_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_38088_, _37656_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor (_38089_, _38088_, _38087_);
  and (_38090_, _37659_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_38091_, _37661_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor (_38092_, _38091_, _38090_);
  and (_38093_, _38092_, _38089_);
  nor (_38095_, _38093_, _37691_);
  and (_38096_, _37653_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_38097_, _37656_, \oc8051_golden_model_1.IRAM[10] [5]);
  nor (_38098_, _38097_, _38096_);
  and (_38099_, _37659_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_38100_, _37661_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor (_38101_, _38100_, _38099_);
  and (_38102_, _38101_, _38098_);
  nor (_38103_, _38102_, _37702_);
  nor (_38104_, _38103_, _38095_);
  and (_38106_, _38104_, _38086_);
  and (_38107_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_38108_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_38109_, _38108_, _38107_);
  and (_38110_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_38111_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_38112_, _38111_, _38110_);
  and (_38113_, _38112_, _38109_);
  and (_38114_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_38115_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_38117_, _38115_, _38114_);
  and (_38118_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_38119_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_38120_, _38119_, _38118_);
  and (_38121_, _38120_, _38117_);
  and (_38122_, _38121_, _38113_);
  and (_38123_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_38124_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_38125_, _38124_, _38123_);
  and (_38126_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_38128_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_38129_, _38128_, _38126_);
  and (_38130_, _38129_, _38125_);
  and (_38131_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_38132_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_38133_, _38132_, _38131_);
  and (_38134_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_38135_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_38136_, _38135_, _38134_);
  and (_38137_, _38136_, _38133_);
  and (_38139_, _38137_, _38130_);
  and (_38140_, _38139_, _38122_);
  nand (_38141_, _38140_, _38106_);
  or (_38142_, _38140_, _38106_);
  and (_38143_, _38142_, _38141_);
  or (_38144_, _38143_, _38067_);
  and (_38145_, _37653_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_38146_, _37656_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor (_38147_, _38146_, _38145_);
  and (_38148_, _37659_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_38150_, _37661_, \oc8051_golden_model_1.IRAM[7] [7]);
  nor (_38151_, _38150_, _38148_);
  and (_38152_, _38151_, _38147_);
  nor (_38153_, _38152_, _37691_);
  and (_38154_, _37653_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_38155_, _37656_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_38156_, _38155_, _38154_);
  and (_38157_, _37659_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_38158_, _37661_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor (_38159_, _38158_, _38157_);
  and (_38161_, _38159_, _38156_);
  nor (_38162_, _38161_, _37678_);
  nor (_38163_, _38162_, _38153_);
  and (_38164_, _37653_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_38165_, _37656_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor (_38166_, _38165_, _38164_);
  and (_38167_, _37659_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_38168_, _37661_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor (_38169_, _38168_, _38167_);
  and (_38170_, _38169_, _38166_);
  nor (_38172_, _38170_, _37667_);
  and (_38173_, _37653_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_38174_, _37656_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor (_38175_, _38174_, _38173_);
  and (_38176_, _37659_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_38177_, _37661_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor (_38178_, _38177_, _38176_);
  and (_38179_, _38178_, _38175_);
  nor (_38180_, _38179_, _37702_);
  nor (_38181_, _38180_, _38172_);
  and (_38183_, _38181_, _38163_);
  and (_38184_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_38185_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_38186_, _38185_, _38184_);
  and (_38187_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_38188_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_38189_, _38188_, _38187_);
  and (_38190_, _38189_, _38186_);
  and (_38191_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_38192_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_38194_, _38192_, _38191_);
  and (_38195_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_38196_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_38197_, _38196_, _38195_);
  and (_38198_, _38197_, _38194_);
  and (_38199_, _38198_, _38190_);
  and (_38200_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_38201_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor (_38202_, _38201_, _38200_);
  and (_38203_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_38205_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_38206_, _38205_, _38203_);
  and (_38207_, _38206_, _38202_);
  and (_38208_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_38209_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_38210_, _38209_, _38208_);
  and (_38211_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_38212_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_38213_, _38212_, _38211_);
  and (_38214_, _38213_, _38210_);
  and (_38216_, _38214_, _38207_);
  and (_38217_, _38216_, _38199_);
  nand (_38218_, _38217_, _38183_);
  or (_38219_, _38217_, _38183_);
  and (_38220_, _38219_, _38218_);
  and (_38221_, _37653_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_38222_, _37656_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor (_38223_, _38222_, _38221_);
  and (_38224_, _37659_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_38225_, _37661_, \oc8051_golden_model_1.IRAM[3] [6]);
  nor (_38227_, _38225_, _38224_);
  and (_38228_, _38227_, _38223_);
  nor (_38229_, _38228_, _37667_);
  and (_38230_, _37653_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_38231_, _37656_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor (_38232_, _38231_, _38230_);
  and (_38233_, _37659_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_38234_, _37661_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor (_38235_, _38234_, _38233_);
  and (_38236_, _38235_, _38232_);
  nor (_38238_, _38236_, _37702_);
  nor (_38239_, _38238_, _38229_);
  and (_38240_, _37653_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_38241_, _37656_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor (_38242_, _38241_, _38240_);
  and (_38243_, _37659_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_38244_, _37661_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor (_38245_, _38244_, _38243_);
  and (_38246_, _38245_, _38242_);
  nor (_38247_, _38246_, _37691_);
  and (_38249_, _37653_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_38250_, _37656_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor (_38251_, _38250_, _38249_);
  and (_38252_, _37659_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_38253_, _37661_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor (_38254_, _38253_, _38252_);
  and (_38255_, _38254_, _38251_);
  nor (_38256_, _38255_, _37678_);
  nor (_38257_, _38256_, _38247_);
  and (_38258_, _38257_, _38239_);
  and (_38260_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_38261_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_38262_, _38261_, _38260_);
  and (_38263_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_38264_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_38265_, _38264_, _38263_);
  and (_38266_, _38265_, _38262_);
  and (_38267_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_38268_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_38269_, _38268_, _38267_);
  and (_38271_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_38272_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_38273_, _38272_, _38271_);
  and (_38274_, _38273_, _38269_);
  and (_38275_, _38274_, _38266_);
  and (_38276_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_38277_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_38278_, _38277_, _38276_);
  and (_38279_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_38280_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_38282_, _38280_, _38279_);
  and (_38283_, _38282_, _38278_);
  and (_38284_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_38285_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_38286_, _38285_, _38284_);
  and (_38287_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_38288_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_38289_, _38288_, _38287_);
  and (_38290_, _38289_, _38286_);
  and (_38291_, _38290_, _38283_);
  and (_38293_, _38291_, _38275_);
  not (_38294_, _38293_);
  nor (_38295_, _38294_, _38258_);
  and (_38296_, _38294_, _38258_);
  or (_38297_, _38296_, _38295_);
  or (_38298_, _38297_, _38220_);
  or (_38299_, _38298_, _38144_);
  or (_38300_, _38299_, _37991_);
  and (property_invalid_iram, _38300_, _37651_);
  nor (_38301_, _09981_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_38303_, _09981_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_38304_, _38303_, _38301_);
  nand (_38305_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_38306_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38307_, _38306_, _38305_);
  or (_38308_, _38307_, _38304_);
  and (_38309_, _05887_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_38310_, _05887_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_38311_, _38310_, _38309_);
  and (_38312_, _05855_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_38314_, \oc8051_golden_model_1.ACC [0], _39264_);
  or (_38315_, _38314_, _38312_);
  or (_38316_, _38315_, _38311_);
  or (_38317_, _38316_, _38308_);
  or (_38318_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_38319_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_38320_, _38319_, _38318_);
  or (_38321_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_38322_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38323_, _38322_, _38321_);
  or (_38325_, _38323_, _38320_);
  nand (_38326_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_38327_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_38328_, _38327_, _38326_);
  and (_38329_, _08430_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_38330_, _08430_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_38331_, _38330_, _38329_);
  or (_38332_, _38331_, _38328_);
  or (_38333_, _38332_, _38325_);
  or (_38334_, _38333_, _38317_);
  and (property_invalid_acc, _38334_, _37651_);
  nor (_38336_, _25393_, _01950_);
  and (_38337_, _26427_, _01962_);
  and (_38338_, _25393_, _01950_);
  or (_38339_, _38338_, _38337_);
  or (_38340_, _38339_, _38336_);
  nor (_38341_, _27478_, _01973_);
  and (_38342_, _27478_, _01973_);
  nor (_38343_, _26780_, _01966_);
  or (_38344_, _38343_, _38342_);
  or (_38346_, _38344_, _38341_);
  nor (_38347_, _26427_, _01962_);
  and (_38348_, _26780_, _01966_);
  nand (_38349_, _27123_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_38350_, _27123_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_38351_, _38350_, _38349_);
  nor (_38352_, _26084_, _01958_);
  and (_38353_, _26084_, _01958_);
  nor (_38354_, _28124_, _38782_);
  and (_38355_, _28124_, _38782_);
  nor (_38357_, _12760_, _38760_);
  nor (_38358_, _28439_, _38787_);
  and (_38359_, _12760_, _38760_);
  or (_38360_, _38359_, _38358_);
  or (_38361_, _38360_, _38357_);
  and (_38362_, _28742_, _38772_);
  nor (_38363_, _28742_, _38772_);
  or (_38364_, _38363_, _38362_);
  and (_38365_, _29365_, _38768_);
  and (_38366_, _28439_, _38787_);
  or (_38368_, _38366_, _38365_);
  or (_38369_, _38368_, _38364_);
  nand (_38370_, _27800_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_38371_, _27800_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38372_, _38371_, _38370_);
  nor (_38373_, _29365_, _38768_);
  nor (_38374_, _29666_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38375_, _29666_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38376_, _25025_, _01946_);
  nor (_38377_, _25025_, _01946_);
  or (_38379_, _38377_, _38376_);
  or (_38380_, _38379_, _38375_);
  or (_38381_, _38380_, _38374_);
  nor (_38382_, _29057_, _38793_);
  and (_38383_, _29057_, _38793_);
  or (_38384_, _38383_, _38382_);
  or (_38385_, _38384_, _38381_);
  or (_38386_, _38385_, _38373_);
  or (_38387_, _38386_, _38372_);
  or (_38388_, _38387_, _38369_);
  or (_38390_, _38388_, _38361_);
  or (_38391_, _38390_, _38355_);
  or (_38392_, _38391_, _38354_);
  or (_38393_, _38392_, _38353_);
  or (_38394_, _38393_, _38352_);
  or (_38395_, _38394_, _38351_);
  or (_38396_, _38395_, _38348_);
  or (_38397_, _38396_, _38347_);
  or (_38398_, _38397_, _38346_);
  or (_38399_, _38398_, _38340_);
  and (_38401_, _25749_, _01954_);
  nor (_38402_, _25749_, _01954_);
  or (_38403_, _38402_, _38401_);
  or (_38404_, _38403_, _38399_);
  and (_38405_, _37650_, _01317_);
  and (property_invalid_pc, _38405_, _38404_);
  buf (_00544_, _43102_);
  buf (_05108_, _43100_);
  buf (_05159_, _43100_);
  buf (_05211_, _43100_);
  buf (_05262_, _43100_);
  buf (_05314_, _43100_);
  buf (_05365_, _43100_);
  buf (_05417_, _43100_);
  buf (_05470_, _43100_);
  buf (_05523_, _43100_);
  buf (_05576_, _43100_);
  buf (_05629_, _43100_);
  buf (_05682_, _43100_);
  buf (_05735_, _43100_);
  buf (_05788_, _43100_);
  buf (_05841_, _43100_);
  buf (_05894_, _43100_);
  buf (_39277_, _39174_);
  buf (_39279_, _39176_);
  buf (_39292_, _39174_);
  buf (_39293_, _39176_);
  buf (_39605_, _39194_);
  buf (_39606_, _39195_);
  buf (_39607_, _39197_);
  buf (_39608_, _39198_);
  buf (_39609_, _39199_);
  buf (_39610_, _39200_);
  buf (_39611_, _39201_);
  buf (_39612_, _39203_);
  buf (_39613_, _39204_);
  buf (_39615_, _39205_);
  buf (_39616_, _39206_);
  buf (_39617_, _39207_);
  buf (_39618_, _39209_);
  buf (_39619_, _39210_);
  buf (_39670_, _39194_);
  buf (_39671_, _39195_);
  buf (_39672_, _39197_);
  buf (_39673_, _39198_);
  buf (_39674_, _39199_);
  buf (_39675_, _39200_);
  buf (_39676_, _39201_);
  buf (_39677_, _39203_);
  buf (_39678_, _39204_);
  buf (_39680_, _39205_);
  buf (_39681_, _39206_);
  buf (_39682_, _39207_);
  buf (_39683_, _39209_);
  buf (_39684_, _39210_);
  buf (_40076_, _39980_);
  buf (_40240_, _39980_);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _05111_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _05115_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _05119_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _05123_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _05127_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _05131_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _05135_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _05105_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _05108_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _05163_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _05167_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _05171_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _05175_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _05179_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _05183_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _05186_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _05156_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _05159_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _05633_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _05637_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _05641_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _05645_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _05649_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _05653_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _05657_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _05626_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _05629_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _05686_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _05690_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _05694_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _05698_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _05702_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _05706_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _05710_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _05679_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _05682_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _05739_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _05743_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _05747_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _05751_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _05755_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _05759_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _05763_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _05732_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _05735_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _05792_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _05796_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _05800_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _05804_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _05808_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _05812_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _05816_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _05785_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _05788_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _05845_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _05849_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _05853_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _05857_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _05861_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _05865_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _05869_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _05838_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _05841_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _05898_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _05902_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _05906_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _05910_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _05914_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _05918_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _05922_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _05891_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _05894_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _05215_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _05219_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _05222_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _05226_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _05230_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _05234_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _05238_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _05208_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _05211_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _05266_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _05270_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _05274_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _05278_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _05282_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _05286_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _05290_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _05259_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _05262_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _05318_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _05322_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _05326_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _05329_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _05333_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _05337_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _05341_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _05311_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _05314_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _05369_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _05373_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _05377_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _05381_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _05385_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _05389_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _05393_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _05363_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _05365_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _05421_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _05425_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _05429_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _05433_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _05437_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _05441_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _05445_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _05414_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _05417_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _05474_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _05478_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _05482_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _05486_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _05490_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _05494_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _05498_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _05467_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _05470_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _05527_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _05531_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _05535_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _05539_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _05543_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _05547_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _05551_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _05520_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _05523_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _05580_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _05584_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _05588_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _05592_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _05596_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _05600_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _05604_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _05573_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _05576_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _41193_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _41194_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _41196_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _41197_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _41198_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _41199_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _41200_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _40979_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _41181_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _41182_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _41184_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _41185_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _41186_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _41187_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _41188_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _41190_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _41169_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _41170_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _41171_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _41173_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _41174_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _41175_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _41176_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _41177_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _41158_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _41159_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _41160_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _41162_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _41163_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _41164_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _41165_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _41166_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _41148_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _41149_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _41150_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _41151_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _41152_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _41153_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _41154_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _41155_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _41136_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _41137_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _41138_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _41139_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _41140_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _41142_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _41143_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _41144_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _41123_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _41124_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _41125_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _41126_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _41127_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _41128_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _41131_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _41132_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _41112_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _41114_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _41115_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _41116_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _41117_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _41118_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _41120_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _41121_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _41100_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _41101_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _41102_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _41103_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _41104_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _41106_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _41107_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _41108_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _41088_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _41089_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _41090_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _41091_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _41092_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _41094_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _41095_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _41096_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _41075_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _41077_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _41078_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _41079_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _41080_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _41081_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _41083_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _41084_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _41063_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _41066_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _41067_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _41068_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _41069_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _41070_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _41071_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _41072_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _41052_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _41053_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _41054_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _41055_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _41056_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _41058_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _41059_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _41060_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _41038_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _41041_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _41042_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _41043_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _41044_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _41045_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _41047_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _41048_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _41027_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _41028_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _41029_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _41030_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _41031_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _41033_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _41034_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _41035_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _41013_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _41014_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _41016_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _41017_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _41018_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _41020_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _41021_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _41022_);
  dff (\oc8051_golden_model_1.B [0], _43594_);
  dff (\oc8051_golden_model_1.B [1], _43595_);
  dff (\oc8051_golden_model_1.B [2], _43596_);
  dff (\oc8051_golden_model_1.B [3], _43598_);
  dff (\oc8051_golden_model_1.B [4], _43599_);
  dff (\oc8051_golden_model_1.B [5], _43600_);
  dff (\oc8051_golden_model_1.B [6], _43601_);
  dff (\oc8051_golden_model_1.B [7], _40980_);
  dff (\oc8051_golden_model_1.ACC [0], _43603_);
  dff (\oc8051_golden_model_1.ACC [1], _43604_);
  dff (\oc8051_golden_model_1.ACC [2], _43605_);
  dff (\oc8051_golden_model_1.ACC [3], _43606_);
  dff (\oc8051_golden_model_1.ACC [4], _43607_);
  dff (\oc8051_golden_model_1.ACC [5], _43608_);
  dff (\oc8051_golden_model_1.ACC [6], _43609_);
  dff (\oc8051_golden_model_1.ACC [7], _40981_);
  dff (\oc8051_golden_model_1.PCON [0], _43611_);
  dff (\oc8051_golden_model_1.PCON [1], _43612_);
  dff (\oc8051_golden_model_1.PCON [2], _43613_);
  dff (\oc8051_golden_model_1.PCON [3], _43614_);
  dff (\oc8051_golden_model_1.PCON [4], _43615_);
  dff (\oc8051_golden_model_1.PCON [5], _43617_);
  dff (\oc8051_golden_model_1.PCON [6], _43618_);
  dff (\oc8051_golden_model_1.PCON [7], _40982_);
  dff (\oc8051_golden_model_1.TMOD [0], _43619_);
  dff (\oc8051_golden_model_1.TMOD [1], _43621_);
  dff (\oc8051_golden_model_1.TMOD [2], _43622_);
  dff (\oc8051_golden_model_1.TMOD [3], _43623_);
  dff (\oc8051_golden_model_1.TMOD [4], _43624_);
  dff (\oc8051_golden_model_1.TMOD [5], _43625_);
  dff (\oc8051_golden_model_1.TMOD [6], _43626_);
  dff (\oc8051_golden_model_1.TMOD [7], _40983_);
  dff (\oc8051_golden_model_1.DPL [0], _43628_);
  dff (\oc8051_golden_model_1.DPL [1], _43629_);
  dff (\oc8051_golden_model_1.DPL [2], _43630_);
  dff (\oc8051_golden_model_1.DPL [3], _43631_);
  dff (\oc8051_golden_model_1.DPL [4], _43632_);
  dff (\oc8051_golden_model_1.DPL [5], _43633_);
  dff (\oc8051_golden_model_1.DPL [6], _43634_);
  dff (\oc8051_golden_model_1.DPL [7], _40985_);
  dff (\oc8051_golden_model_1.DPH [0], _43636_);
  dff (\oc8051_golden_model_1.DPH [1], _43637_);
  dff (\oc8051_golden_model_1.DPH [2], _43638_);
  dff (\oc8051_golden_model_1.DPH [3], _43640_);
  dff (\oc8051_golden_model_1.DPH [4], _43641_);
  dff (\oc8051_golden_model_1.DPH [5], _43642_);
  dff (\oc8051_golden_model_1.DPH [6], _43643_);
  dff (\oc8051_golden_model_1.DPH [7], _40986_);
  dff (\oc8051_golden_model_1.TL1 [0], _43645_);
  dff (\oc8051_golden_model_1.TL1 [1], _43646_);
  dff (\oc8051_golden_model_1.TL1 [2], _43647_);
  dff (\oc8051_golden_model_1.TL1 [3], _43648_);
  dff (\oc8051_golden_model_1.TL1 [4], _43649_);
  dff (\oc8051_golden_model_1.TL1 [5], _43650_);
  dff (\oc8051_golden_model_1.TL1 [6], _43651_);
  dff (\oc8051_golden_model_1.TL1 [7], _40987_);
  dff (\oc8051_golden_model_1.TL0 [0], _43653_);
  dff (\oc8051_golden_model_1.TL0 [1], _43654_);
  dff (\oc8051_golden_model_1.TL0 [2], _43655_);
  dff (\oc8051_golden_model_1.TL0 [3], _43656_);
  dff (\oc8051_golden_model_1.TL0 [4], _43657_);
  dff (\oc8051_golden_model_1.TL0 [5], _43659_);
  dff (\oc8051_golden_model_1.TL0 [6], _43660_);
  dff (\oc8051_golden_model_1.TL0 [7], _40988_);
  dff (\oc8051_golden_model_1.TCON [0], _43661_);
  dff (\oc8051_golden_model_1.TCON [1], _43663_);
  dff (\oc8051_golden_model_1.TCON [2], _43664_);
  dff (\oc8051_golden_model_1.TCON [3], _43665_);
  dff (\oc8051_golden_model_1.TCON [4], _43666_);
  dff (\oc8051_golden_model_1.TCON [5], _43667_);
  dff (\oc8051_golden_model_1.TCON [6], _43668_);
  dff (\oc8051_golden_model_1.TCON [7], _40989_);
  dff (\oc8051_golden_model_1.TH1 [0], _43670_);
  dff (\oc8051_golden_model_1.TH1 [1], _43671_);
  dff (\oc8051_golden_model_1.TH1 [2], _43672_);
  dff (\oc8051_golden_model_1.TH1 [3], _43673_);
  dff (\oc8051_golden_model_1.TH1 [4], _43674_);
  dff (\oc8051_golden_model_1.TH1 [5], _43675_);
  dff (\oc8051_golden_model_1.TH1 [6], _43676_);
  dff (\oc8051_golden_model_1.TH1 [7], _40991_);
  dff (\oc8051_golden_model_1.TH0 [0], _43678_);
  dff (\oc8051_golden_model_1.TH0 [1], _43679_);
  dff (\oc8051_golden_model_1.TH0 [2], _43680_);
  dff (\oc8051_golden_model_1.TH0 [3], _43682_);
  dff (\oc8051_golden_model_1.TH0 [4], _43683_);
  dff (\oc8051_golden_model_1.TH0 [5], _43684_);
  dff (\oc8051_golden_model_1.TH0 [6], _43685_);
  dff (\oc8051_golden_model_1.TH0 [7], _40992_);
  dff (\oc8051_golden_model_1.PC [0], _43687_);
  dff (\oc8051_golden_model_1.PC [1], _43689_);
  dff (\oc8051_golden_model_1.PC [2], _43690_);
  dff (\oc8051_golden_model_1.PC [3], _43691_);
  dff (\oc8051_golden_model_1.PC [4], _43692_);
  dff (\oc8051_golden_model_1.PC [5], _43693_);
  dff (\oc8051_golden_model_1.PC [6], _43694_);
  dff (\oc8051_golden_model_1.PC [7], _43695_);
  dff (\oc8051_golden_model_1.PC [8], _43696_);
  dff (\oc8051_golden_model_1.PC [9], _43697_);
  dff (\oc8051_golden_model_1.PC [10], _43698_);
  dff (\oc8051_golden_model_1.PC [11], _43700_);
  dff (\oc8051_golden_model_1.PC [12], _43701_);
  dff (\oc8051_golden_model_1.PC [13], _43702_);
  dff (\oc8051_golden_model_1.PC [14], _43703_);
  dff (\oc8051_golden_model_1.PC [15], _40993_);
  dff (\oc8051_golden_model_1.P2 [0], _43705_);
  dff (\oc8051_golden_model_1.P2 [1], _43706_);
  dff (\oc8051_golden_model_1.P2 [2], _43707_);
  dff (\oc8051_golden_model_1.P2 [3], _43708_);
  dff (\oc8051_golden_model_1.P2 [4], _43709_);
  dff (\oc8051_golden_model_1.P2 [5], _43710_);
  dff (\oc8051_golden_model_1.P2 [6], _43711_);
  dff (\oc8051_golden_model_1.P2 [7], _40994_);
  dff (\oc8051_golden_model_1.P3 [0], _43713_);
  dff (\oc8051_golden_model_1.P3 [1], _43714_);
  dff (\oc8051_golden_model_1.P3 [2], _43715_);
  dff (\oc8051_golden_model_1.P3 [3], _43716_);
  dff (\oc8051_golden_model_1.P3 [4], _43717_);
  dff (\oc8051_golden_model_1.P3 [5], _43719_);
  dff (\oc8051_golden_model_1.P3 [6], _43720_);
  dff (\oc8051_golden_model_1.P3 [7], _40995_);
  dff (\oc8051_golden_model_1.P0 [0], _43721_);
  dff (\oc8051_golden_model_1.P0 [1], _43723_);
  dff (\oc8051_golden_model_1.P0 [2], _43724_);
  dff (\oc8051_golden_model_1.P0 [3], _43725_);
  dff (\oc8051_golden_model_1.P0 [4], _43726_);
  dff (\oc8051_golden_model_1.P0 [5], _43727_);
  dff (\oc8051_golden_model_1.P0 [6], _43728_);
  dff (\oc8051_golden_model_1.P0 [7], _40997_);
  dff (\oc8051_golden_model_1.P1 [0], _43730_);
  dff (\oc8051_golden_model_1.P1 [1], _43731_);
  dff (\oc8051_golden_model_1.P1 [2], _43732_);
  dff (\oc8051_golden_model_1.P1 [3], _43733_);
  dff (\oc8051_golden_model_1.P1 [4], _43734_);
  dff (\oc8051_golden_model_1.P1 [5], _43735_);
  dff (\oc8051_golden_model_1.P1 [6], _43736_);
  dff (\oc8051_golden_model_1.P1 [7], _40998_);
  dff (\oc8051_golden_model_1.IP [0], _43738_);
  dff (\oc8051_golden_model_1.IP [1], _43739_);
  dff (\oc8051_golden_model_1.IP [2], _43740_);
  dff (\oc8051_golden_model_1.IP [3], _43742_);
  dff (\oc8051_golden_model_1.IP [4], _43743_);
  dff (\oc8051_golden_model_1.IP [5], _43744_);
  dff (\oc8051_golden_model_1.IP [6], _43745_);
  dff (\oc8051_golden_model_1.IP [7], _40999_);
  dff (\oc8051_golden_model_1.IE [0], _43747_);
  dff (\oc8051_golden_model_1.IE [1], _43748_);
  dff (\oc8051_golden_model_1.IE [2], _43749_);
  dff (\oc8051_golden_model_1.IE [3], _43750_);
  dff (\oc8051_golden_model_1.IE [4], _43751_);
  dff (\oc8051_golden_model_1.IE [5], _43752_);
  dff (\oc8051_golden_model_1.IE [6], _43753_);
  dff (\oc8051_golden_model_1.IE [7], _41000_);
  dff (\oc8051_golden_model_1.SCON [0], _43755_);
  dff (\oc8051_golden_model_1.SCON [1], _43756_);
  dff (\oc8051_golden_model_1.SCON [2], _43757_);
  dff (\oc8051_golden_model_1.SCON [3], _43758_);
  dff (\oc8051_golden_model_1.SCON [4], _43759_);
  dff (\oc8051_golden_model_1.SCON [5], _43761_);
  dff (\oc8051_golden_model_1.SCON [6], _43762_);
  dff (\oc8051_golden_model_1.SCON [7], _41001_);
  dff (\oc8051_golden_model_1.SP [0], _43763_);
  dff (\oc8051_golden_model_1.SP [1], _43765_);
  dff (\oc8051_golden_model_1.SP [2], _43766_);
  dff (\oc8051_golden_model_1.SP [3], _43767_);
  dff (\oc8051_golden_model_1.SP [4], _43768_);
  dff (\oc8051_golden_model_1.SP [5], _43769_);
  dff (\oc8051_golden_model_1.SP [6], _43770_);
  dff (\oc8051_golden_model_1.SP [7], _41003_);
  dff (\oc8051_golden_model_1.SBUF [0], _43772_);
  dff (\oc8051_golden_model_1.SBUF [1], _43773_);
  dff (\oc8051_golden_model_1.SBUF [2], _43774_);
  dff (\oc8051_golden_model_1.SBUF [3], _43775_);
  dff (\oc8051_golden_model_1.SBUF [4], _43776_);
  dff (\oc8051_golden_model_1.SBUF [5], _43777_);
  dff (\oc8051_golden_model_1.SBUF [6], _43778_);
  dff (\oc8051_golden_model_1.SBUF [7], _41004_);
  dff (\oc8051_golden_model_1.PSW [0], _43779_);
  dff (\oc8051_golden_model_1.PSW [1], _43780_);
  dff (\oc8051_golden_model_1.PSW [2], _43781_);
  dff (\oc8051_golden_model_1.PSW [3], _43783_);
  dff (\oc8051_golden_model_1.PSW [4], _43784_);
  dff (\oc8051_golden_model_1.PSW [5], _43785_);
  dff (\oc8051_golden_model_1.PSW [6], _43786_);
  dff (\oc8051_golden_model_1.PSW [7], _41005_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02839_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02851_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02873_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02897_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02919_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00957_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _02931_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00927_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _02944_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _02957_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _02969_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _02980_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _02994_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03006_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03020_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00976_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02359_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22218_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02546_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02703_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _02884_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03126_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03363_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03564_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03763_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _03958_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04057_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04156_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04250_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04349_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04447_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04546_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04645_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24376_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _39186_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _39188_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _39189_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _39190_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _39191_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _39192_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _39193_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _39173_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _39194_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _39195_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _39197_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _39198_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _39199_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _39200_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _39201_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _39174_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _39203_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _39204_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _39205_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _39206_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _39207_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _39209_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _39210_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _39176_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _34279_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _34282_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _09718_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _34284_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _34286_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _09721_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _34288_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _09724_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _34290_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _34292_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _34294_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _09727_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _34296_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _09730_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _09733_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09792_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09794_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _09697_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09797_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09800_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _09700_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _09803_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _09703_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _09806_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _09809_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _09812_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _09815_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _09818_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _09821_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _09824_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _09706_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _09709_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _34277_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _09715_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _09827_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _09712_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39980_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _40013_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _40014_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _40015_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _40016_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _40017_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _40018_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _40019_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _39981_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _40021_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _40022_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _40023_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _40024_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _40025_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _40026_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _40027_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _39982_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _40028_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _40029_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _40030_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _40032_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _40033_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _40034_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _40035_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _39983_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _40036_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _40037_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _40038_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _40039_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _40040_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _40041_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _40043_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _39985_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39558_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39559_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39560_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39561_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _39275_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _39347_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _39348_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _39349_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _39350_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _39351_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _39353_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _39354_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _39355_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _39356_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _39357_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _39358_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _39359_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _39360_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39361_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39362_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _39234_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39367_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39368_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39369_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39370_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39371_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39372_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39373_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39374_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39375_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39376_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39378_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39379_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39380_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39381_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39382_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _39235_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39562_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39563_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39564_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39565_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39567_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39568_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39569_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39570_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39571_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39572_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39573_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39574_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39575_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39576_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39578_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39579_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39580_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39581_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39582_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39583_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39584_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39585_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39586_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39587_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39589_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39590_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39591_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39592_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39593_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39594_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39595_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _39300_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _39273_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39596_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39598_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39599_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39600_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39601_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39602_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39604_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _39276_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39605_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39606_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39607_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39608_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39609_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39610_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39611_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _39277_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39612_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39613_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39615_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39616_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39617_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39618_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39619_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _39279_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _39280_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _39281_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39620_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39621_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39622_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39623_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39624_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39626_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39627_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _39282_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39628_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39629_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39630_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39631_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39632_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39633_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39634_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39635_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39636_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39637_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39638_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39639_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39640_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39641_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39642_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _39283_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39643_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39644_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39645_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39647_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39648_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39649_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39650_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39651_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39652_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39653_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39654_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39655_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39656_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39658_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39659_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _39285_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _39286_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _39288_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _39287_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39660_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39661_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39662_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39663_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39664_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39665_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39666_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _39290_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39667_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39669_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _39291_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39670_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39671_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39672_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39673_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39674_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39675_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39676_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _39292_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39677_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39678_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39680_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39681_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39682_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39683_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39684_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _39293_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _39294_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39685_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39686_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39687_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39688_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39689_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39691_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39692_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _39295_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _39297_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _39298_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39693_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39694_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _39299_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39696_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39698_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39699_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39700_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39702_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39703_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39704_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39707_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39708_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39709_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39710_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39711_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39714_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39716_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39717_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39718_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39719_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39720_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39721_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39722_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39724_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39725_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39726_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39727_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39728_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39729_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _39301_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39730_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39731_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39732_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39735_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39736_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39737_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _39302_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _39303_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _39305_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39738_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39739_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39740_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39741_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39742_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39743_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39744_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39746_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39748_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39750_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39751_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39752_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39753_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _39306_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _39307_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _39308_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _39309_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39754_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39755_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39757_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39758_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39759_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39760_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39761_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39762_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39763_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39764_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39765_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39766_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39768_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39769_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39770_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _39310_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _39311_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _40237_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _40258_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _40259_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _40260_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _40261_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _40262_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _40263_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _40264_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _40239_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _40240_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _40265_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _40266_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _40241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _02802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _02807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _02812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _02817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _02822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _02827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _02832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _02834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _02842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _02845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _02848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _02853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _02856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _02859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _02862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _02865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _02871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _02875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _02879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _02882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _02886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _02889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _02893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _02895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _02933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _02937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _02940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _02945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _02949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _02952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _02956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _02959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _02901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _02904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _02907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _02910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _02914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _02917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _02922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _02925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _02992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _02996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _03000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _03003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _03008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _02963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _02966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _02971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _02974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _02977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _02981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _02985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _02987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _02578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _05087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _05089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _05091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _05095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _05097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02567_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _40070_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _40156_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _40157_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _40158_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _40072_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _40073_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _40074_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _40159_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _40161_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _40162_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _40163_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _40164_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _40165_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _40166_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _40075_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _40076_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19875_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19886_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19898_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19910_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19922_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _18000_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08905_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08916_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08927_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08938_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08949_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08960_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08971_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06664_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13660_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13671_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13682_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13693_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13704_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13715_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12715_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13737_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13748_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13769_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13780_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13791_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _43104_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _43102_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _43100_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00131_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00137_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00142_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _43098_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00144_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _43096_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _43094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00146_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00148_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _43093_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _43091_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _43089_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _43087_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _43058_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _43056_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _43054_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _43052_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00157_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _43050_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00166_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _43048_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00175_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00177_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00179_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00181_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00183_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00186_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _43045_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _40808_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _40810_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _40812_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _40814_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _40816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _40818_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _40820_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _31130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _40821_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _40823_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _40825_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _40827_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _40829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _40831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _40833_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _31153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _40835_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _40837_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _40839_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _40841_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _40843_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _40845_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _40847_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _31176_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _40849_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _40851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _40852_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _40854_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _40856_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _40858_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _40860_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _31199_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17376_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17387_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17398_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17420_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17431_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15195_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09521_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10753_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10764_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09542_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _41311_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _41314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _41820_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _41822_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _41823_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _41825_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _41827_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _41829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _41831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _41317_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _41833_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _41835_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _41837_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _41839_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _41840_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _41842_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _41844_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _41320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _41323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _41326_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _41846_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _41848_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _41850_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _41852_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _41854_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _41855_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _41857_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _41329_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _41859_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _41861_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _41863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _41865_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _41867_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _41869_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _41870_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _41332_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _41335_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _41872_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _41874_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _41876_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _41877_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _41879_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _41881_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _41883_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _41338_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01636_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01639_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02112_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02114_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02116_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02117_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02121_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02123_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01642_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02124_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02126_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02128_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02131_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01645_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01648_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02137_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02142_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02144_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01654_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02166_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01660_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01213_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01215_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01217_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01223_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01224_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01226_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01228_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01230_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00568_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00544_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00546_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00552_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00554_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00557_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01232_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01234_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01236_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01238_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00562_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01240_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01242_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01244_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01246_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01248_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01252_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00565_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00576_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00579_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00581_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00584_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01259_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01261_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01263_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01265_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01267_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01269_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01273_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01275_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01277_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00587_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01279_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01281_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01283_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01285_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01287_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01291_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00589_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01304_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00592_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [0], \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [1], \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [2], \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [3], \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [4], \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [5], \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [6], \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [7], \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [0], \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [1], \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [2], \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [3], \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [4], \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [5], \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [6], \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [7], \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [0], \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [1], \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [2], \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [3], \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [4], \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [5], \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [6], \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [7], \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [0], \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [1], \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [2], \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [3], \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [4], \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [5], \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [6], \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [7], \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1237 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1237 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1237 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1257 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1257 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1257 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1276 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1276 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1288 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1288 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1348 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1348 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1348 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1364 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1364 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1364 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1380 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1380 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n1558 [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n1582 [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n1591 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n1747 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n1747 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n1747 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n1760 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n1760 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n1760 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n1773 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n1773 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n1773 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n1773 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n1773 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n1773 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n1789 [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n1801 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n1805 [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n1826 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n1832 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n1838 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n1844 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n1844 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n1909 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0994 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0994 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0994 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0994 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0994 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0994 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0994 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1090 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1090 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1090 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1090 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1092 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1092 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1092 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1092 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1094 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1094 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1094 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1094 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1095 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1095 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1095 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1095 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1096 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1096 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1096 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1096 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1097 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1097 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1097 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1097 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1098 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1098 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1098 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1098 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1099 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1099 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1099 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1099 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1100 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1100 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1100 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1100 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1147 , \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.n1175 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1176 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1176 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1176 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1176 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1176 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1176 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1176 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1176 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1176 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1177 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1177 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1177 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1177 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1177 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1177 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1177 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1177 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1177 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1178 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1178 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1178 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1178 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1178 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1178 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1178 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1178 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1179 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1180 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1181 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1181 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1181 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1182 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1183 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1183 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1184 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1184 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1184 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1184 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1184 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1184 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1184 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1184 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1211 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1211 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1211 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1211 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1211 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1211 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1211 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1211 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1211 [8], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1211 [9], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1211 [10], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1211 [11], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1211 [12], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.n1211 [13], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.n1211 [14], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.n1211 [15], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n1213 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1213 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1213 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1213 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1213 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1213 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1213 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1213 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1215 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1215 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1215 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1215 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1215 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1215 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1215 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1215 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1215 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1219 [8], \oc8051_golden_model_1.n1237 [7]);
  buf(\oc8051_golden_model_1.n1220 , \oc8051_golden_model_1.n1237 [7]);
  buf(\oc8051_golden_model_1.n1221 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1221 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1221 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1221 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1222 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1222 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1222 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1222 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1222 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1226 [4], \oc8051_golden_model_1.n1237 [6]);
  buf(\oc8051_golden_model_1.n1227 , \oc8051_golden_model_1.n1237 [6]);
  buf(\oc8051_golden_model_1.n1228 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1228 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1228 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1228 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1228 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1228 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1228 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1228 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1228 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1236 , \oc8051_golden_model_1.n1237 [2]);
  buf(\oc8051_golden_model_1.n1237 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1237 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1237 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1237 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1237 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1241 [8], \oc8051_golden_model_1.n1257 [7]);
  buf(\oc8051_golden_model_1.n1242 , \oc8051_golden_model_1.n1257 [7]);
  buf(\oc8051_golden_model_1.n1247 [4], \oc8051_golden_model_1.n1257 [6]);
  buf(\oc8051_golden_model_1.n1248 , \oc8051_golden_model_1.n1257 [6]);
  buf(\oc8051_golden_model_1.n1256 , \oc8051_golden_model_1.n1257 [2]);
  buf(\oc8051_golden_model_1.n1257 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1257 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1257 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1257 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1257 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1259 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1259 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1259 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1259 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1259 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1259 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1259 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1259 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1259 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1261 [8], \oc8051_golden_model_1.n1276 [7]);
  buf(\oc8051_golden_model_1.n1262 , \oc8051_golden_model_1.n1276 [7]);
  buf(\oc8051_golden_model_1.n1263 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1263 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1263 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1263 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1264 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.n1267 , \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.n1268 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1268 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1268 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1268 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1268 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1268 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1268 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1268 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1268 [8], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.n1276 [2]);
  buf(\oc8051_golden_model_1.n1276 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1276 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1276 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1276 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1276 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1276 [6], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.n1279 [8], \oc8051_golden_model_1.n1288 [7]);
  buf(\oc8051_golden_model_1.n1280 , \oc8051_golden_model_1.n1288 [7]);
  buf(\oc8051_golden_model_1.n1287 , \oc8051_golden_model_1.n1288 [2]);
  buf(\oc8051_golden_model_1.n1288 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1288 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1288 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1288 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1288 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1290 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1290 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1290 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1290 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1290 [4], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.n1290 [5], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.n1290 [6], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.n1290 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n1290 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1292 [8], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.n1293 , \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.n1294 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1294 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1294 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1294 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1294 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1296 [4], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.n1297 , \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.n1298 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n1305 , \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.n1306 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1306 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1306 [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.n1306 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1306 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1306 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1306 [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.n1306 [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.n1308 [4], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.n1309 , \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.n1310 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1310 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1310 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1310 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1310 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1310 [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.n1312 [8], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.n1313 , \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.n1320 , \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.n1321 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1321 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1321 [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.n1321 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1321 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1321 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1321 [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.n1322 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1322 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1322 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1322 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1322 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1325 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1325 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1325 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1325 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1325 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1325 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1325 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1325 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1326 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1326 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1326 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1326 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1326 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1326 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1326 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1326 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1326 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1327 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1327 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1327 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1327 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1327 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1327 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1327 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1327 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1328 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1329 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1329 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1329 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1329 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1329 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1329 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1329 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1329 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1330 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1330 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1333 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1335 [8], \oc8051_golden_model_1.n1348 [7]);
  buf(\oc8051_golden_model_1.n1336 , \oc8051_golden_model_1.n1348 [7]);
  buf(\oc8051_golden_model_1.n1337 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1337 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1337 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1337 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1337 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1339 [4], \oc8051_golden_model_1.n1348 [6]);
  buf(\oc8051_golden_model_1.n1340 , \oc8051_golden_model_1.n1348 [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.n1348 [2]);
  buf(\oc8051_golden_model_1.n1348 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1348 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1348 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1348 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1348 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1352 [8], \oc8051_golden_model_1.n1364 [7]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.n1364 [7]);
  buf(\oc8051_golden_model_1.n1355 [4], \oc8051_golden_model_1.n1364 [6]);
  buf(\oc8051_golden_model_1.n1356 , \oc8051_golden_model_1.n1364 [6]);
  buf(\oc8051_golden_model_1.n1363 , \oc8051_golden_model_1.n1364 [2]);
  buf(\oc8051_golden_model_1.n1364 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1364 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1364 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1364 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1364 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1368 [8], \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.n1369 , \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.n1371 [4], \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.n1372 , \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.n1379 , \oc8051_golden_model_1.n1380 [2]);
  buf(\oc8051_golden_model_1.n1380 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1380 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1380 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1380 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1380 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1384 [8], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.n1385 , \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.n1387 [4], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.n1388 , \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.n1395 , \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.n1396 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1396 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1396 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1396 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1396 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1556 , \oc8051_golden_model_1.n1558 [7]);
  buf(\oc8051_golden_model_1.n1557 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1557 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1557 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1557 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1557 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1557 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1557 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1558 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1558 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1558 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1558 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1558 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1558 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1558 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1581 , \oc8051_golden_model_1.n1582 [7]);
  buf(\oc8051_golden_model_1.n1582 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1582 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1582 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1582 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1582 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1582 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1582 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1589 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1589 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1589 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1589 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1590 , \oc8051_golden_model_1.n1591 [2]);
  buf(\oc8051_golden_model_1.n1591 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1591 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1591 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1591 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1591 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1591 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1591 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1735 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1738 , \oc8051_golden_model_1.n1747 [7]);
  buf(\oc8051_golden_model_1.n1740 , \oc8051_golden_model_1.n1747 [6]);
  buf(\oc8051_golden_model_1.n1746 , \oc8051_golden_model_1.n1747 [2]);
  buf(\oc8051_golden_model_1.n1747 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1747 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1747 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1747 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1747 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1751 , \oc8051_golden_model_1.n1760 [7]);
  buf(\oc8051_golden_model_1.n1753 , \oc8051_golden_model_1.n1760 [6]);
  buf(\oc8051_golden_model_1.n1759 , \oc8051_golden_model_1.n1760 [2]);
  buf(\oc8051_golden_model_1.n1760 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1760 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1760 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1760 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1760 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1764 , \oc8051_golden_model_1.n1773 [7]);
  buf(\oc8051_golden_model_1.n1766 , \oc8051_golden_model_1.n1773 [6]);
  buf(\oc8051_golden_model_1.n1772 , \oc8051_golden_model_1.n1773 [2]);
  buf(\oc8051_golden_model_1.n1773 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1773 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1773 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1773 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1773 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1777 , \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.n1779 , \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.n1785 , \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.n1786 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1786 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1786 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1786 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1786 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1788 , \oc8051_golden_model_1.n1789 [7]);
  buf(\oc8051_golden_model_1.n1789 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1789 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1789 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1789 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1789 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1789 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1789 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1790 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1790 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1790 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1790 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1790 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1790 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1790 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1794 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n1794 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n1794 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n1794 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n1794 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n1794 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n1794 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n1794 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n1794 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [9], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [10], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [11], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [12], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [13], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [14], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1800 , \oc8051_golden_model_1.n1801 [2]);
  buf(\oc8051_golden_model_1.n1801 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1801 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1801 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1801 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1801 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1801 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1801 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1804 , \oc8051_golden_model_1.n1805 [7]);
  buf(\oc8051_golden_model_1.n1805 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1805 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1805 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1805 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1805 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1805 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1805 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1825 , \oc8051_golden_model_1.n1826 [7]);
  buf(\oc8051_golden_model_1.n1826 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1826 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1826 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1826 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1826 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1826 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1826 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1831 , \oc8051_golden_model_1.n1832 [7]);
  buf(\oc8051_golden_model_1.n1832 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1832 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1832 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1832 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1832 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1832 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1832 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1837 , \oc8051_golden_model_1.n1838 [7]);
  buf(\oc8051_golden_model_1.n1838 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1838 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1838 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1838 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1838 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1838 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1838 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1843 , \oc8051_golden_model_1.n1844 [7]);
  buf(\oc8051_golden_model_1.n1844 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1844 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1844 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1844 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1844 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1844 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1844 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1849 , \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.n1850 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1850 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1850 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1850 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1850 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1850 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1850 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1851 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1851 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1851 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1851 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1851 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1851 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1851 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1851 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1852 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1852 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1852 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1852 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1853 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1853 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1853 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1853 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1853 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1853 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1889 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1889 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1889 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1889 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1889 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1889 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1889 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1889 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1908 , \oc8051_golden_model_1.n1909 [7]);
  buf(\oc8051_golden_model_1.n1909 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1909 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1909 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1909 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1909 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1909 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1909 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1913 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1913 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1913 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1913 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1914 [0], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1914 [1], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1914 [2], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1914 [3], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1915 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1915 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1915 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1915 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
