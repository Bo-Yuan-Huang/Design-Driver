
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_jc, ABINPUT, ABINPUT000, ABINPUT000000);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  input [8:0] ABINPUT;
  input [16:0] ABINPUT000;
  input [16:0] ABINPUT000000;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [16:0] \oc8051_top_1.ABINPUT000 ;
  wire [16:0] \oc8051_top_1.ABINPUT000000 ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT000 ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire \oc8051_top_1.oc8051_alu1.divOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.mulOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pc_log_change_r;
  output property_invalid_jc;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not (_05141_, rst);
  not (_05142_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  not (_05143_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_05144_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _05143_);
  and (_05145_, _05144_, _05142_);
  and (_05146_, _05145_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_05147_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  not (_05148_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_05149_, _05145_, _05148_);
  and (_05150_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_05151_, _05150_, _05147_);
  not (_05152_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  not (_05153_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nand (_05154_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  or (_05155_, _05154_, _05153_);
  and (_05156_, _05155_, _05152_);
  and (_05157_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05143_);
  and (_05158_, _05157_, _05148_);
  and (_05159_, _05158_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  or (_05160_, _05155_, _05152_);
  nand (_05161_, _05160_, _05159_);
  or (_05162_, _05161_, _05156_);
  nor (_05163_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  nor (_05164_, _05163_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_05165_, _05164_, _05144_);
  nand (_05166_, _05165_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  not (_05167_, _05158_);
  nor (_05168_, _05167_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  nand (_05169_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  and (_05170_, _05169_, _05166_);
  and (_05171_, _05170_, _05162_);
  and (_05172_, _05171_, _05151_);
  not (_05173_, _05172_);
  and (_05174_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_05175_, _05174_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_05176_, _05154_, _05153_);
  nor (_05177_, _05176_, _05175_);
  and (_05178_, _05177_, _05159_);
  and (_05179_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_05180_, _05179_, _05178_);
  and (_05181_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand (_05182_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  nand (_05183_, _05165_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  nand (_05184_, _05183_, _05182_);
  nor (_05185_, _05184_, _05181_);
  and (_05186_, _05185_, _05180_);
  and (_05187_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_05188_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_05189_, _05188_, _05187_);
  and (_05190_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not (_05191_, _05190_);
  not (_05192_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_05193_, _05159_, _05192_);
  and (_05194_, _05165_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_05195_, _05194_, _05193_);
  and (_05196_, _05195_, _05191_);
  and (_05197_, _05196_, _05189_);
  nor (_05198_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_05199_, _05198_, _05174_);
  and (_05200_, _05199_, _05159_);
  and (_05201_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_05202_, _05201_, _05200_);
  and (_05203_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand (_05204_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nand (_05205_, _05165_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  nand (_05206_, _05205_, _05204_);
  nor (_05207_, _05206_, _05203_);
  and (_05208_, _05207_, _05202_);
  and (_05209_, _05208_, _05197_);
  and (_05210_, _05209_, _05186_);
  and (_05211_, _05210_, _05173_);
  not (_05212_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_05213_, _05160_, _05212_);
  and (_05214_, _05213_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nand (_05215_, _05214_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  or (_05216_, _05214_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_05217_, _05216_, _05159_);
  nand (_05218_, _05217_, _05215_);
  nand (_05219_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_05220_, _05144_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  nand (_05221_, _05220_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_05222_, _05221_, _05219_);
  nand (_05223_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nand (_05224_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_05225_, _05224_, _05223_);
  and (_05226_, _05225_, _05222_);
  and (_05227_, _05226_, _05218_);
  not (_05228_, _05227_);
  nand (_05229_, _05215_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  or (_05230_, _05215_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand (_05231_, _05230_, _05229_);
  nand (_05232_, _05231_, _05159_);
  nand (_05233_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_05234_, _05233_, _05221_);
  nand (_05236_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nand (_05237_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_05239_, _05237_, _05236_);
  and (_05240_, _05239_, _05234_);
  nand (_05241_, _05240_, _05232_);
  nor (_05242_, _05241_, _05228_);
  not (_05243_, _05159_);
  and (_05244_, _05160_, _05212_);
  or (_05245_, _05244_, _05243_);
  or (_05246_, _05245_, _05213_);
  nand (_05247_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_05248_, _05247_, _05221_);
  nand (_05249_, _05165_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nand (_05250_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  and (_05252_, _05250_, _05249_);
  nand (_05253_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_05254_, _05253_, _05252_);
  and (_05255_, _05254_, _05248_);
  and (_05256_, _05255_, _05246_);
  or (_05257_, _05213_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_05258_, _05214_, _05243_);
  nand (_05259_, _05258_, _05257_);
  nand (_05260_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_05261_, _05260_, _05221_);
  nand (_05262_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  nand (_05263_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_05264_, _05263_, _05262_);
  and (_05265_, _05264_, _05261_);
  and (_05266_, _05265_, _05259_);
  and (_05267_, _05266_, _05256_);
  and (_05268_, _05267_, _05242_);
  and (_05269_, _05268_, _05211_);
  not (_05270_, _05269_);
  and (_05271_, _05186_, _05172_);
  and (_05272_, _05209_, _05271_);
  and (_05273_, _05272_, _05268_);
  not (_05274_, _05208_);
  nor (_05275_, _05274_, _05197_);
  and (_05276_, _05271_, _05275_);
  and (_05277_, _05268_, _05276_);
  nor (_05278_, _05277_, _05273_);
  and (_05279_, _05278_, _05270_);
  not (_05280_, _05266_);
  nor (_05281_, _05280_, _05256_);
  and (_05282_, _05281_, _05242_);
  and (_05283_, _05282_, _05276_);
  and (_05284_, _05211_, _05282_);
  nor (_05285_, _05284_, _05283_);
  not (_05286_, _05197_);
  and (_05287_, _05186_, _05208_);
  and (_05288_, _05287_, _05286_);
  and (_05289_, _05288_, _05173_);
  and (_05290_, _05289_, _05268_);
  and (_05291_, _05272_, _05282_);
  nor (_05292_, _05291_, _05290_);
  and (_05293_, _05292_, _05285_);
  and (_05294_, _05293_, _05279_);
  not (_05295_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_05296_, _05143_, \oc8051_top_1.oc8051_decoder1.wr );
  and (_05297_, _05296_, _05295_);
  nand (_05298_, _05297_, _05279_);
  or (_05299_, _05298_, _05294_);
  and (_05300_, _05299_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  not (_05301_, _05290_);
  nor (_05302_, _05291_, _05283_);
  nand (_05303_, _05302_, _05301_);
  and (_05305_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_05306_, _05305_, _05303_);
  not (_05307_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  not (_05308_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or (_05309_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_05310_, _05309_, _05308_);
  nor (_05311_, _05310_, _05307_);
  not (_05312_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nand (_05313_, _05308_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_05314_, _05313_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nor (_05315_, _05314_, _05312_);
  nor (_05316_, _05315_, _05311_);
  not (_05317_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_05318_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand (_05319_, _05318_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nor (_05320_, _05319_, _05317_);
  not (_05321_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_05322_, _05313_, _05321_);
  not (_05323_, _05322_);
  and (_05324_, _05323_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_05325_, _05324_, _05320_);
  and (_05326_, _05325_, _05316_);
  nor (_05327_, _05309_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  not (_05328_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_05330_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05328_);
  nor (_05331_, _05330_, ABINPUT[5]);
  nand (_05332_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05328_);
  nor (_05333_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor (_05334_, _05333_, _05331_);
  and (_05335_, _05334_, _05327_);
  and (_05336_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_05337_, _05336_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_05338_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  not (_05339_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_05341_, _05336_, _05321_);
  nor (_05342_, _05341_, _05339_);
  nor (_05343_, _05342_, _05338_);
  not (_05344_, _05343_);
  nor (_05345_, _05344_, _05335_);
  and (_05346_, _05345_, _05326_);
  and (_05347_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _05143_);
  and (_05348_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _05143_);
  nor (_05349_, _05348_, _05347_);
  not (_05350_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or (_05351_, _05350_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_05352_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _05143_);
  not (_05353_, _05352_);
  and (_05354_, _05353_, _05351_);
  and (_05355_, _05354_, _05349_);
  not (_05356_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_05357_, _05347_, _05356_);
  nand (_05358_, _05357_, _05350_);
  nand (_05359_, _05349_, _05352_);
  nand (_05360_, _05359_, _05358_);
  nor (_05361_, _05360_, _05355_);
  and (_05362_, _05348_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_05363_, _05362_, _05350_);
  not (_05364_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_05365_, _05348_, _05364_);
  not (_05366_, _05365_);
  nor (_05367_, _05366_, _05351_);
  nor (_05368_, _05367_, _05363_);
  and (_05370_, _05368_, _05361_);
  nor (_05371_, _05370_, _05346_);
  not (_05372_, _05371_);
  not (_05373_, _05346_);
  and (_05374_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_05375_, _05374_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_05376_, _05375_);
  or (_05377_, _05330_, ABINPUT[0]);
  or (_05378_, _05332_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_05379_, _05378_, _05377_);
  or (_05380_, _05379_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_05381_, _05380_, _05376_);
  not (_05382_, _05381_);
  not (_05383_, _05310_);
  and (_05384_, _05383_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  not (_05385_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_05386_, _05314_, _05385_);
  nor (_05387_, _05386_, _05384_);
  not (_05388_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_05389_, _05322_, _05388_);
  not (_05390_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_05391_, _05319_, _05390_);
  nor (_05392_, _05391_, _05389_);
  and (_05393_, _05392_, _05387_);
  not (_05394_, _05327_);
  or (_05395_, _05330_, ABINPUT[4]);
  or (_05396_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_05397_, _05396_, _05395_);
  or (_05398_, _05397_, _05394_);
  not (_05399_, _05341_);
  and (_05400_, _05399_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_05401_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_05402_, _05401_, _05400_);
  and (_05403_, _05402_, _05398_);
  and (_05404_, _05403_, _05393_);
  not (_05405_, _05404_);
  not (_05406_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or (_05407_, _05314_, _05406_);
  not (_05408_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  or (_05409_, _05310_, _05408_);
  and (_05410_, _05409_, _05407_);
  not (_05411_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_05412_, _05319_, _05411_);
  nand (_05413_, _05323_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_05414_, _05413_, _05412_);
  and (_05415_, _05414_, _05410_);
  or (_05416_, _05330_, ABINPUT[1]);
  or (_05417_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_05418_, _05417_, _05416_);
  or (_05419_, _05418_, _05394_);
  not (_05420_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_05421_, _05341_, _05420_);
  nand (_05422_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_05423_, _05422_, _05421_);
  and (_05424_, _05423_, _05419_);
  and (_05425_, _05424_, _05415_);
  or (_05426_, _05330_, ABINPUT[2]);
  or (_05427_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_05428_, _05427_, _05426_);
  or (_05429_, _05428_, _05394_);
  not (_05430_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_05431_, _05314_, _05430_);
  not (_05432_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  or (_05433_, _05310_, _05432_);
  and (_05434_, _05433_, _05431_);
  and (_05435_, _05434_, _05429_);
  not (_05436_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_05437_, _05319_, _05436_);
  not (_05438_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_05439_, _05322_, _05438_);
  and (_05440_, _05439_, _05437_);
  not (_05441_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_05442_, _05341_, _05441_);
  nand (_05443_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_05444_, _05443_, _05442_);
  and (_05445_, _05444_, _05440_);
  and (_05446_, _05445_, _05435_);
  not (_05447_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_05448_, _05314_, _05447_);
  not (_05449_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  or (_05450_, _05310_, _05449_);
  and (_05452_, _05450_, _05448_);
  not (_05453_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_05454_, _05322_, _05453_);
  not (_05455_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_05456_, _05319_, _05455_);
  and (_05457_, _05456_, _05454_);
  and (_05458_, _05457_, _05452_);
  or (_05459_, _05330_, ABINPUT[3]);
  or (_05460_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_05461_, _05460_, _05459_);
  or (_05462_, _05461_, _05394_);
  nand (_05463_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  not (_05464_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_05465_, _05341_, _05464_);
  and (_05466_, _05465_, _05463_);
  and (_05467_, _05466_, _05462_);
  and (_05469_, _05467_, _05458_);
  and (_05470_, _05469_, _05446_);
  nand (_05471_, _05470_, _05425_);
  or (_05472_, _05471_, _05405_);
  or (_05473_, _05472_, _05382_);
  or (_05474_, _05446_, _05425_);
  nor (_05475_, _05474_, _05469_);
  nand (_05476_, _05475_, _05405_);
  or (_05477_, _05476_, _05381_);
  nand (_05478_, _05477_, _05473_);
  nand (_05479_, _05478_, _05373_);
  nor (_05480_, _05351_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_05481_, _05362_, _05480_);
  or (_05482_, _05478_, _05373_);
  and (_05483_, _05482_, _05481_);
  nand (_05484_, _05483_, _05479_);
  and (_05485_, _05365_, _05354_);
  nor (_05486_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_05487_, _05486_, _05334_);
  not (_05488_, _05487_);
  and (_05489_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_05490_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not (_05491_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_05492_, _05491_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_05493_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_05494_, _05493_, _05490_);
  and (_05495_, _05494_, _05488_);
  nor (_05496_, _05495_, _05346_);
  and (_05497_, _05495_, _05346_);
  nor (_05498_, _05497_, _05496_);
  nand (_05499_, _05498_, _05485_);
  and (_05500_, _05352_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_05501_, _05500_, _05357_);
  and (_05503_, _05501_, _05496_);
  and (_05504_, _05480_, _05357_);
  and (_05505_, _05504_, _05346_);
  nor (_05506_, _05505_, _05503_);
  and (_05507_, _05382_, _05346_);
  not (_05508_, _05507_);
  and (_05509_, _05362_, _05500_);
  not (_05510_, _05509_);
  and (_05511_, _05495_, _05381_);
  nor (_05512_, _05511_, _05510_);
  and (_05513_, _05512_, _05508_);
  and (_05514_, _05352_, _05350_);
  and (_05515_, _05365_, _05514_);
  not (_05516_, _05515_);
  nor (_05517_, _05516_, _05497_);
  nor (_05518_, _05517_, _05513_);
  and (_05519_, _05518_, _05506_);
  and (_05520_, _05519_, _05499_);
  and (_05521_, _05520_, _05484_);
  nand (_05522_, _05521_, _05372_);
  and (_05523_, _05297_, _05284_);
  and (_05524_, _05523_, _05522_);
  or (_05525_, _05524_, _05306_);
  or (_05526_, _05525_, _05300_);
  and (_09109_, _05526_, _05141_);
  not (_05527_, _05486_);
  or (_05528_, _05527_, _05461_);
  and (_05529_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_05530_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_05531_, _05530_, _05529_);
  and (_05532_, _05531_, _05528_);
  nor (_05533_, _05532_, _05510_);
  not (_05534_, _05469_);
  nand (_05535_, _05424_, _05415_);
  and (_05536_, _05535_, _05381_);
  nand (_05537_, _05445_, _05435_);
  or (_05538_, _05537_, _05382_);
  and (_05539_, _05538_, _05474_);
  nor (_05540_, _05539_, _05536_);
  nand (_05541_, _05540_, _05534_);
  or (_05542_, _05540_, _05534_);
  and (_05543_, _05542_, _05481_);
  and (_05544_, _05543_, _05541_);
  nor (_05545_, _05544_, _05533_);
  nor (_05546_, _05469_, _05370_);
  not (_05547_, _05546_);
  nor (_05548_, _05532_, _05469_);
  and (_05549_, _05548_, _05501_);
  and (_05550_, _05504_, _05469_);
  nor (_05551_, _05550_, _05549_);
  and (_05552_, _05532_, _05469_);
  nor (_05553_, _05552_, _05548_);
  and (_05554_, _05553_, _05485_);
  nor (_05555_, _05552_, _05516_);
  nor (_05556_, _05555_, _05554_);
  and (_05557_, _05556_, _05551_);
  and (_05559_, _05557_, _05547_);
  and (_05560_, _05559_, _05545_);
  not (_05561_, _05560_);
  and (_05562_, _05561_, _05284_);
  or (_05563_, _05303_, _05299_);
  and (_05564_, _05563_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or (_05565_, _05564_, _05562_);
  or (_05566_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_05567_, _05566_, _05141_);
  and (_10437_, _05567_, _05565_);
  not (_05568_, _05291_);
  nand (_05569_, _05568_, _05285_);
  and (_05570_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_05571_, _05570_, _05569_);
  not (_05572_, _05297_);
  nand (_05573_, _05282_, _05287_);
  or (_05574_, _05573_, _05572_);
  and (_05575_, _05574_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_05576_, _05289_, _05282_);
  or (_05577_, _05527_, _05418_);
  nand (_05578_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nand (_05579_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_05580_, _05579_, _05578_);
  and (_05581_, _05580_, _05577_);
  and (_05582_, _05581_, _05425_);
  not (_05583_, _05485_);
  not (_05584_, _05581_);
  and (_05585_, _05584_, _05535_);
  or (_05586_, _05585_, _05583_);
  and (_05587_, _05586_, _05516_);
  or (_05588_, _05587_, _05582_);
  not (_05589_, _05501_);
  or (_05590_, _05581_, _05425_);
  or (_05591_, _05590_, _05589_);
  not (_05592_, _05504_);
  or (_05593_, _05592_, _05535_);
  and (_05594_, _05593_, _05591_);
  or (_05595_, _05581_, _05510_);
  not (_05597_, _05481_);
  or (_05598_, _05597_, _05535_);
  and (_05600_, _05598_, _05595_);
  or (_05601_, _05425_, _05370_);
  and (_05602_, _05601_, _05600_);
  and (_05603_, _05602_, _05594_);
  and (_05604_, _05603_, _05588_);
  nor (_05605_, _05604_, _05572_);
  and (_05606_, _05605_, _05576_);
  or (_05607_, _05606_, _05575_);
  or (_05608_, _05607_, _05571_);
  and (_00002_, _05608_, _05141_);
  and (_05609_, _05292_, _05270_);
  not (_05610_, _05609_);
  nand (_05611_, _05268_, _05287_);
  and (_05612_, _05611_, _05302_);
  nand (_05613_, _05297_, _05278_);
  or (_05614_, _05613_, _05612_);
  or (_05615_, _05614_, _05610_);
  and (_05616_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_05617_, _05297_, _05283_);
  and (_05618_, _05617_, _05522_);
  or (_05619_, _05618_, _05616_);
  and (_02660_, _05619_, _05141_);
  and (_05620_, _05605_, _05290_);
  not (_05621_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_05622_, _05297_, _05290_);
  nor (_05623_, _05622_, _05621_);
  or (_05624_, _05623_, _05620_);
  and (_06673_, _05624_, _05141_);
  nor (_05625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_05626_, _05625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  not (_05627_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_05628_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_05629_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_05630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_05631_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _05630_);
  nor (_05632_, _05631_, _05629_);
  nor (_05633_, _05632_, _05628_);
  nor (_05634_, _05633_, _05627_);
  and (_05635_, _05630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_05636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_05637_, _05636_, _05635_);
  and (_05638_, _05637_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_05639_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_05640_, _05630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor (_05641_, _05640_, _05639_);
  and (_05642_, _05641_, _05638_);
  nand (_05643_, _05642_, _05634_);
  and (_05644_, _05643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nor (_05645_, _05644_, _05626_);
  and (_05646_, _05296_, _05167_);
  and (_05647_, _05646_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_05648_, _05241_, _05227_);
  and (_05649_, _05648_, _05267_);
  nor (_05650_, _05208_, _05197_);
  nor (_05651_, _05186_, _05172_);
  and (_05652_, _05651_, _05650_);
  and (_05653_, _05652_, _05649_);
  and (_05654_, _05653_, _05647_);
  or (_05655_, _05654_, _05645_);
  and (_05656_, _05480_, _05349_);
  not (_05657_, _05656_);
  not (_05658_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_05659_, _05310_, _05658_);
  not (_05660_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_05661_, _05314_, _05660_);
  nor (_05662_, _05661_, _05659_);
  not (_05663_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_05664_, _05319_, _05663_);
  not (_05665_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_05666_, _05322_, _05665_);
  nor (_05667_, _05666_, _05664_);
  and (_05668_, _05667_, _05662_);
  nor (_05669_, _05330_, ABINPUT[8]);
  nor (_05670_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nor (_05671_, _05670_, _05669_);
  and (_05672_, _05671_, _05327_);
  not (_05673_, _05672_);
  and (_05674_, _05399_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_05675_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_05676_, _05675_, _05674_);
  and (_05677_, _05676_, _05673_);
  and (_05678_, _05677_, _05668_);
  and (_05679_, _05671_, _05486_);
  not (_05680_, _05679_);
  and (_05681_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_05682_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_05683_, _05682_, _05681_);
  and (_05684_, _05683_, _05680_);
  not (_05685_, _05684_);
  and (_05686_, _05685_, _05678_);
  nor (_05688_, _05684_, _05678_);
  and (_05689_, _05684_, _05678_);
  nor (_05691_, _05689_, _05688_);
  not (_05692_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_05693_, _05314_, _05692_);
  not (_05694_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor (_05695_, _05310_, _05694_);
  nor (_05696_, _05695_, _05693_);
  and (_05697_, _05323_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_05699_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_05700_, _05319_, _05699_);
  nor (_05701_, _05700_, _05697_);
  and (_05702_, _05701_, _05696_);
  nor (_05703_, _05330_, ABINPUT[7]);
  nor (_05704_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nor (_05705_, _05704_, _05703_);
  and (_05706_, _05705_, _05327_);
  not (_05708_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_05709_, _05341_, _05708_);
  and (_05710_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_05711_, _05710_, _05709_);
  not (_05712_, _05711_);
  nor (_05713_, _05712_, _05706_);
  and (_05715_, _05713_, _05702_);
  not (_05716_, _05715_);
  and (_05718_, _05705_, _05486_);
  not (_05719_, _05718_);
  and (_05721_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_05722_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_05723_, _05722_, _05721_);
  and (_05724_, _05723_, _05719_);
  and (_05725_, _05724_, _05716_);
  nor (_05727_, _05724_, _05715_);
  and (_05728_, _05724_, _05715_);
  nor (_05730_, _05728_, _05727_);
  not (_05731_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_05733_, _05314_, _05731_);
  not (_05734_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor (_05736_, _05310_, _05734_);
  nor (_05737_, _05736_, _05733_);
  not (_05739_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_05740_, _05319_, _05739_);
  not (_05742_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_05743_, _05322_, _05742_);
  nor (_05745_, _05743_, _05740_);
  and (_05746_, _05745_, _05737_);
  nor (_05747_, _05330_, ABINPUT[6]);
  nor (_05748_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nor (_05749_, _05748_, _05747_);
  and (_05750_, _05749_, _05327_);
  not (_05751_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_05752_, _05341_, _05751_);
  and (_05753_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  nor (_05754_, _05753_, _05752_);
  not (_05755_, _05754_);
  nor (_05757_, _05755_, _05750_);
  and (_05758_, _05757_, _05746_);
  not (_05759_, _05758_);
  and (_05761_, _05749_, _05486_);
  not (_05762_, _05761_);
  and (_05763_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_05765_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_05766_, _05765_, _05763_);
  and (_05768_, _05766_, _05762_);
  and (_05769_, _05768_, _05759_);
  not (_05771_, _05495_);
  and (_05772_, _05771_, _05346_);
  nor (_05773_, _05768_, _05758_);
  and (_05774_, _05768_, _05758_);
  nor (_05775_, _05774_, _05773_);
  nor (_05776_, _05775_, _05772_);
  nor (_05777_, _05776_, _05769_);
  nor (_05778_, _05777_, _05730_);
  nor (_05779_, _05778_, _05725_);
  and (_05781_, _05777_, _05730_);
  nor (_05782_, _05781_, _05778_);
  and (_05784_, _05775_, _05772_);
  nor (_05785_, _05784_, _05776_);
  not (_05786_, _05785_);
  not (_05787_, _05498_);
  nor (_05788_, _05527_, _05397_);
  not (_05789_, _05788_);
  and (_05791_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_05792_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_05794_, _05792_, _05791_);
  and (_05795_, _05794_, _05789_);
  nor (_05796_, _05795_, _05404_);
  and (_05797_, _05795_, _05404_);
  nor (_05798_, _05797_, _05796_);
  not (_05799_, _05532_);
  nor (_05800_, _05799_, _05469_);
  not (_05801_, _05553_);
  and (_05802_, _05584_, _05425_);
  or (_05803_, _05527_, _05428_);
  nand (_05804_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand (_05805_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_05806_, _05805_, _05804_);
  and (_05807_, _05806_, _05803_);
  and (_05808_, _05807_, _05446_);
  nand (_05809_, _05806_, _05803_);
  and (_05810_, _05809_, _05537_);
  nor (_05811_, _05810_, _05808_);
  or (_05812_, _05811_, _05802_);
  or (_05813_, _05809_, _05446_);
  nand (_05814_, _05813_, _05812_);
  and (_05815_, _05814_, _05801_);
  nor (_05816_, _05815_, _05800_);
  nor (_05817_, _05816_, _05798_);
  and (_05818_, _05816_, _05798_);
  or (_05819_, _05818_, _05817_);
  nor (_05820_, _05814_, _05801_);
  or (_05821_, _05820_, _05815_);
  and (_05822_, _05811_, _05802_);
  not (_05823_, _05822_);
  nand (_05824_, _05823_, _05812_);
  nor (_05825_, _05585_, _05582_);
  nor (_05826_, _05825_, _05382_);
  and (_05827_, _05826_, _05824_);
  and (_05828_, _05827_, _05821_);
  and (_05829_, _05828_, _05819_);
  not (_05830_, _05795_);
  or (_05831_, _05830_, _05404_);
  and (_05832_, _05830_, _05404_);
  or (_05833_, _05816_, _05832_);
  and (_05834_, _05833_, _05831_);
  or (_05835_, _05834_, _05829_);
  and (_05836_, _05835_, _05787_);
  and (_05837_, _05836_, _05786_);
  not (_05838_, _05837_);
  nor (_05839_, _05838_, _05782_);
  nor (_05840_, _05839_, _05779_);
  nor (_05841_, _05840_, _05691_);
  nor (_05842_, _05841_, _05686_);
  or (_05843_, _05842_, _05657_);
  and (_05844_, _05514_, _05349_);
  not (_05845_, _05844_);
  not (_05846_, _05688_);
  not (_05847_, _05548_);
  and (_05848_, _05811_, _05585_);
  or (_05849_, _05848_, _05810_);
  nand (_05850_, _05849_, _05553_);
  nand (_05851_, _05850_, _05847_);
  or (_05852_, _05851_, _05798_);
  nand (_05853_, _05851_, _05798_);
  and (_05854_, _05853_, _05852_);
  and (_05855_, _05825_, _05381_);
  and (_05856_, _05855_, _05811_);
  or (_05857_, _05849_, _05553_);
  and (_05858_, _05857_, _05850_);
  and (_05859_, _05858_, _05856_);
  and (_05860_, _05859_, _05854_);
  not (_05861_, _05797_);
  and (_05862_, _05851_, _05861_);
  or (_05863_, _05862_, _05796_);
  or (_05864_, _05863_, _05860_);
  nand (_05865_, _05864_, _05498_);
  and (_05866_, _05775_, _05496_);
  nor (_05867_, _05775_, _05496_);
  nor (_05868_, _05867_, _05866_);
  not (_05869_, _05868_);
  or (_05870_, _05869_, _05865_);
  not (_05871_, _05730_);
  nor (_05872_, _05866_, _05773_);
  nor (_05873_, _05872_, _05871_);
  and (_05874_, _05872_, _05871_);
  nor (_05875_, _05874_, _05873_);
  not (_05876_, _05875_);
  or (_05877_, _05876_, _05870_);
  nor (_05878_, _05873_, _05727_);
  and (_05879_, _05878_, _05877_);
  or (_05880_, _05879_, _05689_);
  and (_05881_, _05880_, _05846_);
  or (_05882_, _05881_, _05845_);
  and (_05883_, _05514_, _05357_);
  and (_05884_, _05758_, _05715_);
  nor (_05885_, _05884_, _05678_);
  and (_05886_, _05885_, _05382_);
  nor (_05887_, _05470_, _05404_);
  nor (_05888_, _05885_, _05382_);
  or (_05889_, _05888_, _05887_);
  or (_05890_, _05889_, _05886_);
  and (_05891_, _05890_, _05883_);
  and (_05892_, _05365_, _05500_);
  not (_05893_, _05892_);
  nor (_05894_, _05678_, _05893_);
  and (_05895_, _05379_, _05375_);
  and (_05896_, _05365_, _05480_);
  and (_05897_, _05501_, _05379_);
  nor (_05898_, _05897_, _05896_);
  nor (_05899_, _05898_, _05895_);
  nor (_05900_, _05899_, _05894_);
  nor (_05901_, _05381_, _05379_);
  and (_05902_, _05379_, _05376_);
  nor (_05903_, _05902_, _05583_);
  nor (_05904_, _05903_, _05515_);
  nor (_05905_, _05904_, _05901_);
  not (_05906_, _05905_);
  and (_05907_, _05362_, _05514_);
  and (_05908_, _05535_, _05907_);
  and (_05909_, _05362_, _05354_);
  not (_05910_, _05379_);
  and (_05911_, _05910_, _05909_);
  nor (_05912_, _05911_, _05355_);
  and (_05913_, _05912_, _05381_);
  nor (_05914_, _05504_, _05381_);
  nor (_05915_, _05914_, _05913_);
  nor (_05916_, _05915_, _05908_);
  and (_05917_, _05916_, _05906_);
  and (_05918_, _05917_, _05900_);
  not (_05919_, _05918_);
  nor (_05920_, _05919_, _05891_);
  and (_05921_, _05920_, _05882_);
  nand (_05922_, _05921_, _05843_);
  nand (_05923_, _05654_, _05922_);
  and (_05924_, _05923_, _05655_);
  and (_05925_, _05297_, _05167_);
  and (_05926_, _05925_, _05211_);
  and (_05927_, _05926_, _05649_);
  not (_05928_, _05927_);
  nand (_05929_, _05928_, _05924_);
  and (_05930_, _05678_, _05382_);
  not (_05931_, _05930_);
  and (_05933_, _05684_, _05381_);
  nor (_05934_, _05933_, _05510_);
  and (_05935_, _05934_, _05931_);
  not (_05936_, _05678_);
  nor (_05937_, _05472_, _05373_);
  and (_05938_, _05884_, _05937_);
  nor (_05939_, _05938_, _05382_);
  nor (_05940_, _05476_, _05346_);
  and (_05941_, _05940_, _05759_);
  nand (_05942_, _05941_, _05716_);
  and (_05943_, _05942_, _05382_);
  nor (_05944_, _05943_, _05939_);
  and (_05945_, _05944_, _05936_);
  nor (_05946_, _05944_, _05936_);
  nor (_05947_, _05946_, _05945_);
  and (_05948_, _05947_, _05481_);
  nor (_05949_, _05948_, _05935_);
  and (_05950_, _05691_, _05485_);
  and (_05951_, _05688_, _05501_);
  nor (_05952_, _05689_, _05516_);
  and (_05953_, _05678_, _05504_);
  or (_05954_, _05953_, _05952_);
  or (_05955_, _05954_, _05951_);
  nor (_05956_, _05955_, _05950_);
  nor (_05957_, _05678_, _05370_);
  not (_05958_, _05957_);
  and (_05959_, _05958_, _05956_);
  and (_05960_, _05959_, _05949_);
  nand (_05961_, _05960_, _05927_);
  and (_05962_, _05961_, _05141_);
  and (_07206_, _05962_, _05929_);
  not (_05963_, _05922_);
  and (_05964_, _05651_, _05275_);
  and (_05965_, _05964_, _05649_);
  and (_05966_, _05965_, _05647_);
  nand (_05967_, _05966_, _05963_);
  not (_05968_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_05969_, _05968_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not (_05970_, _05634_);
  nor (_05971_, _05641_, _05628_);
  not (_05972_, _05971_);
  or (_05973_, _05972_, _05638_);
  or (_05974_, _05973_, _05970_);
  and (_05975_, _05974_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_05976_, _05975_, _05969_);
  or (_05977_, _05976_, _05966_);
  and (_05978_, _05977_, _05928_);
  and (_05979_, _05978_, _05967_);
  nor (_05980_, _05758_, _05381_);
  nor (_05981_, _05768_, _05382_);
  or (_05982_, _05981_, _05980_);
  and (_05983_, _05982_, _05509_);
  not (_05984_, _05937_);
  nand (_05985_, _05984_, _05477_);
  and (_05986_, _05985_, _05508_);
  nand (_05987_, _05986_, _05759_);
  or (_05988_, _05986_, _05759_);
  and (_05989_, _05988_, _05481_);
  and (_05990_, _05989_, _05987_);
  nor (_05991_, _05990_, _05983_);
  nor (_05992_, _05758_, _05370_);
  not (_05993_, _05992_);
  and (_05994_, _05775_, _05485_);
  not (_05995_, _05994_);
  nor (_05996_, _05774_, _05516_);
  not (_05997_, _05996_);
  and (_05998_, _05773_, _05501_);
  and (_05999_, _05758_, _05504_);
  nor (_06000_, _05999_, _05998_);
  and (_06001_, _06000_, _05997_);
  and (_06002_, _06001_, _05995_);
  and (_06003_, _06002_, _05993_);
  nand (_06004_, _06003_, _05991_);
  and (_06005_, _06004_, _05927_);
  or (_06006_, _06005_, _05979_);
  and (_07277_, _06006_, _05141_);
  not (_06007_, _05186_);
  and (_06008_, _05650_, _06007_);
  and (_06009_, _05280_, _05227_);
  and (_06010_, _05647_, _05241_);
  nor (_06011_, _05256_, _05172_);
  and (_06012_, _06011_, _06010_);
  and (_06013_, _06012_, _06009_);
  and (_06014_, _06013_, _06008_);
  nand (_06015_, _06014_, _05963_);
  nor (_06016_, _05266_, _05256_);
  and (_06017_, _06016_, _05648_);
  and (_06018_, _05925_, _05172_);
  and (_06019_, _06018_, _06008_);
  and (_06020_, _06019_, _06017_);
  not (_06021_, _06020_);
  or (_06022_, _06014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_06023_, _06022_, _06021_);
  and (_06024_, _06023_, _06015_);
  nor (_06025_, _06021_, _05960_);
  or (_06026_, _06025_, _06024_);
  and (_07297_, _06026_, _05141_);
  and (_06027_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand (_06028_, _05633_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_06030_, _06028_, _05973_);
  and (_06031_, _06030_, _06027_);
  and (_06032_, _05650_, _05186_);
  and (_06033_, _06032_, _05173_);
  and (_06034_, _06033_, _05649_);
  and (_06035_, _06034_, _05647_);
  or (_06036_, _06035_, _06031_);
  and (_06037_, _06036_, _05928_);
  nand (_06038_, _06035_, _05963_);
  and (_06039_, _06038_, _06037_);
  nor (_06040_, _05795_, _05510_);
  nand (_06041_, _05471_, _05381_);
  or (_06042_, _05475_, _05381_);
  nand (_06043_, _06042_, _06041_);
  nand (_06044_, _06043_, _05404_);
  or (_06045_, _06043_, _05404_);
  and (_06046_, _06045_, _05481_);
  and (_06047_, _06046_, _06044_);
  nor (_06048_, _06047_, _06040_);
  nor (_06049_, _05404_, _05370_);
  not (_06050_, _06049_);
  and (_06051_, _05798_, _05485_);
  not (_06052_, _06051_);
  nor (_06053_, _05797_, _05516_);
  not (_06054_, _06053_);
  and (_06055_, _05796_, _05501_);
  and (_06056_, _05504_, _05404_);
  nor (_06057_, _06056_, _06055_);
  and (_06059_, _06057_, _06054_);
  and (_06060_, _06059_, _06052_);
  and (_06061_, _06060_, _06050_);
  and (_06062_, _06061_, _06048_);
  nor (_06063_, _06062_, _05928_);
  or (_06064_, _06063_, _06039_);
  and (_07616_, _06064_, _05141_);
  and (_06065_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_06066_, _06065_);
  and (_06067_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _05630_);
  and (_06068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_06069_, _06068_, _06067_);
  and (_06070_, _06069_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_06071_, _06070_, _05628_);
  and (_06072_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_06073_, _06072_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_06074_, _06073_);
  and (_06075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_06076_, _06075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_06077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_06078_, _06077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_06080_, _06078_, _06076_);
  and (_06081_, _06080_, _06074_);
  not (_06082_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_06083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_06084_, _06083_, _06082_);
  nand (_06085_, _06084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_06086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_06087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_06088_, _06087_, _06086_);
  and (_06089_, _06088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_06090_, _06089_);
  and (_06091_, _06090_, _06085_);
  and (_06092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_06093_, _06092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_06094_, _06093_);
  and (_06095_, _06094_, _06091_);
  and (_06096_, _06095_, _06081_);
  nor (_06097_, _06096_, _06071_);
  and (_06098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _05628_);
  not (_06099_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_06100_, _06084_, _06099_);
  not (_06101_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_06102_, _06088_, _06101_);
  nor (_06103_, _06102_, _06100_);
  not (_06104_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_06105_, _06092_, _06104_);
  not (_06106_, _06105_);
  not (_06107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_06109_, _06072_, _06107_);
  not (_06110_, _06109_);
  not (_06111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_06112_, _06075_, _06111_);
  not (_06113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_06114_, _06077_, _06113_);
  nor (_06115_, _06114_, _06112_);
  and (_06116_, _06115_, _06110_);
  and (_06117_, _06116_, _06106_);
  nand (_06118_, _06117_, _06103_);
  nand (_06119_, _06118_, _06098_);
  not (_06120_, _06119_);
  nor (_06121_, _06120_, _06097_);
  and (_06122_, _06121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not (_06123_, _06097_);
  nor (_06124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _05630_);
  and (_06125_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _05630_);
  nor (_06126_, _06125_, _06124_);
  nor (_06127_, _06126_, _06123_);
  or (_06128_, _06127_, _06122_);
  and (_06129_, _06128_, _06066_);
  and (_06130_, _06126_, _06065_);
  or (_06131_, _06130_, _06129_);
  and (_07816_, _06131_, _05141_);
  or (_06132_, _06081_, _06071_);
  nor (_06133_, _06119_, _06097_);
  not (_06134_, _06133_);
  or (_06135_, _06134_, _06116_);
  and (_06136_, _06135_, _06132_);
  nor (_06137_, _06065_, _05630_);
  not (_06138_, _06137_);
  or (_06139_, _06138_, _06136_);
  not (_06140_, _06103_);
  and (_06141_, _06140_, _06098_);
  and (_06142_, _06105_, _06098_);
  or (_06143_, _06142_, _06141_);
  or (_06144_, _06143_, _06097_);
  not (_06145_, _06095_);
  or (_06146_, _06132_, _06145_);
  and (_06147_, _06146_, _06137_);
  and (_06148_, _06147_, _06144_);
  or (_06150_, _06148_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_06151_, _06150_, _05141_);
  and (_07981_, _06151_, _06139_);
  nor (_06152_, _05277_, _05269_);
  and (_06153_, _05292_, _06152_);
  or (_06154_, _06153_, _05572_);
  and (_06155_, _06154_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nand (_06156_, _05301_, _06152_);
  and (_06157_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_06158_, _06157_, _06156_);
  nor (_06159_, _05446_, _05370_);
  not (_06160_, _06159_);
  or (_06161_, _05446_, _05381_);
  and (_06162_, _05538_, _06161_);
  or (_06163_, _06162_, _05425_);
  nand (_06164_, _06162_, _05425_);
  and (_06165_, _06164_, _05481_);
  nand (_06166_, _06165_, _06163_);
  or (_06167_, _05810_, _05808_);
  or (_06168_, _06167_, _05583_);
  or (_06169_, _05808_, _05516_);
  nand (_06170_, _05810_, _05501_);
  and (_06171_, _05809_, _05509_);
  and (_06172_, _05504_, _05446_);
  nor (_06173_, _06172_, _06171_);
  and (_06174_, _06173_, _06170_);
  and (_06175_, _06174_, _06169_);
  and (_06176_, _06175_, _06168_);
  and (_06177_, _06176_, _06166_);
  and (_06178_, _06177_, _06160_);
  not (_06179_, _06178_);
  and (_06180_, _05297_, _05291_);
  and (_06181_, _06180_, _06179_);
  or (_06182_, _06181_, _06158_);
  or (_06183_, _06182_, _06155_);
  and (_08821_, _06183_, _05141_);
  and (_06184_, _05649_, _05289_);
  and (_06185_, _06184_, _05647_);
  nand (_06186_, _06185_, _05963_);
  not (_06187_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_06188_, _05971_, _05638_);
  or (_06189_, _06188_, _06028_);
  and (_06190_, _06189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_06191_, _06190_, _06187_);
  or (_06192_, _06191_, _06185_);
  and (_06193_, _06192_, _05928_);
  and (_06194_, _06193_, _06186_);
  nor (_06195_, _06178_, _05928_);
  or (_06197_, _06195_, _06194_);
  and (_08859_, _06197_, _05141_);
  and (_09119_, _05141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nand (_06198_, _06119_, _05628_);
  or (_06199_, _06198_, _06097_);
  nand (_06200_, _06124_, _06065_);
  and (_06201_, _06200_, _05141_);
  and (_10115_, _06201_, _06199_);
  and (_06202_, _05266_, _05227_);
  and (_06203_, _05256_, _05173_);
  and (_06204_, _06010_, _06203_);
  and (_06205_, _06204_, _06202_);
  and (_06206_, _05274_, _05197_);
  and (_06207_, _06206_, _06007_);
  and (_06208_, _05922_, _06207_);
  nor (_06209_, _05186_, _05208_);
  nand (_06210_, _05197_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_06211_, _06210_, _06209_);
  or (_06212_, _06211_, _06208_);
  and (_06213_, _06212_, _06205_);
  nand (_06214_, _06205_, _05197_);
  and (_06215_, _06214_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_06216_, _06215_, _05927_);
  or (_06217_, _06216_, _06213_);
  nor (_06218_, _05724_, _05382_);
  nor (_06219_, _05715_, _05381_);
  or (_06220_, _06219_, _06218_);
  and (_06221_, _06220_, _05509_);
  or (_06222_, _05941_, _05716_);
  nand (_06223_, _06222_, _05943_);
  nand (_06224_, _05758_, _05937_);
  and (_06225_, _06224_, _05716_);
  or (_06226_, _06225_, _05938_);
  nand (_06227_, _06226_, _05381_);
  nand (_06228_, _06227_, _06223_);
  and (_06229_, _06228_, _05481_);
  nor (_06230_, _06229_, _06221_);
  nor (_06231_, _05715_, _05370_);
  not (_06233_, _06231_);
  and (_06234_, _05730_, _05485_);
  not (_06235_, _06234_);
  nor (_06236_, _05728_, _05516_);
  not (_06237_, _06236_);
  and (_06238_, _05727_, _05501_);
  and (_06239_, _05715_, _05504_);
  nor (_06240_, _06239_, _06238_);
  and (_06241_, _06240_, _06237_);
  and (_06242_, _06241_, _06235_);
  and (_06243_, _06242_, _06233_);
  and (_06244_, _06243_, _06230_);
  nand (_06245_, _06244_, _05927_);
  and (_06246_, _06245_, _05141_);
  and (_10153_, _06246_, _06217_);
  nor (_06247_, _06065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_06248_, _06247_);
  or (_06249_, _06248_, _06136_);
  and (_06250_, _06247_, _06146_);
  and (_06251_, _06250_, _06144_);
  or (_06253_, _06251_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_06254_, _06253_, _05141_);
  and (_10191_, _06254_, _06249_);
  and (_06255_, _06204_, _06009_);
  and (_06256_, _06255_, _06008_);
  nand (_06257_, _06256_, _05963_);
  or (_06259_, _06256_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_06260_, _05280_, _05256_);
  and (_06261_, _06260_, _05648_);
  and (_06262_, _06261_, _05926_);
  not (_06263_, _06262_);
  and (_06264_, _06263_, _06259_);
  and (_06265_, _06264_, _06257_);
  nor (_06266_, _06263_, _05960_);
  or (_06267_, _06266_, _06265_);
  and (_10239_, _06267_, _05141_);
  or (_06268_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_06269_, _06268_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor (_06270_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_06271_, _06270_, _05143_);
  and (_06272_, _06271_, _06269_);
  and (pc_log_change, _06272_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_06273_, _06004_, _05576_);
  not (_06274_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_06275_, _05576_, _05297_);
  nor (_06276_, _06275_, _06274_);
  or (_06277_, _06276_, _06273_);
  or (_06278_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_06279_, _06278_, _05141_);
  and (_12316_, _06279_, _06277_);
  and (_06280_, _05569_, _05297_);
  or (_06281_, _06280_, _05574_);
  and (_06282_, _06281_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  not (_06283_, _06244_);
  and (_06284_, _06275_, _06283_);
  or (_06285_, _06284_, _06282_);
  and (_12641_, _06285_, _05141_);
  and (_06286_, _06281_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_06287_, _06275_, _05522_);
  or (_06288_, _06287_, _06286_);
  and (_12994_, _06288_, _05141_);
  and (_06289_, _06281_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  not (_06290_, _06062_);
  and (_06291_, _06275_, _06290_);
  or (_06292_, _06291_, _06289_);
  and (_00302_, _06292_, _05141_);
  and (_06293_, _05141_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06295_, _06293_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_06296_, _06271_, _05141_);
  and (_06297_, _06269_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_06298_, _06297_, _06272_);
  not (_06299_, _06298_);
  not (_06300_, _06272_);
  not (_06301_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  not (_06302_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or (_06303_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or (_06304_, _06303_, _06302_);
  or (_06305_, _06304_, _06301_);
  not (_06306_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nand (_06307_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or (_06308_, _06307_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or (_06309_, _06308_, _06306_);
  and (_06310_, _06309_, _06305_);
  not (_06311_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  not (_06312_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_06313_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _06302_);
  nand (_06314_, _06313_, _06312_);
  or (_06315_, _06314_, _06311_);
  and (_06316_, _06315_, _06310_);
  not (_06317_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_06318_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_06319_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], _06318_);
  nand (_06320_, _06319_, _06302_);
  not (_06321_, _06320_);
  nand (_06322_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_06323_, _06322_, _06317_);
  not (_06324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_06325_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or (_06326_, _06325_, _06302_);
  or (_06327_, _06326_, _06324_);
  and (_06328_, _06325_, _06302_);
  nand (_06329_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_06330_, _06329_, _06327_);
  and (_06331_, _06330_, _06323_);
  nand (_06332_, _06331_, _06316_);
  or (_06333_, _06332_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_06334_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_06335_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _06334_);
  not (_06336_, _06335_);
  and (_06337_, _06336_, _06333_);
  or (_06338_, _06337_, _06300_);
  nand (_06339_, _06338_, _06299_);
  and (_06340_, _06269_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_06341_, _06340_, _06272_);
  not (_06342_, _06341_);
  not (_06343_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_06344_, _06308_, _06343_);
  nand (_06345_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_06346_, _06345_, _06344_);
  not (_06347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_06348_, _06326_, _06347_);
  nand (_06349_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_06350_, _06349_, _06348_);
  not (_06351_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_06352_, _06304_, _06351_);
  not (_06353_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_06354_, _06314_, _06353_);
  and (_06355_, _06354_, _06352_);
  and (_06356_, _06355_, _06350_);
  nand (_06357_, _06356_, _06346_);
  nand (_06358_, _06357_, _06317_);
  nand (_06360_, _06358_, _06334_);
  nor (_06361_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _06334_);
  not (_06362_, _06361_);
  and (_06363_, _06362_, _06360_);
  or (_06364_, _06363_, _06300_);
  nand (_06365_, _06364_, _06342_);
  and (_06366_, _06365_, _06339_);
  and (_06367_, _06269_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_06368_, _06367_, _06272_);
  not (_06369_, _06368_);
  not (_06370_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_06371_, _06314_, _06370_);
  nand (_06372_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_06373_, _06372_, _06371_);
  not (_06374_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_06375_, _06308_, _06374_);
  not (_06376_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_06377_, _06304_, _06376_);
  and (_06378_, _06377_, _06375_);
  not (_06379_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_06380_, _06326_, _06379_);
  nand (_06381_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_06382_, _06381_, _06380_);
  and (_06383_, _06382_, _06378_);
  nand (_06384_, _06383_, _06373_);
  nand (_06385_, _06384_, _06317_);
  nand (_06386_, _06385_, _06334_);
  nor (_06387_, _06334_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  not (_06388_, _06387_);
  and (_06389_, _06388_, _06386_);
  or (_06390_, _06389_, _06300_);
  and (_06391_, _06390_, _06369_);
  and (_06392_, _06269_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_06393_, _06392_, _06272_);
  not (_06394_, _06393_);
  not (_06395_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_06396_, _06308_, _06395_);
  nand (_06397_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_06398_, _06397_, _06396_);
  not (_06399_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_06400_, _06326_, _06399_);
  nand (_06401_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_06402_, _06401_, _06400_);
  not (_06403_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or (_06404_, _06304_, _06403_);
  not (_06406_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_06407_, _06314_, _06406_);
  and (_06408_, _06407_, _06404_);
  and (_06409_, _06408_, _06402_);
  and (_06410_, _06409_, _06398_);
  or (_06411_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_06412_, _06411_, _06410_);
  and (_06413_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  not (_06414_, _06413_);
  and (_06415_, _06414_, _06412_);
  nand (_06416_, _06415_, _06272_);
  and (_06417_, _06416_, _06394_);
  not (_06418_, _06417_);
  and (_06419_, _06418_, _06391_);
  and (_06420_, _06419_, _06366_);
  and (_06421_, _06269_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_06422_, _06421_, _06272_);
  not (_06423_, _06422_);
  not (_06425_, _06326_);
  and (_06426_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  not (_06427_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_06428_, _06304_, _06427_);
  not (_06429_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_06430_, _06308_, _06429_);
  nand (_06431_, _06430_, _06428_);
  nor (_06432_, _06431_, _06426_);
  nand (_06433_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not (_06434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_06436_, _06320_, _06434_);
  and (_06437_, _06436_, _06433_);
  not (_06438_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_06439_, _06314_, _06438_);
  and (_06440_, _06439_, _06317_);
  and (_06441_, _06440_, _06437_);
  nand (_06442_, _06441_, _06432_);
  or (_06444_, _06442_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_06445_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _06334_);
  not (_06446_, _06445_);
  and (_06447_, _06446_, _06444_);
  or (_06448_, _06447_, _06300_);
  and (_06449_, _06448_, _06423_);
  not (_06450_, _06449_);
  and (_06451_, _06269_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_06452_, _06451_, _06272_);
  not (_06453_, _06452_);
  nand (_06454_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_06455_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_06456_, _06455_, _06454_);
  not (_06457_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_06458_, _06326_, _06457_);
  not (_06459_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or (_06460_, _06304_, _06459_);
  and (_06461_, _06460_, _06458_);
  not (_06462_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_06463_, _06308_, _06462_);
  not (_06464_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_06465_, _06314_, _06464_);
  and (_06466_, _06465_, _06463_);
  and (_06467_, _06466_, _06461_);
  and (_06468_, _06467_, _06456_);
  or (_06469_, _06468_, _06411_);
  and (_06470_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  not (_06471_, _06470_);
  and (_06472_, _06471_, _06469_);
  nand (_06473_, _06472_, _06272_);
  and (_06474_, _06473_, _06453_);
  and (_06475_, _06269_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_06476_, _06475_, _06272_);
  not (_06477_, _06476_);
  nor (_06478_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_06479_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand (_06480_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_06481_, _06480_, _06479_);
  not (_06482_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_06483_, _06326_, _06482_);
  not (_06484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_06485_, _06308_, _06484_);
  and (_06486_, _06485_, _06483_);
  not (_06487_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or (_06488_, _06304_, _06487_);
  not (_06489_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_06490_, _06314_, _06489_);
  and (_06491_, _06490_, _06488_);
  and (_06492_, _06491_, _06486_);
  nand (_06493_, _06492_, _06481_);
  nand (_06494_, _06493_, _06478_);
  and (_06495_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  not (_06496_, _06495_);
  nand (_06497_, _06496_, _06494_);
  or (_06498_, _06497_, _06300_);
  and (_06499_, _06498_, _06477_);
  and (_06500_, _06269_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_06501_, _06500_, _06272_);
  not (_06502_, _06501_);
  nand (_06504_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_06505_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_06506_, _06505_, _06504_);
  not (_06508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_06509_, _06326_, _06508_);
  not (_06510_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_06511_, _06308_, _06510_);
  and (_06512_, _06511_, _06509_);
  not (_06514_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_06515_, _06304_, _06514_);
  not (_06516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_06517_, _06314_, _06516_);
  and (_06518_, _06517_, _06515_);
  and (_06519_, _06518_, _06512_);
  and (_06520_, _06519_, _06506_);
  or (_06521_, _06520_, _06411_);
  and (_06522_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  not (_06523_, _06522_);
  nand (_06524_, _06523_, _06521_);
  or (_06525_, _06524_, _06300_);
  and (_06526_, _06525_, _06502_);
  and (_06527_, _06526_, _06499_);
  and (_06528_, _06527_, _06474_);
  and (_06529_, _06528_, _06450_);
  and (_06530_, _06529_, _06420_);
  and (_06531_, _06364_, _06342_);
  and (_06532_, _06338_, _06299_);
  nand (_06533_, _06390_, _06369_);
  and (_06534_, _06533_, _06532_);
  and (_06535_, _06534_, _06418_);
  and (_06536_, _06535_, _06531_);
  nand (_06537_, _06498_, _06477_);
  nand (_06538_, _06525_, _06502_);
  and (_06539_, _06538_, _06537_);
  and (_06540_, _06539_, _06474_);
  and (_06541_, _06540_, _06536_);
  and (_06542_, _06541_, _06450_);
  or (_06543_, _06542_, _06530_);
  and (_06544_, _06535_, _06365_);
  and (_06545_, _06526_, _06537_);
  and (_06546_, _06545_, _06474_);
  and (_06547_, _06546_, _06450_);
  and (_06548_, _06547_, _06544_);
  and (_06549_, _06418_, _06533_);
  and (_06550_, _06549_, _06366_);
  not (_06551_, _06474_);
  and (_06552_, _06539_, _06551_);
  and (_06553_, _06552_, _06449_);
  and (_06554_, _06553_, _06550_);
  and (_06555_, _06538_, _06499_);
  and (_06556_, _06555_, _06551_);
  and (_06557_, _06556_, _06450_);
  and (_06558_, _06557_, _06550_);
  or (_06559_, _06558_, _06554_);
  and (_06560_, _06547_, _06536_);
  or (_06561_, _06560_, _06559_);
  or (_06562_, _06561_, _06548_);
  and (_06563_, _06545_, _06551_);
  and (_06564_, _06563_, _06449_);
  and (_06565_, _06563_, _06450_);
  and (_06566_, _06556_, _06449_);
  or (_06567_, _06566_, _06565_);
  or (_06568_, _06567_, _06564_);
  and (_06569_, _06568_, _06550_);
  and (_06570_, _06546_, _06449_);
  and (_06571_, _06570_, _06535_);
  and (_06572_, _06540_, _06450_);
  and (_06573_, _06550_, _06572_);
  and (_06574_, _06527_, _06551_);
  and (_06575_, _06574_, _06550_);
  or (_06576_, _06575_, _06573_);
  or (_06577_, _06576_, _06571_);
  or (_06578_, _06577_, _06569_);
  or (_06579_, _06578_, _06562_);
  or (_06580_, _06579_, _06543_);
  and (_06581_, _06580_, _06296_);
  or (_00855_, _06581_, _06295_);
  nor (_06582_, _05858_, _05856_);
  not (_06583_, _06582_);
  nor (_06584_, _05859_, _05845_);
  and (_06585_, _06584_, _06583_);
  not (_06586_, _06585_);
  nor (_06587_, _05827_, _05821_);
  nor (_06588_, _06587_, _05828_);
  nor (_06589_, _06588_, _05657_);
  not (_06590_, _06589_);
  not (_06591_, _05883_);
  nor (_06592_, _05887_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_06593_, _06592_, _05537_);
  nor (_06594_, _06593_, _05469_);
  and (_06595_, _05470_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_06596_, _06595_, _06594_);
  nor (_06597_, _06596_, _06591_);
  not (_06598_, _05355_);
  nor (_06599_, _05469_, _06598_);
  and (_06600_, _05354_, _05357_);
  and (_06601_, _06600_, ABINPUT000000[3]);
  nor (_06602_, _06601_, _06599_);
  not (_06603_, _05363_);
  or (_06604_, _05404_, _06603_);
  and (_06605_, _05537_, _05367_);
  and (_06606_, _05500_, _05349_);
  and (_06607_, _06606_, ABINPUT000[3]);
  nor (_06608_, _06607_, _06605_);
  and (_06610_, _06608_, _06604_);
  and (_06611_, _06610_, _06602_);
  and (_06612_, _06611_, _05557_);
  not (_06613_, _06612_);
  nor (_06614_, _06613_, _06597_);
  and (_06615_, _06614_, _05545_);
  and (_06616_, _06615_, _06590_);
  and (_06617_, _06616_, _06586_);
  and (_06618_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05143_);
  and (_06619_, _06618_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_06620_, _06206_, _05186_);
  and (_06621_, _06018_, _05649_);
  and (_06622_, _06621_, _06620_);
  nor (_06623_, _06622_, _06619_);
  not (_06624_, _06623_);
  nand (_06625_, _06624_, _06617_);
  or (_06626_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_06627_, _06626_, _05141_);
  and (_01188_, _06627_, _06625_);
  nor (_06628_, _05715_, _06598_);
  or (_06629_, _05678_, _06603_);
  nand (_06630_, _06230_, _06629_);
  not (_06631_, _05367_);
  nor (_06632_, _05758_, _06631_);
  or (_06633_, _06236_, _06234_);
  or (_06634_, _06633_, _06632_);
  or (_06635_, _06634_, _06630_);
  not (_06636_, _05885_);
  and (_06637_, _05887_, _05883_);
  nor (_06638_, _06637_, _05381_);
  and (_06639_, _06638_, _06636_);
  not (_06640_, _06639_);
  and (_06641_, _06637_, _05373_);
  and (_06642_, _06641_, _05759_);
  nor (_06643_, _06642_, _05716_);
  nor (_06644_, _06643_, _06640_);
  nor (_06645_, _06641_, _05759_);
  nor (_06646_, _06639_, _06645_);
  and (_06647_, _06646_, _05716_);
  not (_06648_, _05884_);
  nor (_06649_, _06641_, _06648_);
  and (_06650_, _06640_, _06649_);
  or (_06651_, _06650_, _06647_);
  nor (_06652_, _06651_, _06644_);
  nor (_06653_, _06652_, _06591_);
  and (_06654_, _06600_, ABINPUT000000[7]);
  nor (_06655_, _06654_, _06653_);
  nand (_06656_, _06655_, _06240_);
  and (_06657_, _05876_, _05870_);
  not (_06658_, _06657_);
  and (_06659_, _05877_, _05844_);
  and (_06660_, _06659_, _06658_);
  and (_06661_, _05838_, _05782_);
  nor (_06662_, _06661_, _05839_);
  nor (_06663_, _06662_, _05657_);
  and (_06664_, _06606_, ABINPUT000[7]);
  or (_06665_, _06664_, _06663_);
  or (_06666_, _06665_, _06660_);
  or (_06667_, _06666_, _06656_);
  or (_06668_, _06667_, _06635_);
  or (_06669_, _06668_, _06628_);
  or (_06670_, _06669_, _06623_);
  or (_06671_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_06672_, _06671_, _05141_);
  and (_01207_, _06672_, _06670_);
  or (_06674_, _05572_, _05279_);
  and (_06675_, _06674_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nand (_06676_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_06677_, _06676_, _05278_);
  and (_06678_, _05297_, _05269_);
  and (_06679_, _06678_, _06179_);
  or (_06680_, _06679_, _06677_);
  or (_06681_, _06680_, _06675_);
  and (_02780_, _06681_, _05141_);
  not (_06682_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_06683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nor (_06684_, _06683_, _06682_);
  and (_06685_, _06684_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_06686_, _06685_);
  and (_06687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_06688_, _06687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor (_06689_, _06688_, _06686_);
  not (_06690_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not (_06691_, _06683_);
  and (_06692_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_06693_, _06692_, _06691_);
  nor (_06694_, _06693_, _06685_);
  or (_06695_, _06694_, _06690_);
  or (_06696_, _06695_, _06689_);
  and (_06697_, _06685_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_06698_, _06697_, _06687_);
  or (_06699_, _06698_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_06700_, _06699_, _05141_);
  and (_03603_, _06700_, _06696_);
  not (_06701_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_06702_, _06678_, _06701_);
  not (_06703_, _05604_);
  and (_06705_, _06678_, _06703_);
  or (_06706_, _06705_, _06702_);
  and (_03622_, _06706_, _05141_);
  and (_06707_, _05297_, _05273_);
  not (_06708_, _06707_);
  or (_06709_, _06708_, _06004_);
  or (_06710_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_06711_, _06710_, _05141_);
  and (_03936_, _06711_, _06709_);
  nor (_06713_, rst, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_06714_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_06715_, _05141_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_06716_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_04037_, _06716_, _06714_);
  and (_06718_, _05522_, _05277_);
  not (_06719_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_06720_, _05277_, _06719_);
  or (_06721_, _06720_, _05572_);
  or (_06722_, _06721_, _06718_);
  or (_06723_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_06724_, _06723_, _05141_);
  and (_04141_, _06724_, _06722_);
  and (_06725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_06726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_06727_, _06726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_06728_, _06727_, _06725_);
  or (_06729_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  not (_06730_, _06728_);
  or (_06731_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_06732_, _06731_, _06729_);
  and (_06733_, _05241_, _05228_);
  and (_06734_, _06733_, _05267_);
  not (_06735_, _05925_);
  nor (_06736_, _06735_, _05172_);
  and (_06737_, _06736_, _06620_);
  and (_06738_, _06737_, _06734_);
  or (_06739_, _06738_, _06732_);
  nand (_06740_, _06738_, _06178_);
  and (_06741_, _06740_, _06739_);
  and (_06742_, _06033_, _05925_);
  and (_06743_, _06742_, _06734_);
  or (_06744_, _06743_, _06741_);
  not (_06745_, _06743_);
  or (_06746_, _06745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_06747_, _06746_, _05141_);
  and (_05132_, _06747_, _06744_);
  or (_06748_, _06708_, _05522_);
  or (_06749_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_06750_, _06749_, _05141_);
  and (_05139_, _06750_, _06748_);
  nand (_06751_, _06678_, _05560_);
  or (_06752_, _06678_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_06753_, _06752_, _05141_);
  and (_05140_, _06753_, _06751_);
  and (_06754_, _06293_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_06755_, _06419_, _06339_);
  and (_06756_, _06755_, _06553_);
  and (_06757_, _06552_, _06450_);
  and (_06758_, _06757_, _06420_);
  and (_06759_, _06531_, _06339_);
  and (_06760_, _06759_, _06419_);
  or (_06761_, _06757_, _06570_);
  and (_06762_, _06761_, _06760_);
  or (_06763_, _06762_, _06758_);
  or (_06764_, _06763_, _06756_);
  and (_06765_, _06540_, _06449_);
  and (_06766_, _06555_, _06474_);
  and (_06767_, _06766_, _06449_);
  or (_06768_, _06767_, _06765_);
  and (_06769_, _06768_, _06420_);
  and (_06770_, _06391_, _06532_);
  and (_06771_, _06770_, _06418_);
  and (_06772_, _06771_, _06552_);
  or (_06773_, _06770_, _06417_);
  and (_06774_, _06773_, _06767_);
  or (_06775_, _06774_, _06772_);
  or (_06776_, _06775_, _06769_);
  and (_06777_, _06761_, _06417_);
  and (_06778_, _06449_, _06417_);
  and (_06779_, _06778_, _06552_);
  or (_06780_, _06779_, _06777_);
  and (_06781_, _06550_, _06765_);
  and (_06782_, _06766_, _06450_);
  and (_06784_, _06782_, _06536_);
  or (_06785_, _06784_, _06781_);
  or (_06786_, _06785_, _06780_);
  or (_06787_, _06786_, _06776_);
  or (_06788_, _06787_, _06764_);
  and (_06789_, _06788_, _06296_);
  or (_05235_, _06789_, _06754_);
  not (_06790_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_06791_, \oc8051_top_1.oc8051_decoder1.state [0], _05143_);
  and (_06792_, _06791_, _06790_);
  and (_06793_, _06782_, _06420_);
  and (_06795_, _06572_, _06420_);
  nor (_06796_, _06795_, _06793_);
  not (_06797_, _06796_);
  and (_06798_, _06797_, _06792_);
  and (_06799_, _06760_, _06572_);
  and (_06800_, _06799_, _06270_);
  or (_06801_, _06800_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_06802_, _06801_, _06798_);
  or (_06803_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05143_);
  and (_06804_, _06803_, _05141_);
  and (_05238_, _06804_, _06802_);
  not (_06805_, _06541_);
  and (_06806_, _06550_, _06529_);
  nor (_06807_, _06449_, _06417_);
  and (_06808_, _06807_, _06534_);
  and (_06809_, _06808_, _06528_);
  nor (_06810_, _06809_, _06806_);
  and (_06811_, _06810_, _06805_);
  not (_06812_, _06811_);
  and (_06813_, _06812_, _06792_);
  or (_06814_, _06813_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_06815_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_06816_, _06759_, _06549_);
  and (_06818_, _06816_, _06449_);
  and (_06819_, _06553_, _06544_);
  or (_06820_, _06819_, _06818_);
  or (_06821_, _06270_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06822_, _06821_, _06542_);
  or (_06823_, _06822_, _06820_);
  and (_06824_, _06823_, _06815_);
  or (_06825_, _06824_, _06814_);
  or (_06826_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05143_);
  and (_06827_, _06826_, _05141_);
  and (_05251_, _06827_, _06825_);
  and (_06828_, _06528_, _06449_);
  nand (_06829_, _06828_, _06550_);
  and (_06830_, _06829_, _06811_);
  not (_06831_, _06296_);
  and (_06832_, _06535_, _06528_);
  or (_06833_, _06832_, _06831_);
  or (_05304_, _06833_, _06830_);
  not (_06834_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_06835_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05143_);
  and (_06836_, _06835_, _06834_);
  not (_06837_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_06838_, _06618_, _06837_);
  and (_06839_, _06733_, _06260_);
  and (_06840_, _06839_, _05272_);
  and (_06841_, _06840_, _05925_);
  nor (_06842_, _06841_, _06838_);
  not (_06843_, _05691_);
  and (_06844_, _05840_, _06843_);
  nor (_06845_, _05840_, _06843_);
  nor (_06846_, _06845_, _06844_);
  and (_06847_, _06846_, _05656_);
  not (_06848_, _06847_);
  nor (_06849_, _05879_, _06843_);
  and (_06850_, _05879_, _06843_);
  nor (_06851_, _06850_, _06849_);
  and (_06852_, _06851_, _05844_);
  nor (_06853_, _06639_, _06649_);
  and (_06854_, _06853_, _05678_);
  nor (_06855_, _06853_, _05678_);
  or (_06856_, _06855_, _06854_);
  and (_06857_, _06856_, _05883_);
  nor (_06858_, _05715_, _06631_);
  and (_06859_, _05535_, _05909_);
  and (_06860_, _05381_, _05907_);
  and (_06861_, _06600_, ABINPUT000000[8]);
  or (_06862_, _06861_, _06860_);
  or (_06863_, _06862_, _06859_);
  nor (_06864_, _06863_, _06858_);
  nor (_06865_, _05678_, _06598_);
  and (_06866_, _06606_, ABINPUT000[8]);
  nor (_06867_, _06866_, _06865_);
  and (_06868_, _06867_, _05956_);
  and (_06869_, _06868_, _06864_);
  not (_06870_, _06869_);
  nor (_06871_, _06870_, _06857_);
  and (_06872_, _06871_, _05949_);
  not (_06873_, _06872_);
  nor (_06874_, _06873_, _06852_);
  and (_06875_, _06874_, _06848_);
  nor (_06876_, _06875_, _06842_);
  and (_06877_, _05241_, _05172_);
  and (_06878_, _06877_, _05256_);
  nor (_06879_, _05266_, _05227_);
  and (_06880_, _06879_, _05647_);
  and (_06881_, _06880_, _06878_);
  and (_06882_, _06881_, _06008_);
  and (_06883_, _06882_, _05963_);
  not (_06884_, _06842_);
  nor (_06885_, _06882_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_06886_, _06885_, _06884_);
  nor (_06888_, _06886_, _06883_);
  nor (_06889_, _06888_, _06876_);
  or (_06890_, _06889_, _06836_);
  nor (_06891_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_06892_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05663_);
  nor (_06893_, _06892_, _06891_);
  nor (_06894_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_06895_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05699_);
  nor (_06896_, _06895_, _06894_);
  not (_06897_, _06896_);
  nor (_06898_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_06899_, _05390_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_06900_, _06899_, _06898_);
  nand (_06901_, _05880_, _05846_);
  nor (_06902_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_06904_, _05411_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_06905_, _06904_, _06902_);
  and (_06906_, _06905_, _06901_);
  nor (_06907_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_06908_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05436_);
  nor (_06909_, _06908_, _06907_);
  and (_06910_, _06909_, _06906_);
  nor (_06911_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_06912_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05455_);
  nor (_06913_, _06912_, _06911_);
  and (_06914_, _06913_, _06910_);
  and (_06915_, _06914_, _06900_);
  nor (_06916_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_06917_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05739_);
  nor (_06918_, _06917_, _06916_);
  nor (_06919_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_06920_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05317_);
  nor (_06921_, _06920_, _06919_);
  and (_06922_, _06921_, _06918_);
  nand (_06923_, _06922_, _06915_);
  or (_06924_, _06923_, _06897_);
  nor (_06925_, _06924_, _06893_);
  and (_06926_, _06924_, _06893_);
  or (_06927_, _06926_, _06925_);
  and (_06928_, _06927_, _05844_);
  and (_06929_, _05768_, _05382_);
  not (_06930_, _06929_);
  nand (_06931_, _05495_, _05382_);
  nor (_06932_, _05942_, _05678_);
  and (_06933_, _06932_, _05584_);
  and (_06934_, _06933_, _05809_);
  and (_06935_, _06934_, _05799_);
  and (_06936_, _06935_, _05830_);
  or (_06937_, _06936_, _05381_);
  and (_06938_, _06937_, _06931_);
  and (_06939_, _06938_, _06930_);
  and (_06940_, _05678_, _05581_);
  and (_06941_, _06940_, _05938_);
  and (_06942_, _06941_, _05807_);
  and (_06943_, _06942_, _05532_);
  and (_06944_, _06943_, _05795_);
  and (_06945_, _06944_, _05495_);
  and (_06946_, _06945_, _05768_);
  nor (_06947_, _06946_, _05382_);
  not (_06948_, _06947_);
  and (_06949_, _06948_, _06939_);
  and (_06950_, _05724_, _05382_);
  nor (_06951_, _06950_, _06218_);
  and (_06952_, _06951_, _06949_);
  or (_06953_, _06952_, _05685_);
  nand (_06954_, _06952_, _05685_);
  and (_06955_, _06954_, _06953_);
  and (_06956_, _06955_, _05481_);
  nor (_06958_, _05678_, _05382_);
  nor (_06959_, _05684_, _05381_);
  or (_06961_, _06959_, _06958_);
  and (_06963_, _06961_, _05509_);
  nor (_06964_, _05404_, _05893_);
  nor (_06965_, _05684_, _06598_);
  and (_06967_, _06600_, ABINPUT000000[16]);
  and (_06968_, _06606_, ABINPUT000[16]);
  or (_06969_, _06968_, _06967_);
  or (_06970_, _06969_, _06965_);
  or (_06972_, _06970_, _06964_);
  or (_06973_, _06972_, _06963_);
  or (_06974_, _06973_, _06956_);
  or (_06975_, _06974_, _06928_);
  nand (_06976_, _06975_, _06836_);
  nand (_06977_, _06976_, _06890_);
  and (_05329_, _06977_, _05141_);
  and (_06978_, _06293_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_06979_, _06771_, _06546_);
  and (_06980_, _06979_, _06450_);
  and (_06981_, _06760_, _06570_);
  and (_06982_, _06772_, _06449_);
  or (_06983_, _06982_, _06981_);
  or (_06985_, _06983_, _06980_);
  or (_06986_, _06756_, _06571_);
  or (_06987_, _06986_, _06784_);
  and (_06988_, _06778_, _06546_);
  or (_06989_, _06988_, _06779_);
  and (_06990_, _06782_, _06544_);
  or (_06992_, _06990_, _06989_);
  and (_06993_, _06767_, _06544_);
  and (_06994_, _06760_, _06547_);
  and (_06995_, _06450_, _06417_);
  and (_06996_, _06995_, _06545_);
  and (_06997_, _06996_, _06474_);
  or (_06998_, _06997_, _06994_);
  or (_06999_, _06998_, _06993_);
  or (_07000_, _06999_, _06992_);
  or (_07001_, _07000_, _06987_);
  or (_07002_, _07001_, _06985_);
  and (_07003_, _07002_, _06296_);
  or (_05340_, _07003_, _06978_);
  and (_07004_, _06269_, _05143_);
  and (_07005_, _07004_, _06815_);
  not (_07006_, _06497_);
  nor (_07007_, _06524_, _06472_);
  and (_07008_, _07007_, _07006_);
  not (_07009_, _06415_);
  nor (_07010_, _07009_, _06389_);
  and (_07011_, _07010_, _06337_);
  and (_07012_, _07011_, _06363_);
  and (_07013_, _07012_, _07008_);
  not (_07014_, _06472_);
  nor (_07015_, _06524_, _07014_);
  and (_07016_, _07015_, _06497_);
  not (_07017_, _06363_);
  and (_07018_, _07011_, _07017_);
  and (_07019_, _07018_, _07016_);
  nor (_07020_, _07009_, _06337_);
  and (_07021_, _07020_, _06389_);
  and (_07022_, _07021_, _07017_);
  not (_07023_, _06447_);
  and (_07025_, _07007_, _07023_);
  and (_07026_, _07025_, _07022_);
  or (_07028_, _07026_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_07029_, _07028_, _07019_);
  or (_07030_, _07029_, _07013_);
  and (_07031_, _07030_, _07005_);
  nor (_07032_, _07004_, _06815_);
  or (_07033_, _07032_, rst);
  or (_05369_, _07033_, _07031_);
  nor (_07034_, _06993_, _06548_);
  and (_07035_, _06760_, _06553_);
  or (_07036_, _06981_, _07035_);
  and (_07037_, _06565_, _06535_);
  nor (_07039_, _07037_, _07036_);
  nand (_07040_, _07039_, _07034_);
  and (_07041_, _06527_, _06449_);
  and (_07042_, _07041_, _06760_);
  or (_07043_, _07042_, _06799_);
  and (_07044_, _06550_, _06546_);
  or (_07045_, _07044_, _07043_);
  or (_07046_, _07045_, _06819_);
  and (_07047_, _06544_, _06765_);
  or (_07048_, _07047_, _06994_);
  nand (_07049_, _06535_, _06365_);
  not (_07050_, _06570_);
  or (_07051_, _07050_, _07049_);
  nand (_07052_, _06757_, _06760_);
  and (_07053_, _06574_, _06450_);
  nand (_07054_, _07053_, _06535_);
  and (_07055_, _07054_, _07052_);
  nand (_07056_, _07055_, _07051_);
  or (_07057_, _07056_, _07048_);
  or (_07058_, _07057_, _07046_);
  or (_07059_, _07058_, _07040_);
  or (_07060_, _06997_, _06979_);
  and (_07062_, _06778_, _06527_);
  and (_07063_, _06995_, _06766_);
  or (_07064_, _07063_, _07062_);
  or (_07065_, _07064_, _07060_);
  or (_07066_, _07065_, _06780_);
  and (_07067_, _06782_, _06771_);
  and (_07068_, _06449_, _06418_);
  and (_07069_, _07068_, _06770_);
  and (_07070_, _07069_, _06527_);
  or (_07071_, _07070_, _06772_);
  or (_07072_, _07071_, _07067_);
  and (_07073_, _06564_, _06535_);
  and (_07074_, _06807_, _06770_);
  and (_07076_, _07074_, _06540_);
  or (_07077_, _07076_, _07073_);
  and (_07078_, _06995_, _06540_);
  or (_07079_, _07078_, _06818_);
  or (_07080_, _07079_, _07077_);
  or (_07081_, _07080_, _07072_);
  or (_07083_, _07081_, _07066_);
  or (_07084_, _07083_, _07059_);
  and (_07085_, _07084_, _06271_);
  and (_07086_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.wr );
  and (_07087_, \oc8051_top_1.oc8051_decoder1.state [1], _05143_);
  and (_07088_, _07087_, _06815_);
  and (_07089_, _07088_, _06820_);
  or (_07090_, _07089_, _06798_);
  and (_07091_, _07088_, _06554_);
  or (_07092_, _07091_, _07090_);
  or (_07093_, _07092_, _07086_);
  or (_07094_, _07093_, _07085_);
  and (_05451_, _07094_, _05141_);
  not (_07096_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor (_07097_, _05291_, _07096_);
  and (_07099_, _06004_, _05291_);
  or (_07100_, _07099_, _05572_);
  or (_07101_, _07100_, _07097_);
  or (_07102_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_07103_, _07102_, _05141_);
  and (_05468_, _07103_, _07101_);
  or (_07104_, _06556_, _06765_);
  and (_07105_, _06755_, _06556_);
  or (_07106_, _07105_, _06773_);
  and (_07107_, _07106_, _07104_);
  and (_07108_, _06765_, _06420_);
  and (_07109_, _06760_, _06765_);
  or (_07110_, _07109_, _07108_);
  or (_07111_, _07110_, _07107_);
  and (_07112_, _07111_, _06271_);
  and (_07113_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_07114_, _06796_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_07115_, _07114_, _07113_);
  or (_07116_, _07115_, _07112_);
  and (_05502_, _07116_, _05141_);
  not (_07117_, _06270_);
  or (_07118_, _06337_, _07117_);
  or (_07119_, _06270_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_07120_, _07119_, _05141_);
  and (_05558_, _07120_, _07118_);
  nor (_05596_, _06472_, rst);
  nor (_07121_, _06271_, _05660_);
  nor (_07123_, _06308_, _06459_);
  nor (_07124_, _06314_, _06462_);
  nor (_07125_, _07124_, _07123_);
  and (_07126_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_07127_, _06320_, _06464_);
  nor (_07128_, _07127_, _07126_);
  and (_07129_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_07130_, _06304_, _06457_);
  nor (_07131_, _07130_, _07129_);
  and (_07132_, _07131_, _07128_);
  and (_07133_, _07132_, _07125_);
  and (_07134_, _06271_, _06317_);
  not (_07135_, _07134_);
  nor (_07136_, _07135_, _07133_);
  nor (_07137_, _07136_, _07121_);
  nor (_05599_, _07137_, rst);
  not (_07138_, _06619_);
  not (_07139_, _06918_);
  nand (_07140_, _06921_, _06915_);
  nand (_07141_, _07140_, _07139_);
  or (_07142_, _07140_, _07139_);
  and (_07143_, _07142_, _05844_);
  and (_07144_, _07143_, _07141_);
  nor (_07145_, _06945_, _05382_);
  not (_07146_, _07145_);
  and (_07147_, _07146_, _06938_);
  and (_07148_, _07147_, _05768_);
  nor (_07149_, _07147_, _05768_);
  or (_07150_, _07149_, _07148_);
  and (_07151_, _07150_, _05481_);
  nand (_07152_, _05758_, _05381_);
  nor (_07153_, _06929_, _05510_);
  and (_07154_, _07153_, _07152_);
  and (_07155_, _05537_, _05892_);
  nor (_07156_, _05768_, _06598_);
  and (_07157_, _06600_, ABINPUT000000[14]);
  and (_07158_, _06606_, ABINPUT000[14]);
  or (_07159_, _07158_, _07157_);
  or (_07161_, _07159_, _07156_);
  or (_07162_, _07161_, _07155_);
  or (_07163_, _07162_, _07154_);
  or (_07164_, _07163_, _07151_);
  or (_07166_, _07164_, _07144_);
  or (_07167_, _07166_, _07138_);
  and (_07168_, _06621_, _06032_);
  not (_07169_, _07168_);
  nor (_07170_, _05836_, _05786_);
  nor (_07171_, _07170_, _05837_);
  nor (_07172_, _07171_, _05657_);
  not (_07173_, _07172_);
  and (_07174_, _05869_, _05865_);
  not (_07175_, _07174_);
  and (_07176_, _05870_, _05844_);
  and (_07177_, _07176_, _07175_);
  nor (_07178_, _06642_, _06645_);
  nor (_07179_, _07178_, _06640_);
  and (_07180_, _07178_, _06640_);
  or (_07181_, _07180_, _06591_);
  nor (_07182_, _07181_, _07179_);
  nor (_07183_, _06631_, _05346_);
  and (_07184_, _06600_, ABINPUT000000[6]);
  and (_07185_, _06606_, ABINPUT000[6]);
  nor (_07186_, _07185_, _07184_);
  not (_07187_, _07186_);
  nor (_07188_, _07187_, _07183_);
  nor (_07189_, _05758_, _06598_);
  not (_07190_, _07189_);
  or (_07191_, _05715_, _06603_);
  and (_07192_, _07191_, _07190_);
  and (_07193_, _07192_, _07188_);
  and (_07194_, _07193_, _06002_);
  not (_07195_, _07194_);
  nor (_07196_, _07195_, _07182_);
  and (_07197_, _07196_, _05991_);
  not (_07198_, _07197_);
  nor (_07199_, _07198_, _07177_);
  and (_07200_, _07199_, _07173_);
  nor (_07201_, _07200_, _07169_);
  and (_07202_, _07169_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_07203_, _07202_, _06619_);
  or (_07204_, _07203_, _07201_);
  and (_07205_, _07204_, _05141_);
  and (_05687_, _07205_, _07167_);
  or (_07207_, _06921_, _06915_);
  and (_07208_, _07140_, _05844_);
  and (_07209_, _07208_, _07207_);
  nor (_07210_, _06944_, _05382_);
  not (_07211_, _07210_);
  and (_07212_, _07211_, _06937_);
  nand (_07213_, _07212_, _05771_);
  or (_07214_, _07212_, _05771_);
  and (_07215_, _07214_, _07213_);
  and (_07216_, _07215_, _05481_);
  nand (_07217_, _05381_, _05346_);
  and (_07218_, _06931_, _05509_);
  and (_07219_, _07218_, _07217_);
  and (_07220_, _05535_, _05892_);
  nor (_07221_, _05495_, _06598_);
  and (_07222_, _06600_, ABINPUT000000[13]);
  and (_07223_, _06606_, ABINPUT000[13]);
  or (_07224_, _07223_, _07222_);
  or (_07225_, _07224_, _07221_);
  or (_07226_, _07225_, _07220_);
  or (_07227_, _07226_, _07219_);
  or (_07228_, _07227_, _07216_);
  or (_07229_, _07228_, _07209_);
  or (_07230_, _07229_, _07138_);
  nor (_07231_, _05835_, _05498_);
  and (_07232_, _05835_, _05498_);
  nor (_07233_, _07232_, _07231_);
  and (_07234_, _07233_, _05656_);
  not (_07235_, _07234_);
  nor (_07236_, _05864_, _05498_);
  nor (_07237_, _07236_, _05845_);
  and (_07238_, _07237_, _05865_);
  nor (_07239_, _05887_, _06591_);
  nor (_07240_, _07239_, _05355_);
  nor (_07241_, _07240_, _05346_);
  not (_07242_, _07241_);
  and (_07243_, _06637_, _05346_);
  or (_07244_, _05758_, _06603_);
  nor (_07245_, _05404_, _06631_);
  and (_07246_, _06600_, ABINPUT000000[5]);
  and (_07248_, _06606_, ABINPUT000[5]);
  nor (_07249_, _07248_, _07246_);
  not (_07250_, _07249_);
  nor (_07251_, _07250_, _07245_);
  and (_07252_, _07251_, _07244_);
  not (_07253_, _07252_);
  nor (_07254_, _07253_, _07243_);
  and (_07255_, _07254_, _07242_);
  and (_07256_, _07255_, _05521_);
  not (_07257_, _07256_);
  nor (_07258_, _07257_, _07238_);
  and (_07259_, _07258_, _07235_);
  nor (_07260_, _07259_, _07169_);
  and (_07261_, _07169_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_07262_, _07261_, _06619_);
  or (_07263_, _07262_, _07260_);
  and (_07264_, _07263_, _05141_);
  and (_05690_, _07264_, _07230_);
  or (_07265_, _06923_, _06896_);
  nand (_07266_, _06923_, _06896_);
  nand (_07267_, _07266_, _07265_);
  nand (_07268_, _07267_, _05844_);
  and (_07269_, _06949_, _05724_);
  nor (_07270_, _06949_, _05724_);
  nor (_07271_, _07270_, _07269_);
  nor (_07272_, _07271_, _05597_);
  and (_07273_, _06606_, ABINPUT000[15]);
  and (_07274_, _05715_, _05381_);
  not (_07275_, _07274_);
  nor (_07276_, _06950_, _05510_);
  and (_07278_, _07276_, _07275_);
  nor (_07279_, _05469_, _05893_);
  nor (_07280_, _05724_, _06598_);
  and (_07281_, _06600_, ABINPUT000000[15]);
  or (_07282_, _07281_, _07280_);
  or (_07283_, _07282_, _07279_);
  or (_07284_, _07283_, _07278_);
  nor (_07285_, _07284_, _07273_);
  not (_07286_, _07285_);
  nor (_07287_, _07286_, _07272_);
  nand (_07288_, _07287_, _07268_);
  or (_07289_, _07288_, _07138_);
  and (_07290_, _07168_, _06669_);
  and (_07291_, _07169_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_07292_, _07291_, _06619_);
  or (_07293_, _07292_, _07290_);
  and (_07294_, _07293_, _05141_);
  and (_05698_, _07294_, _07289_);
  or (_07295_, _06914_, _06900_);
  nor (_07296_, _06915_, _05845_);
  nand (_07298_, _07296_, _07295_);
  not (_07299_, _05894_);
  or (_07300_, _06935_, _05381_);
  nor (_07301_, _06943_, _05382_);
  not (_07302_, _07301_);
  and (_07303_, _07302_, _07300_);
  nor (_07304_, _07303_, _05830_);
  and (_07305_, _07303_, _05830_);
  or (_07306_, _07305_, _05597_);
  nor (_07307_, _07306_, _07304_);
  nor (_07308_, _05510_, _05404_);
  not (_07309_, _07308_);
  nor (_07310_, _05795_, _06598_);
  and (_07311_, _06600_, ABINPUT000000[12]);
  and (_07312_, _06606_, ABINPUT000[12]);
  nor (_07313_, _07312_, _07311_);
  not (_07314_, _07313_);
  nor (_07315_, _07314_, _07310_);
  nand (_07316_, _07315_, _07309_);
  nor (_07317_, _07316_, _07307_);
  and (_07318_, _07317_, _07299_);
  nand (_07319_, _07318_, _07298_);
  or (_07320_, _07319_, _07138_);
  nor (_07321_, _05828_, _05819_);
  nor (_07322_, _07321_, _05829_);
  nor (_07323_, _07322_, _05657_);
  not (_07324_, _07323_);
  nor (_07325_, _05859_, _05854_);
  or (_07326_, _07325_, _05845_);
  nor (_07327_, _07326_, _05860_);
  not (_07328_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_07329_, _05470_, _07328_);
  nor (_07330_, _07329_, _05405_);
  not (_07331_, _07330_);
  and (_07332_, _07331_, _07239_);
  nor (_07333_, _05404_, _06598_);
  and (_07334_, _06600_, ABINPUT000000[4]);
  and (_07335_, _06606_, ABINPUT000[4]);
  nor (_07336_, _07335_, _07334_);
  not (_07337_, _07336_);
  nor (_07338_, _07337_, _07333_);
  or (_07339_, _06603_, _05346_);
  nor (_07340_, _05469_, _06631_);
  not (_07341_, _07340_);
  and (_07342_, _07341_, _07339_);
  and (_07343_, _07342_, _07338_);
  not (_07344_, _07343_);
  nor (_07345_, _07344_, _07332_);
  and (_07346_, _07345_, _06060_);
  and (_07347_, _07346_, _06048_);
  not (_07348_, _07347_);
  nor (_07349_, _07348_, _07327_);
  and (_07350_, _07349_, _07324_);
  nand (_07351_, _07350_, _07168_);
  or (_07352_, _07168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_07353_, _07352_, _07351_);
  or (_07354_, _07353_, _06619_);
  and (_07355_, _07354_, _05141_);
  and (_05707_, _07355_, _07320_);
  or (_07356_, _06913_, _06910_);
  nor (_07357_, _06914_, _05845_);
  nand (_07358_, _07357_, _07356_);
  or (_07359_, _06934_, _05381_);
  nor (_07360_, _06942_, _05382_);
  not (_07361_, _07360_);
  and (_07362_, _07361_, _07359_);
  and (_07363_, _07362_, _05799_);
  nor (_07364_, _07362_, _05799_);
  nor (_07365_, _07364_, _07363_);
  and (_07366_, _07365_, _05481_);
  nor (_07367_, _05715_, _05893_);
  nor (_07368_, _05532_, _06598_);
  and (_07369_, _06600_, ABINPUT000000[11]);
  or (_07370_, _07369_, _07368_);
  nor (_07371_, _07370_, _07367_);
  nor (_07372_, _05510_, _05469_);
  and (_07373_, _06606_, ABINPUT000[11]);
  nor (_07374_, _07373_, _07372_);
  and (_07375_, _07374_, _07371_);
  not (_07376_, _07375_);
  nor (_07377_, _07376_, _07366_);
  nand (_07378_, _07377_, _07358_);
  or (_07379_, _07378_, _07138_);
  or (_07380_, _07168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nand (_07381_, _07168_, _06617_);
  and (_07382_, _07381_, _07380_);
  or (_07383_, _07382_, _06619_);
  and (_07384_, _07383_, _05141_);
  and (_05714_, _07384_, _07379_);
  or (_07385_, _06909_, _06906_);
  nor (_07386_, _06910_, _05845_);
  nand (_07387_, _07386_, _07385_);
  nor (_07388_, _06933_, _05381_);
  nor (_07389_, _06941_, _05382_);
  nor (_07390_, _07389_, _07388_);
  and (_07391_, _07390_, _05807_);
  nor (_07392_, _07390_, _05807_);
  or (_07393_, _07392_, _07391_);
  and (_07394_, _07393_, _05481_);
  nor (_07395_, _05758_, _05893_);
  and (_07396_, _05809_, _05355_);
  and (_07397_, _06600_, ABINPUT000000[10]);
  or (_07398_, _07397_, _07396_);
  nor (_07399_, _07398_, _07395_);
  and (_07400_, _05509_, _05537_);
  and (_07401_, _06606_, ABINPUT000[10]);
  nor (_07402_, _07401_, _07400_);
  and (_07403_, _07402_, _07399_);
  not (_07404_, _07403_);
  nor (_07405_, _07404_, _07394_);
  nand (_07406_, _07405_, _07387_);
  or (_07407_, _07406_, _07138_);
  or (_07408_, _07168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_07409_, _05826_, _05824_);
  nor (_07410_, _07409_, _05827_);
  nor (_07411_, _07410_, _05657_);
  not (_07412_, _07411_);
  or (_07413_, _05469_, _06603_);
  and (_07414_, _06600_, ABINPUT000000[2]);
  and (_07415_, _06606_, ABINPUT000[2]);
  nor (_07416_, _07415_, _07414_);
  and (_07417_, _07416_, _07413_);
  and (_07418_, _05535_, _05367_);
  and (_07419_, _05537_, _05355_);
  nor (_07420_, _07419_, _07418_);
  and (_07421_, _07420_, _07417_);
  and (_07422_, _07421_, _06177_);
  and (_07423_, _06592_, _05537_);
  nor (_07424_, _07423_, _06593_);
  nor (_07425_, _07424_, _06591_);
  and (_07426_, _06167_, _05590_);
  or (_07427_, _07426_, _05848_);
  and (_07428_, _07427_, _05855_);
  nor (_07429_, _07427_, _05855_);
  or (_07430_, _07429_, _07428_);
  and (_07431_, _07430_, _05844_);
  nor (_07432_, _07431_, _07425_);
  and (_07433_, _07432_, _07422_);
  and (_07434_, _07433_, _07412_);
  nand (_07435_, _07434_, _07168_);
  and (_07436_, _07435_, _07408_);
  or (_07437_, _07436_, _06619_);
  and (_07438_, _07437_, _05141_);
  and (_05717_, _07438_, _07407_);
  or (_07439_, _06905_, _06901_);
  nor (_07440_, _06906_, _05845_);
  nand (_07441_, _07440_, _07439_);
  nor (_07442_, _05930_, _06958_);
  and (_07444_, _07442_, _05944_);
  nor (_07445_, _07444_, _05584_);
  and (_07447_, _07444_, _05584_);
  nor (_07448_, _07447_, _07445_);
  and (_07450_, _07448_, _05481_);
  nor (_07451_, _05893_, _05346_);
  nor (_07452_, _05581_, _06598_);
  and (_07453_, _06600_, ABINPUT000000[9]);
  or (_07455_, _07453_, _07452_);
  nor (_07456_, _07455_, _07451_);
  and (_07458_, _05509_, _05535_);
  and (_07459_, _06606_, ABINPUT000[9]);
  nor (_07461_, _07459_, _07458_);
  and (_07462_, _07461_, _07456_);
  not (_07463_, _07462_);
  nor (_07464_, _07463_, _07450_);
  nand (_07466_, _07464_, _07441_);
  or (_07467_, _07466_, _07138_);
  or (_07468_, _07168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_07469_, _05883_, _05535_);
  and (_07471_, _05936_, _05896_);
  nor (_07472_, _07471_, _07469_);
  and (_07473_, _05535_, _05355_);
  not (_07474_, _07473_);
  and (_07476_, _06606_, ABINPUT000[1]);
  and (_07478_, _05381_, _05892_);
  and (_07479_, _06600_, ABINPUT000000[1]);
  or (_07480_, _07479_, _07478_);
  nor (_07481_, _07480_, _07476_);
  and (_07482_, _07481_, _07474_);
  and (_07483_, _07482_, _07472_);
  and (_07484_, _07483_, _05588_);
  nor (_07485_, _05825_, _05381_);
  nor (_07486_, _07485_, _05855_);
  not (_07487_, _07486_);
  nor (_07488_, _05844_, _05656_);
  nor (_07489_, _07488_, _07487_);
  or (_07490_, _05446_, _06603_);
  and (_07491_, _07490_, _05600_);
  and (_07492_, _07491_, _05594_);
  not (_07494_, _07492_);
  nor (_07495_, _07494_, _07489_);
  and (_07496_, _07495_, _07484_);
  nand (_07497_, _07496_, _07168_);
  and (_07498_, _07497_, _07468_);
  or (_07499_, _07498_, _06619_);
  and (_07500_, _07499_, _05141_);
  and (_05720_, _07500_, _07467_);
  and (_05726_, _06363_, _05141_);
  and (_05729_, _06337_, _05141_);
  and (_05732_, _06389_, _05141_);
  nor (_05735_, _06415_, rst);
  and (_05738_, _06447_, _05141_);
  and (_05741_, _06497_, _05141_);
  and (_05744_, _06524_, _05141_);
  nor (_07501_, _06271_, _05731_);
  nor (_07502_, _06308_, _06487_);
  nor (_07503_, _06314_, _06484_);
  nor (_07504_, _07503_, _07502_);
  and (_07505_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_07506_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_07507_, _07506_, _07505_);
  nor (_07508_, _06304_, _06482_);
  nor (_07509_, _06320_, _06489_);
  nor (_07510_, _07509_, _07508_);
  and (_07511_, _07510_, _07507_);
  and (_07512_, _07511_, _07504_);
  nor (_07513_, _07512_, _07135_);
  nor (_07514_, _07513_, _07501_);
  nor (_05756_, _07514_, rst);
  nor (_07515_, _06271_, _05408_);
  not (_07516_, _06271_);
  and (_07517_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_07518_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor (_07519_, _06320_, _06343_);
  nor (_07520_, _07519_, _07518_);
  nor (_07521_, _06308_, _06347_);
  and (_07522_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_07523_, _07522_, _07521_);
  not (_07524_, _06304_);
  and (_07525_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_07526_, _06314_, _06351_);
  nor (_07527_, _07526_, _07525_);
  and (_07528_, _07527_, _07523_);
  and (_07529_, _07528_, _07520_);
  nor (_07530_, _07529_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07531_, _07530_, _07517_);
  nor (_07532_, _07531_, _07516_);
  nor (_07533_, _07532_, _07515_);
  nor (_05760_, _07533_, rst);
  nor (_07534_, _06271_, _05449_);
  and (_07535_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07536_, _06308_, _06379_);
  nor (_07537_, _06320_, _06374_);
  nor (_07538_, _07537_, _07536_);
  and (_07539_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor (_07540_, _06314_, _06376_);
  nor (_07541_, _07540_, _07539_);
  and (_07542_, _07541_, _07538_);
  and (_07543_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_07544_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_07545_, _07544_, _07543_);
  and (_07546_, _07545_, _07542_);
  nor (_07547_, _07546_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07548_, _07547_, _07535_);
  nor (_07549_, _07548_, _07516_);
  nor (_07550_, _07549_, _07534_);
  nor (_05764_, _07550_, rst);
  and (_07551_, _07516_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_07552_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_07554_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_07555_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_07556_, _07555_, _07554_);
  and (_07557_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor (_07559_, _06314_, _06403_);
  nor (_07560_, _07559_, _07557_);
  nor (_07561_, _06320_, _06395_);
  nor (_07563_, _06308_, _06399_);
  nor (_07564_, _07563_, _07561_);
  and (_07566_, _07564_, _07560_);
  and (_07567_, _07566_, _07556_);
  nor (_07568_, _07567_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07570_, _07568_, _07552_);
  nor (_07571_, _07570_, _07516_);
  nor (_07572_, _07571_, _07551_);
  nor (_05767_, _07572_, rst);
  nor (_07574_, _06271_, _05307_);
  and (_07576_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_07577_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor (_07579_, _06320_, _06429_);
  nor (_07580_, _07579_, _07577_);
  not (_07581_, _06308_);
  and (_07582_, _07581_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_07583_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_07584_, _07583_, _07582_);
  and (_07585_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_07586_, _06314_, _06427_);
  nor (_07587_, _07586_, _07585_);
  and (_07588_, _07587_, _07584_);
  and (_07589_, _07588_, _07580_);
  nor (_07590_, _07589_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07591_, _07590_, _07576_);
  nor (_07592_, _07591_, _07516_);
  nor (_07593_, _07592_, _07574_);
  nor (_05770_, _07593_, rst);
  nand (_07594_, _07200_, _06624_);
  or (_07595_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_07596_, _07595_, _05141_);
  and (_05780_, _07596_, _07594_);
  or (_07597_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand (_07598_, _07434_, _06624_);
  and (_07599_, _07598_, _05141_);
  and (_05783_, _07599_, _07597_);
  or (_07600_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_07601_, _07496_, _06624_);
  and (_07602_, _07601_, _05141_);
  and (_05790_, _07602_, _07600_);
  nand (_07603_, _07259_, _06624_);
  or (_07604_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_07605_, _07604_, _05141_);
  and (_05793_, _07605_, _07603_);
  and (_07606_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_07607_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_07608_, pc_log_change, _07607_);
  or (_07609_, _07608_, _07606_);
  and (_05932_, _07609_, _05141_);
  nor (_07610_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  not (_07611_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_07612_, _07611_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor (_07613_, _07612_, _07610_);
  not (_07614_, \oc8051_symbolic_cxrom1.regvalid [13]);
  not (_07615_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_07617_, _06307_, _06302_);
  nor (_07618_, _07617_, _07516_);
  nor (_07619_, _07618_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_07620_, _07619_, _07615_);
  nor (_07621_, _07620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_07622_, _07620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_07623_, _07622_, _07621_);
  nor (_07624_, _07623_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_07625_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _07611_);
  nor (_07626_, _07625_, _07624_);
  and (_07627_, _07626_, _07614_);
  nor (_07628_, _07626_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_07629_, _07628_, _07627_);
  not (_07630_, _07629_);
  nor (_07631_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_07632_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _07611_);
  nor (_07633_, _07632_, _07631_);
  not (_07634_, _07633_);
  and (_07635_, _07619_, _07615_);
  nor (_07636_, _07635_, _07620_);
  nor (_07637_, _07636_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_07638_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _07611_);
  nor (_07639_, _07638_, _07637_);
  and (_07640_, _07639_, _07634_);
  nand (_07641_, _07640_, _07630_);
  and (_07642_, _07641_, _07613_);
  nor (_07643_, _07639_, _07634_);
  not (_07644_, _07643_);
  not (_07645_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_07646_, _07626_, _07645_);
  and (_07647_, _07626_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_07648_, _07647_, _07646_);
  nor (_07649_, _07648_, _07644_);
  and (_07650_, _07639_, _07633_);
  not (_07651_, _07650_);
  not (_07652_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_07653_, _07626_, _07652_);
  and (_07654_, _07626_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_07656_, _07654_, _07653_);
  nor (_07657_, _07656_, _07651_);
  nor (_07659_, _07657_, _07649_);
  not (_07661_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_07662_, _07626_, _07661_);
  nor (_07663_, _07626_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_07665_, _07663_);
  nor (_07666_, _07639_, _07633_);
  nand (_07668_, _07666_, _07665_);
  or (_07669_, _07668_, _07662_);
  and (_07671_, _07669_, _07659_);
  and (_07673_, _07671_, _07642_);
  and (_07674_, _07626_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_07675_, _07674_, _07643_);
  not (_07676_, _07626_);
  and (_07678_, _07643_, _07676_);
  and (_07679_, _07678_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_07681_, _07679_, _07613_);
  or (_07683_, _07681_, _07675_);
  not (_07684_, _07666_);
  and (_07685_, _07626_, \oc8051_symbolic_cxrom1.regvalid [8]);
  not (_07686_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_07688_, _07626_, _07686_);
  nor (_07689_, _07688_, _07685_);
  nor (_07690_, _07689_, _07684_);
  not (_07691_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_07692_, _07626_, _07691_);
  nor (_07693_, _07626_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_07694_, _07693_, _07692_);
  nor (_07695_, _07694_, _07651_);
  not (_07696_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_07697_, _07626_, _07696_);
  nor (_07698_, _07626_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_07699_, _07698_, _07697_);
  not (_07700_, _07699_);
  and (_07701_, _07700_, _07640_);
  or (_07702_, _07701_, _07695_);
  or (_07703_, _07702_, _07690_);
  nor (_07704_, _07703_, _07683_);
  nor (_07705_, _07704_, _07673_);
  not (_07706_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_07707_, _07613_, _07706_);
  or (_07708_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_07709_, _07708_, _07707_);
  and (_07710_, _07709_, _07650_);
  not (_07711_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_07712_, _07613_, _07711_);
  or (_07713_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_07714_, _07713_, _07712_);
  and (_07715_, _07714_, _07643_);
  or (_07716_, _07715_, _07710_);
  not (_07717_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_07718_, _07613_, _07717_);
  or (_07719_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_07720_, _07719_, _07718_);
  and (_07721_, _07720_, _07640_);
  not (_07722_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_07723_, _07613_, _07722_);
  or (_07724_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_07725_, _07724_, _07723_);
  and (_07726_, _07725_, _07666_);
  or (_07727_, _07726_, _07721_);
  or (_07728_, _07727_, _07716_);
  and (_07729_, _07728_, _07626_);
  not (_07730_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_07731_, _07613_, _07730_);
  or (_07732_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_07733_, _07732_, _07731_);
  and (_07734_, _07733_, _07643_);
  not (_07735_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_07736_, _07613_, _07735_);
  or (_07737_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_07738_, _07737_, _07736_);
  and (_07739_, _07738_, _07650_);
  or (_07740_, _07739_, _07734_);
  not (_07741_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_07742_, _07613_, _07741_);
  or (_07743_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_07744_, _07743_, _07742_);
  and (_07745_, _07744_, _07640_);
  not (_07746_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_07747_, _07613_, _07746_);
  or (_07748_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_07750_, _07748_, _07747_);
  and (_07751_, _07750_, _07666_);
  or (_07752_, _07751_, _07745_);
  or (_07753_, _07752_, _07740_);
  and (_07754_, _07753_, _07676_);
  or (_07756_, _07754_, _07729_);
  and (_07757_, _07756_, _07705_);
  not (_07758_, _07705_);
  and (_07759_, _07758_, word_in[7]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _07759_, _07757_);
  nor (_07761_, _07633_, _07613_);
  not (_07763_, _07761_);
  and (_07765_, _07633_, _07613_);
  and (_07766_, _07765_, _07639_);
  nor (_07768_, _07765_, _07639_);
  nor (_07769_, _07768_, _07766_);
  not (_07771_, _07769_);
  nor (_07772_, _07771_, _07629_);
  not (_07773_, _07766_);
  and (_07774_, _07773_, _07626_);
  not (_07776_, _07639_);
  nor (_07777_, _07776_, _07626_);
  and (_07779_, _07777_, _07765_);
  nor (_07780_, _07779_, _07774_);
  and (_07781_, _07780_, _07771_);
  and (_07782_, _07781_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_07783_, _07780_, _07769_);
  and (_07784_, _07783_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_07785_, _07784_, _07782_);
  nor (_07786_, _07785_, _07772_);
  nor (_07787_, _07786_, _07763_);
  and (_07788_, _07634_, _07613_);
  not (_07789_, _07788_);
  nor (_07790_, _07771_, _07694_);
  and (_07791_, _07781_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_07792_, _07783_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_07793_, _07792_, _07791_);
  nor (_07794_, _07793_, _07790_);
  nor (_07795_, _07794_, _07789_);
  nor (_07796_, _07795_, _07787_);
  not (_07797_, _07613_);
  and (_07798_, _07633_, _07797_);
  not (_07799_, _07798_);
  nor (_07800_, _07771_, _07656_);
  and (_07801_, _07781_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_07802_, _07783_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_07803_, _07802_, _07801_);
  nor (_07804_, _07803_, _07800_);
  nor (_07805_, _07804_, _07799_);
  not (_07806_, _07765_);
  and (_07807_, _07769_, _07676_);
  and (_07808_, _07807_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_07809_, _07783_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_07810_, _07781_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_07811_, _07769_, _07626_);
  and (_07812_, _07811_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_07813_, _07812_, _07810_);
  or (_07814_, _07813_, _07809_);
  nor (_07815_, _07814_, _07808_);
  nor (_07817_, _07815_, _07806_);
  nor (_07818_, _07817_, _07805_);
  and (_07819_, _07818_, _07796_);
  or (_07820_, _07761_, _07765_);
  not (_07821_, _07820_);
  not (_07822_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_07823_, _07613_, _07822_);
  or (_07824_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_07825_, _07824_, _07823_);
  and (_07826_, _07825_, _07821_);
  not (_07827_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_07828_, _07613_, _07827_);
  or (_07829_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_07830_, _07829_, _07828_);
  and (_07831_, _07830_, _07820_);
  or (_07832_, _07831_, _07826_);
  and (_07833_, _07832_, _07783_);
  not (_07834_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_07835_, _07613_, _07834_);
  or (_07836_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_07837_, _07836_, _07835_);
  and (_07838_, _07837_, _07821_);
  not (_07839_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_07840_, _07613_, _07839_);
  or (_07841_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_07842_, _07841_, _07840_);
  and (_07843_, _07842_, _07820_);
  or (_07844_, _07843_, _07838_);
  and (_07845_, _07844_, _07781_);
  not (_07846_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_07847_, _07613_, _07846_);
  or (_07848_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_07849_, _07848_, _07847_);
  and (_07850_, _07849_, _07821_);
  not (_07851_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_07852_, _07613_, _07851_);
  or (_07853_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_07854_, _07853_, _07852_);
  and (_07855_, _07854_, _07820_);
  or (_07856_, _07855_, _07850_);
  and (_07857_, _07856_, _07807_);
  not (_07858_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_07859_, _07613_, _07858_);
  or (_07860_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_07861_, _07860_, _07859_);
  and (_07862_, _07861_, _07821_);
  not (_07864_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_07865_, _07613_, _07864_);
  or (_07867_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_07868_, _07867_, _07865_);
  and (_07870_, _07868_, _07820_);
  or (_07871_, _07870_, _07862_);
  and (_07872_, _07871_, _07811_);
  or (_07874_, _07872_, _07857_);
  or (_07875_, _07874_, _07845_);
  nor (_07877_, _07875_, _07833_);
  nor (_07878_, _07877_, _07819_);
  and (_07880_, _07819_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _07880_, _07878_);
  nor (_07882_, _07666_, _07650_);
  not (_07883_, _07882_);
  nor (_07884_, _07883_, _07629_);
  nor (_07886_, _07650_, _07626_);
  and (_07887_, _07650_, _07626_);
  nor (_07888_, _07887_, _07886_);
  and (_07889_, _07888_, _07883_);
  and (_07890_, _07889_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_07891_, _07888_, _07882_);
  and (_07892_, _07891_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_07893_, _07892_, _07890_);
  nor (_07894_, _07893_, _07884_);
  nor (_07895_, _07894_, _07806_);
  and (_07896_, _07891_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_07897_, _07896_);
  nor (_07898_, _07883_, _07656_);
  and (_07899_, _07889_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_07900_, _07899_, _07898_);
  and (_07901_, _07900_, _07897_);
  nor (_07902_, _07901_, _07789_);
  nor (_07903_, _07902_, _07895_);
  nor (_07904_, _07883_, _07694_);
  and (_07905_, _07889_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_07906_, _07891_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_07907_, _07906_, _07905_);
  nor (_07908_, _07907_, _07904_);
  nor (_07909_, _07908_, _07763_);
  nor (_07910_, _07883_, _07699_);
  and (_07911_, _07889_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_07912_, _07891_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_07913_, _07912_, _07911_);
  nor (_07914_, _07913_, _07910_);
  nor (_07915_, _07914_, _07799_);
  nor (_07916_, _07915_, _07909_);
  and (_07917_, _07916_, _07903_);
  and (_07918_, _07917_, word_in[23]);
  and (_07919_, _07744_, _07643_);
  and (_07920_, _07733_, _07666_);
  or (_07921_, _07920_, _07919_);
  and (_07922_, _07738_, _07640_);
  and (_07923_, _07750_, _07650_);
  or (_07924_, _07923_, _07922_);
  or (_07925_, _07924_, _07921_);
  or (_07926_, _07925_, _07888_);
  not (_07927_, _07888_);
  and (_07928_, _07720_, _07643_);
  and (_07929_, _07714_, _07666_);
  or (_07930_, _07929_, _07928_);
  and (_07931_, _07709_, _07640_);
  and (_07932_, _07725_, _07650_);
  or (_07933_, _07932_, _07931_);
  or (_07934_, _07933_, _07930_);
  or (_07935_, _07934_, _07927_);
  nand (_07936_, _07935_, _07926_);
  nor (_07937_, _07936_, _07917_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _07937_, _07918_);
  nor (_07938_, _07763_, _07639_);
  not (_07939_, _07938_);
  nand (_07940_, _07763_, _07639_);
  and (_07941_, _07940_, _07939_);
  not (_07942_, _07941_);
  nor (_07943_, _07699_, _07942_);
  nor (_07944_, _07940_, _07626_);
  and (_07945_, _07940_, _07626_);
  nor (_07946_, _07945_, _07944_);
  and (_07947_, _07946_, _07942_);
  and (_07948_, _07947_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_07949_, _07946_, _07941_);
  and (_07950_, _07949_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_07951_, _07950_, _07948_);
  nor (_07952_, _07951_, _07943_);
  nor (_07954_, _07952_, _07789_);
  and (_07955_, _07938_, _07646_);
  nor (_07956_, _07942_, _07656_);
  and (_07958_, _07949_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_07959_, _07958_, _07956_);
  and (_07960_, _07959_, _07761_);
  nor (_07962_, _07960_, _07955_);
  not (_07963_, _07962_);
  nor (_07964_, _07963_, _07954_);
  nor (_07966_, _07694_, _07942_);
  and (_07967_, _07949_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_07968_, _07947_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_07970_, _07968_, _07967_);
  nor (_07972_, _07970_, _07966_);
  nor (_07973_, _07972_, _07806_);
  nor (_07975_, _07942_, _07629_);
  and (_07977_, _07949_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_07978_, _07947_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_07979_, _07978_, _07977_);
  nor (_07980_, _07979_, _07975_);
  nor (_07982_, _07980_, _07799_);
  nor (_07983_, _07982_, _07973_);
  and (_07984_, _07983_, _07964_);
  and (_07985_, _07842_, _07821_);
  and (_07986_, _07837_, _07820_);
  or (_07987_, _07986_, _07985_);
  and (_07988_, _07987_, _07947_);
  and (_07989_, _07830_, _07821_);
  and (_07990_, _07825_, _07820_);
  or (_07991_, _07990_, _07989_);
  and (_07992_, _07991_, _07949_);
  and (_07993_, _07941_, _07676_);
  and (_07994_, _07854_, _07821_);
  and (_07995_, _07849_, _07820_);
  or (_07996_, _07995_, _07994_);
  and (_07997_, _07996_, _07993_);
  and (_07998_, _07868_, _07821_);
  and (_07999_, _07861_, _07820_);
  or (_08000_, _07999_, _07998_);
  and (_08001_, _07945_, _07939_);
  and (_08002_, _08001_, _08000_);
  or (_08003_, _08002_, _07997_);
  or (_08004_, _08003_, _07992_);
  nor (_08005_, _08004_, _07988_);
  nor (_08006_, _08005_, _07984_);
  and (_08007_, _07984_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08007_, _08006_);
  and (_08008_, _07639_, _07626_);
  or (_08009_, _08008_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_06029_, _08009_, _05141_);
  and (_08010_, _07984_, _05141_);
  and (_08011_, _08010_, word_in[31]);
  and (_08012_, _08008_, _07761_);
  and (_08013_, _08010_, _08012_);
  and (_08014_, _08013_, _08011_);
  not (_08015_, _08013_);
  and (_08016_, _07917_, _05141_);
  and (_08017_, _08016_, _07882_);
  and (_08018_, _08017_, _07888_);
  and (_08019_, _08018_, _07788_);
  not (_08020_, _08019_);
  and (_08021_, _07819_, _05141_);
  and (_08022_, _08021_, _07798_);
  and (_08023_, _08022_, _07811_);
  and (_08024_, _07673_, _05141_);
  and (_08025_, _08024_, _07633_);
  nor (_08026_, _07705_, rst);
  and (_08027_, _08026_, _08008_);
  and (_08028_, _08027_, _08025_);
  and (_08029_, _08026_, word_in[7]);
  and (_08030_, _08029_, _08028_);
  nor (_08031_, _08028_, _07706_);
  nor (_08032_, _08031_, _08030_);
  nor (_08033_, _08032_, _08023_);
  and (_08034_, _08023_, word_in[15]);
  or (_08035_, _08034_, _08033_);
  and (_08036_, _08035_, _08020_);
  and (_08037_, _08016_, word_in[23]);
  and (_08038_, _08037_, _08019_);
  or (_08039_, _08038_, _08036_);
  and (_08040_, _08039_, _08015_);
  or (_06058_, _08040_, _08014_);
  or (_08041_, _07947_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_06079_, _08041_, _05141_);
  and (_08043_, _07798_, _07947_);
  and (_08044_, _07766_, _07626_);
  and (_08046_, _07666_, _07676_);
  or (_08047_, _08046_, _08044_);
  or (_08049_, _08047_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08050_, _08049_, _08043_);
  and (_06108_, _08050_, _05141_);
  and (_08052_, _07993_, _07798_);
  or (_08054_, _08052_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08055_, _08054_, _08047_);
  and (_06149_, _08055_, _05141_);
  or (_08057_, _07639_, _07626_);
  nand (_08059_, _08057_, _07645_);
  and (_06196_, _08059_, _05141_);
  or (_08061_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand (_08062_, _07619_, _06347_);
  and (_08063_, _08062_, _05141_);
  and (_06232_, _08063_, _08061_);
  and (_08064_, _07993_, _07765_);
  and (_08065_, _07777_, _07761_);
  or (_08066_, _08065_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_08067_, _08066_, _08057_);
  nor (_08068_, _08067_, _08064_);
  nor (_08069_, _08068_, _07781_);
  and (_08070_, _07821_, _07993_);
  and (_08071_, _07938_, _07676_);
  or (_08072_, _08071_, _08044_);
  and (_08073_, _08072_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_08074_, _08073_, _08070_);
  or (_08075_, _08074_, _08069_);
  and (_06252_, _08075_, _05141_);
  not (_08076_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_08077_, _05622_, _08076_);
  not (_08078_, _05622_);
  nor (_08079_, _06062_, _08078_);
  or (_08080_, _08079_, _08077_);
  and (_06258_, _08080_, _05141_);
  not (_08081_, _08057_);
  nor (_08082_, _08081_, _08044_);
  not (_08083_, _07886_);
  or (_08084_, _08065_, _08064_);
  or (_08085_, _08084_, _08083_);
  and (_08086_, _08085_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08087_, _07788_, _07777_);
  and (_08088_, _08046_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08089_, _08052_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08090_, _08089_, _08088_);
  or (_08091_, _08090_, _08087_);
  or (_08092_, _08091_, _08086_);
  or (_08093_, _07774_, _07944_);
  and (_08094_, _08093_, _08092_);
  and (_08095_, _07993_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08096_, _08095_, _08065_);
  or (_08097_, _08096_, _08094_);
  and (_08098_, _08097_, _08082_);
  and (_08099_, _08092_, _08044_);
  and (_08100_, _08071_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08101_, _07788_, _07993_);
  and (_08102_, _08101_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08103_, _08102_, _08052_);
  or (_08104_, _08103_, _08100_);
  or (_08105_, _08104_, _08064_);
  or (_08106_, _08105_, _08099_);
  or (_08107_, _08106_, _08098_);
  and (_06294_, _08107_, _05141_);
  nand (_08108_, _07639_, _07613_);
  nand (_08109_, _07886_, _08108_);
  and (_08110_, _07798_, _07777_);
  or (_08111_, _08110_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08112_, _08111_, _08109_);
  and (_08113_, _08112_, _08083_);
  and (_08114_, _08084_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08115_, _08114_, _08087_);
  or (_08116_, _08115_, _08113_);
  and (_08117_, _08116_, _08093_);
  and (_08118_, _08111_, _08044_);
  and (_08119_, _08052_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08121_, _08046_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08122_, _08121_, _08064_);
  or (_08124_, _08122_, _08119_);
  or (_08125_, _08124_, _08065_);
  or (_08126_, _08125_, _08118_);
  or (_08127_, _08126_, _08117_);
  and (_06359_, _08127_, _05141_);
  and (_08128_, _05622_, _05522_);
  not (_08129_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_08130_, _05622_, _08129_);
  or (_08131_, _08130_, _08128_);
  and (_06405_, _08131_, _05141_);
  not (_08132_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_08133_, _05622_, _08132_);
  nor (_08134_, _08078_, _05560_);
  or (_08135_, _08134_, _08133_);
  and (_06424_, _08135_, _05141_);
  and (_08136_, _07821_, _07777_);
  and (_08137_, _07941_, _07653_);
  and (_08138_, _07938_, _07653_);
  or (_08139_, _08138_, _08065_);
  or (_08140_, _08139_, _08137_);
  or (_08142_, _07766_, _07626_);
  and (_08143_, _07653_, _07776_);
  or (_08144_, _08110_, _07626_);
  and (_08145_, _08144_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_08146_, _07633_, _07652_);
  and (_08147_, _08146_, _07777_);
  or (_08148_, _08147_, _07779_);
  or (_08149_, _08148_, _08145_);
  or (_08150_, _08149_, _08143_);
  and (_08151_, _08150_, _08142_);
  or (_08152_, _08151_, _08140_);
  or (_08153_, _08152_, _08136_);
  and (_06435_, _08153_, _05141_);
  and (_08154_, _06179_, _05622_);
  not (_08155_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_08156_, _05622_, _08155_);
  or (_08157_, _08156_, _08154_);
  and (_06443_, _08157_, _05141_);
  not (_08158_, _06836_);
  nor (_08159_, _06207_, _05708_);
  or (_08160_, _08159_, _06208_);
  or (_08161_, _06838_, _06836_);
  nor (_08162_, _08161_, _06841_);
  and (_08163_, _08162_, _06881_);
  nand (_08164_, _08163_, _08160_);
  and (_08165_, _06884_, _06669_);
  and (_08166_, _05256_, _05172_);
  and (_08167_, _08166_, _06879_);
  and (_08168_, _08167_, _05241_);
  and (_08169_, _08168_, _05647_);
  not (_08170_, _08169_);
  and (_08171_, _08170_, _08162_);
  and (_08172_, _08171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_08173_, _08172_, _08165_);
  nand (_08174_, _08173_, _08164_);
  nand (_08175_, _08174_, _08158_);
  nand (_08176_, _07288_, _06836_);
  nand (_08177_, _08176_, _08175_);
  and (_06503_, _08177_, _05141_);
  and (_08178_, _05922_, _05288_);
  nor (_08179_, _05288_, _05441_);
  or (_08180_, _08179_, _08178_);
  nand (_08181_, _08180_, _08163_);
  and (_08182_, _08171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_08183_, _07434_, _06842_);
  nor (_08184_, _08183_, _08182_);
  and (_08185_, _08184_, _08158_);
  nand (_08186_, _08185_, _08181_);
  or (_08187_, _07406_, _08158_);
  and (_08188_, _08187_, _08186_);
  and (_06507_, _08188_, _05141_);
  and (_08189_, _07938_, _07626_);
  or (_08190_, _08189_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08191_, _08190_, _07626_);
  not (_08192_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_08193_, _08057_, _08192_);
  and (_08194_, _08065_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_08195_, _08087_, _07779_);
  or (_08196_, _08195_, _08194_);
  or (_08197_, _08196_, _08193_);
  or (_08198_, _08197_, _08191_);
  or (_08199_, _08198_, _08110_);
  and (_06513_, _08199_, _05141_);
  and (_08200_, _07886_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08201_, _07939_, _07626_);
  and (_08202_, _08201_, _07773_);
  and (_08203_, _08001_, _07788_);
  nor (_08204_, _07886_, _07661_);
  or (_08205_, _08204_, _08203_);
  and (_08206_, _08205_, _08202_);
  and (_08207_, _07650_, _07676_);
  and (_08208_, _08207_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_08209_, _08208_, _08189_);
  or (_08211_, _08209_, _08206_);
  and (_08212_, _08211_, _07774_);
  and (_08213_, _08205_, _08044_);
  or (_08214_, _08213_, _08207_);
  or (_08215_, _08214_, _08212_);
  or (_08216_, _08215_, _08200_);
  and (_06609_, _08216_, _05141_);
  and (_08217_, _07798_, _07945_);
  not (_08218_, _07768_);
  and (_08220_, _08218_, _07674_);
  or (_08221_, _08220_, _08217_);
  and (_08222_, _08046_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08223_, _07882_, _07676_);
  and (_08225_, _08223_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08226_, _08110_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08227_, _08226_, _07779_);
  or (_08228_, _08227_, _08225_);
  or (_08230_, _08228_, _08222_);
  or (_08231_, _08230_, _08203_);
  or (_08232_, _08231_, _08189_);
  or (_08233_, _08232_, _08221_);
  and (_06704_, _08233_, _05141_);
  and (_08235_, _06004_, _05622_);
  not (_08237_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_08238_, _05622_, _08237_);
  or (_08239_, _08238_, _08235_);
  and (_06712_, _08239_, _05141_);
  and (_08241_, _05648_, _05281_);
  and (_08242_, _06736_, _05288_);
  and (_08243_, _08242_, _08241_);
  and (_08245_, _06691_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_08246_, _08245_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or (_08247_, _08246_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_08248_, _08246_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_08249_, _08248_, rst);
  nand (_08250_, _08249_, _08247_);
  nor (_06717_, _08250_, _08243_);
  and (_08251_, _06281_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_08252_, _06275_, _05561_);
  or (_08253_, _08252_, _08251_);
  and (_06783_, _08253_, _05141_);
  and (_08254_, _07945_, _07765_);
  and (_08255_, _08008_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08256_, _08255_, _08254_);
  not (_08257_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08258_, _07626_, _08257_);
  or (_08259_, _08189_, _08217_);
  or (_08260_, _08259_, _08258_);
  or (_08261_, _08260_, _08203_);
  or (_08262_, _08261_, _08256_);
  and (_06794_, _08262_, _05141_);
  and (_08263_, _08248_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_08264_, _08263_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_08265_, _08263_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_08266_, _08265_, _08264_);
  nand (_08267_, _08266_, _05141_);
  nor (_06817_, _08267_, _08243_);
  and (_08268_, _08008_, _07763_);
  and (_08269_, _08268_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08270_, _07678_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_08271_, _08189_, _08046_);
  or (_08272_, _08271_, _07777_);
  and (_08273_, _08272_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_08274_, _08273_, _08001_);
  or (_08275_, _08274_, _08270_);
  or (_08276_, _08275_, _08269_);
  and (_06887_, _08276_, _05141_);
  or (_08277_, _08248_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_08278_, _08263_, rst);
  nand (_08279_, _08278_, _08277_);
  nor (_06903_, _08279_, _08243_);
  and (_08280_, _06012_, _06202_);
  and (_08281_, _05922_, _06032_);
  or (_08282_, _05650_, _06007_);
  not (_08283_, _08282_);
  and (_08284_, _08283_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_08285_, _08284_, _08281_);
  and (_08286_, _08285_, _08280_);
  nand (_08287_, _08280_, _05186_);
  and (_08288_, _08287_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_08289_, _08241_, _05926_);
  or (_08290_, _08289_, _08288_);
  or (_08291_, _08290_, _08286_);
  nand (_08292_, _08289_, _06062_);
  and (_08293_, _08292_, _05141_);
  and (_06957_, _08293_, _08291_);
  not (_08294_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_08295_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_08296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _08295_);
  nand (_08297_, _08296_, _08294_);
  or (_08298_, _08296_, rxd_i);
  and (_08299_, _08298_, _08297_);
  nor (_08300_, _06683_, _06690_);
  and (_08301_, _08300_, _06686_);
  and (_08302_, _08301_, _08299_);
  nor (_08303_, _08301_, _08294_);
  or (_08304_, _08303_, rst);
  or (_06960_, _08304_, _08302_);
  and (_08305_, _06621_, _06008_);
  not (_08306_, _08305_);
  or (_08307_, _08306_, _06004_);
  or (_08308_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_08309_, _08308_, _05141_);
  and (_06962_, _08309_, _08307_);
  nand (_08311_, _08305_, _05604_);
  or (_08313_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_08315_, _08313_, _05141_);
  and (_06966_, _08315_, _08311_);
  nor (_08316_, _07634_, _07626_);
  or (_08318_, _08316_, _07887_);
  and (_08319_, _08318_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_08320_, _07643_, _07626_);
  or (_08322_, _08012_, _08320_);
  nor (_08323_, _08008_, _07614_);
  or (_08324_, _08323_, _08268_);
  and (_08326_, _08324_, _07634_);
  or (_08327_, _08326_, _08322_);
  or (_08328_, _08327_, _08319_);
  and (_06971_, _08328_, _05141_);
  not (_08330_, _06821_);
  and (_08332_, _06765_, _06536_);
  and (_08333_, _06574_, _06449_);
  and (_08334_, _08333_, _06536_);
  or (_08336_, _08334_, _06784_);
  nor (_08337_, _08336_, _08332_);
  or (_08338_, _08337_, _08330_);
  nor (_08339_, _06538_, _06474_);
  and (_08340_, _08339_, _06550_);
  and (_08341_, _08340_, _07088_);
  not (_08342_, _08341_);
  and (_08343_, _08342_, _06796_);
  nand (_08344_, _08343_, _08338_);
  and (_06984_, _08344_, _05141_);
  not (_08345_, _06738_);
  nor (_08346_, _08345_, _06244_);
  and (_08347_, _06736_, _06032_);
  and (_08348_, _08347_, _06734_);
  and (_08349_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_08350_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_08351_, _08350_, _08349_);
  nor (_08352_, _08351_, _06738_);
  or (_08353_, _08352_, _08348_);
  or (_08354_, _08353_, _08346_);
  not (_08355_, _08348_);
  or (_08356_, _08355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_08357_, _08356_, _05141_);
  and (_06991_, _08357_, _08354_);
  and (_08358_, _08280_, _06207_);
  nand (_08359_, _08358_, _05963_);
  not (_08360_, _08289_);
  or (_08361_, _08358_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_08362_, _08361_, _08360_);
  and (_08363_, _08362_, _08359_);
  nor (_08364_, _08360_, _06244_);
  or (_08365_, _08364_, _08363_);
  and (_07024_, _08365_, _05141_);
  not (_08366_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand (_08367_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _08366_);
  or (_08368_, _08367_, _06683_);
  nor (_08369_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_08370_, _08369_, _08368_);
  or (_08371_, _08370_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_08372_, _08371_, _08280_);
  and (_08373_, _05922_, _05210_);
  not (_08374_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_08375_, _05210_, _08374_);
  nand (_08376_, _08375_, _08280_);
  or (_08377_, _08376_, _08373_);
  and (_08378_, _08377_, _08372_);
  or (_08379_, _08378_, _08289_);
  nand (_08380_, _08289_, _05604_);
  and (_08381_, _08380_, _05141_);
  and (_07027_, _08381_, _08379_);
  and (_08382_, _08243_, _06683_);
  and (_08383_, _08382_, _05561_);
  and (_08384_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_08385_, _08384_, _06683_);
  nor (_08386_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_08387_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_08388_, _08387_, _08386_);
  and (_08389_, _08388_, _08246_);
  nor (_08390_, _08389_, _08385_);
  not (_08391_, _08390_);
  and (_08392_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_08393_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_08394_, _08393_, _08392_);
  nor (_08395_, _08394_, _08243_);
  and (_08396_, _08243_, _06691_);
  and (_08397_, _08396_, _06179_);
  or (_08398_, _08397_, _08395_);
  or (_08399_, _08398_, _08383_);
  and (_07038_, _08399_, _05141_);
  and (_08401_, _07319_, _06836_);
  and (_08402_, _06881_, _06032_);
  nand (_08404_, _08402_, _05963_);
  not (_08405_, _08162_);
  nor (_08406_, _08402_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_08408_, _08406_, _08405_);
  and (_08409_, _08408_, _08404_);
  nor (_08411_, _07350_, _06842_);
  or (_08412_, _08411_, _08409_);
  and (_08414_, _08412_, _08158_);
  or (_08415_, _08414_, _08401_);
  and (_07061_, _08415_, _05141_);
  nor (_08417_, _06738_, _06730_);
  or (_08418_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  not (_08420_, _08417_);
  or (_08422_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_08423_, _08422_, _08418_);
  and (_08424_, _08423_, _08355_);
  nor (_08425_, _08355_, _06062_);
  or (_08426_, _08425_, _08424_);
  and (_07075_, _08426_, _05141_);
  or (_08427_, _07811_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_07082_, _08427_, _05141_);
  nand (_08428_, _06743_, _06244_);
  or (_08429_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_08430_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_08431_, _08430_, _08429_);
  or (_08432_, _08431_, _06743_);
  and (_08433_, _08432_, _05141_);
  and (_07095_, _08433_, _08428_);
  and (_08434_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not (_08435_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_08436_, \oc8051_top_1.oc8051_sfr1.pres_ow , _08435_);
  nor (_08437_, _08436_, _08434_);
  not (_08438_, _08437_);
  and (_08439_, _08438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_08440_, _08439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  not (_08441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor (_08442_, _06727_, _08441_);
  and (_08443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_08444_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_08445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_08446_, _08445_, _08444_);
  and (_08447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_08448_, _08447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_08449_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_08450_, _08449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_08451_, _08450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_08452_, _08451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_08453_, _08452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_08454_, _08453_, _08446_);
  and (_08455_, _08454_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_08456_, _08455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_08457_, _08456_, _08443_);
  nand (_08458_, _08457_, _08442_);
  nand (_08459_, _08458_, _08440_);
  not (_08460_, _06726_);
  not (_08461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_08462_, _06725_, _08461_);
  nor (_08463_, _08462_, _08460_);
  not (_08464_, _08463_);
  or (_08465_, _08439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_08466_, _08465_, _08464_);
  and (_08467_, _08466_, _08459_);
  and (_08468_, _08463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_08469_, _05209_, _06007_);
  and (_08470_, _06736_, _08469_);
  and (_08471_, _08470_, _06734_);
  or (_08472_, _08471_, _08468_);
  or (_08474_, _08472_, _08467_);
  nand (_08475_, _08471_, _05604_);
  and (_08476_, _05964_, _05925_);
  and (_08478_, _08476_, _06734_);
  not (_08479_, _08478_);
  and (_08480_, _08479_, _08475_);
  and (_08481_, _08480_, _08474_);
  and (_08482_, _08478_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_08483_, _08482_, _08481_);
  and (_07098_, _08483_, _05141_);
  not (_08484_, _05277_);
  nor (_08485_, _06062_, _08484_);
  not (_08487_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_08488_, _05277_, _08487_);
  or (_08489_, _08488_, _05572_);
  or (_08491_, _08489_, _08485_);
  or (_08492_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_08494_, _08492_, _05141_);
  and (_07122_, _08494_, _08491_);
  nand (_08496_, _07466_, _06836_);
  nor (_08497_, _05210_, _05420_);
  or (_08499_, _08497_, _08373_);
  nand (_08500_, _08499_, _08163_);
  nor (_08501_, _06881_, _05420_);
  nor (_08503_, _08501_, _06884_);
  and (_08504_, _08503_, _08500_);
  nor (_08505_, _07496_, _06836_);
  nor (_08507_, _08505_, _08162_);
  or (_08508_, _08507_, _08504_);
  nand (_08509_, _08508_, _08496_);
  and (_07160_, _08509_, _05141_);
  and (_08511_, _08396_, _06703_);
  and (_08512_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_08513_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_08514_, _08513_, _08512_);
  nor (_08515_, _08514_, _08243_);
  and (_08516_, _08382_, _06179_);
  or (_08518_, _08516_, _08515_);
  or (_08519_, _08518_, _08511_);
  and (_07165_, _08519_, _05141_);
  and (_08520_, _05299_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_08521_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_08522_, _08521_, _05303_);
  and (_08523_, _06179_, _05523_);
  or (_08524_, _08523_, _08522_);
  or (_08525_, _08524_, _08520_);
  and (_07247_, _08525_, _05141_);
  and (_08526_, _08016_, _08043_);
  not (_08527_, _08526_);
  and (_08528_, _08021_, _08044_);
  not (_08529_, _08528_);
  and (_08530_, _08026_, _07633_);
  nor (_08531_, _08530_, _08024_);
  and (_08532_, _08026_, _08081_);
  and (_08533_, _08532_, _08531_);
  and (_08534_, _08533_, word_in[0]);
  not (_08535_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_08536_, _08533_, _08535_);
  or (_08537_, _08536_, _08534_);
  and (_08538_, _08537_, _08529_);
  and (_08539_, _08528_, word_in[8]);
  or (_08540_, _08539_, _08538_);
  and (_08541_, _08540_, _08527_);
  and (_08542_, _07788_, _08008_);
  and (_08543_, _08010_, _08542_);
  and (_08544_, _08016_, word_in[16]);
  and (_08545_, _08544_, _08043_);
  or (_08546_, _08545_, _08543_);
  or (_08547_, _08546_, _08541_);
  not (_08548_, _08543_);
  or (_08549_, _08548_, word_in[24]);
  and (_07443_, _08549_, _08547_);
  or (_08550_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not (_08551_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_08552_, pc_log_change, _08551_);
  and (_08553_, _08552_, _05141_);
  and (_07446_, _08553_, _08550_);
  not (_08554_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_08555_, _08533_, _08554_);
  and (_08556_, _08026_, word_in[1]);
  and (_08557_, _08556_, _08533_);
  or (_08558_, _08557_, _08555_);
  or (_08559_, _08558_, _08528_);
  or (_08560_, _08529_, word_in[9]);
  and (_08561_, _08560_, _08559_);
  or (_08562_, _08561_, _08526_);
  nor (_08563_, _08527_, word_in[17]);
  nor (_08564_, _08563_, _08543_);
  and (_08565_, _08564_, _08562_);
  and (_08566_, _08010_, word_in[25]);
  and (_08567_, _08566_, _08543_);
  or (_07449_, _08567_, _08565_);
  and (_08568_, _08010_, word_in[26]);
  and (_08569_, _08568_, _08543_);
  not (_08570_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_08571_, _08533_, _08570_);
  and (_08572_, _08026_, word_in[2]);
  and (_08573_, _08572_, _08533_);
  or (_08574_, _08573_, _08571_);
  or (_08575_, _08574_, _08528_);
  or (_08576_, _08529_, word_in[10]);
  and (_08577_, _08576_, _08575_);
  or (_08578_, _08577_, _08526_);
  nor (_08579_, _08527_, word_in[18]);
  nor (_08580_, _08579_, _08543_);
  and (_08581_, _08580_, _08578_);
  or (_07454_, _08581_, _08569_);
  nor (_07457_, _05625_, rst);
  and (_08582_, _08010_, word_in[27]);
  and (_08583_, _08582_, _08543_);
  not (_08584_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_08585_, _08533_, _08584_);
  and (_08586_, _08026_, word_in[3]);
  and (_08587_, _08586_, _08533_);
  or (_08588_, _08587_, _08585_);
  and (_08589_, _08588_, _08529_);
  and (_08590_, _08528_, word_in[11]);
  or (_08591_, _08590_, _08589_);
  or (_08592_, _08591_, _08526_);
  nor (_08593_, _08527_, word_in[19]);
  nor (_08594_, _08593_, _08543_);
  and (_08595_, _08594_, _08592_);
  or (_07460_, _08595_, _08583_);
  not (_08596_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_08597_, _08533_, _08596_);
  and (_08598_, _08026_, word_in[4]);
  and (_08599_, _08598_, _08533_);
  or (_08600_, _08599_, _08597_);
  or (_08601_, _08600_, _08528_);
  or (_08602_, _08529_, word_in[12]);
  and (_08603_, _08602_, _08601_);
  or (_08604_, _08603_, _08526_);
  nor (_08605_, _08527_, word_in[20]);
  nor (_08606_, _08605_, _08543_);
  and (_08607_, _08606_, _08604_);
  and (_08608_, _08010_, word_in[28]);
  and (_08609_, _08608_, _08543_);
  or (_07465_, _08609_, _08607_);
  not (_08610_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_08611_, _08533_, _08610_);
  and (_08612_, _08026_, word_in[5]);
  and (_08613_, _08612_, _08533_);
  or (_08614_, _08613_, _08611_);
  or (_08615_, _08614_, _08528_);
  or (_08616_, _08529_, word_in[13]);
  and (_08617_, _08616_, _08615_);
  or (_08618_, _08617_, _08526_);
  nor (_08619_, _08527_, word_in[21]);
  nor (_08620_, _08619_, _08543_);
  and (_08621_, _08620_, _08618_);
  and (_08622_, _08010_, word_in[29]);
  and (_08623_, _08622_, _08543_);
  or (_07470_, _08623_, _08621_);
  and (_08624_, _08010_, word_in[30]);
  and (_08625_, _08624_, _08543_);
  not (_08626_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_08627_, _08533_, _08626_);
  and (_08628_, _08026_, word_in[6]);
  and (_08629_, _08628_, _08533_);
  or (_08630_, _08629_, _08627_);
  or (_08631_, _08630_, _08528_);
  or (_08632_, _08529_, word_in[14]);
  and (_08633_, _08632_, _08631_);
  or (_08634_, _08633_, _08526_);
  nor (_08635_, _08527_, word_in[22]);
  nor (_08636_, _08635_, _08543_);
  and (_08637_, _08636_, _08634_);
  or (_07475_, _08637_, _08625_);
  nor (_08638_, _08533_, _07839_);
  and (_08639_, _08533_, _08029_);
  or (_08640_, _08639_, _08638_);
  or (_08641_, _08640_, _08528_);
  not (_08642_, word_in[15]);
  nand (_08643_, _08528_, _08642_);
  and (_08644_, _08643_, _08641_);
  or (_08645_, _08644_, _08526_);
  or (_08646_, _08527_, word_in[23]);
  and (_08647_, _08646_, _08548_);
  and (_08648_, _08647_, _08645_);
  and (_08649_, _08543_, word_in[31]);
  or (_07477_, _08649_, _08648_);
  and (_08650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_08651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_08652_, _05626_, _08651_);
  not (_08653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_08654_, _08653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_08655_, _08654_, _08652_);
  nor (_08656_, _08655_, _08650_);
  or (_08657_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_08658_, _08657_, _05141_);
  nor (_07493_, _08658_, _08656_);
  and (_08659_, _08010_, _08043_);
  not (_08660_, _08659_);
  and (_08661_, _08016_, _07765_);
  and (_08662_, _08661_, _07891_);
  not (_08663_, _08662_);
  and (_08664_, _08021_, _07761_);
  and (_08665_, _08664_, _07781_);
  and (_08666_, _08026_, word_in[0]);
  and (_08667_, _08026_, _08057_);
  and (_08668_, _08024_, _07634_);
  not (_08669_, _08668_);
  nor (_08670_, _08669_, _08667_);
  and (_08671_, _08670_, _08666_);
  not (_08672_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_08673_, _08670_, _08672_);
  nor (_08674_, _08673_, _08671_);
  nor (_08675_, _08674_, _08665_);
  and (_08676_, _08665_, word_in[8]);
  or (_08677_, _08676_, _08675_);
  and (_08678_, _08677_, _08663_);
  and (_08680_, _08662_, _08544_);
  or (_08681_, _08680_, _08678_);
  and (_08683_, _08681_, _08660_);
  and (_08684_, _08659_, word_in[24]);
  or (_07553_, _08684_, _08683_);
  not (_08685_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_08686_, _08670_, _08685_);
  and (_08687_, _08670_, _08556_);
  nor (_08688_, _08687_, _08686_);
  nor (_08689_, _08688_, _08665_);
  and (_08690_, _08665_, word_in[9]);
  or (_08692_, _08690_, _08689_);
  and (_08693_, _08692_, _08663_);
  and (_08694_, _08016_, word_in[17]);
  and (_08695_, _08662_, _08694_);
  or (_08696_, _08695_, _08693_);
  and (_08697_, _08696_, _08660_);
  and (_08698_, _08659_, word_in[25]);
  or (_07558_, _08698_, _08697_);
  and (_08699_, _08670_, _08572_);
  not (_08700_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_08701_, _08670_, _08700_);
  nor (_08702_, _08701_, _08699_);
  nor (_08703_, _08702_, _08665_);
  and (_08704_, _08665_, word_in[10]);
  or (_08705_, _08704_, _08703_);
  and (_08706_, _08705_, _08663_);
  and (_08707_, _08016_, word_in[18]);
  and (_08708_, _08662_, _08707_);
  or (_08709_, _08708_, _08706_);
  and (_08710_, _08709_, _08660_);
  and (_08711_, _08659_, word_in[26]);
  or (_07562_, _08711_, _08710_);
  and (_08712_, _08016_, word_in[19]);
  and (_08713_, _08662_, _08712_);
  not (_08714_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_08715_, _08670_, _08714_);
  and (_08716_, _08670_, _08586_);
  nor (_08717_, _08716_, _08715_);
  nor (_08718_, _08717_, _08665_);
  and (_08719_, _08665_, word_in[11]);
  or (_08720_, _08719_, _08718_);
  and (_08721_, _08720_, _08663_);
  or (_08722_, _08721_, _08713_);
  and (_08723_, _08722_, _08660_);
  and (_08724_, _08659_, word_in[27]);
  or (_07565_, _08724_, _08723_);
  and (_08725_, _08670_, _08598_);
  not (_08726_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_08727_, _08670_, _08726_);
  nor (_08728_, _08727_, _08725_);
  nor (_08729_, _08728_, _08665_);
  and (_08730_, _08665_, word_in[12]);
  or (_08731_, _08730_, _08729_);
  and (_08732_, _08731_, _08663_);
  and (_08733_, _08016_, word_in[20]);
  and (_08734_, _08662_, _08733_);
  or (_08735_, _08734_, _08732_);
  and (_08736_, _08735_, _08660_);
  and (_08737_, _08659_, word_in[28]);
  or (_07569_, _08737_, _08736_);
  and (_08738_, _08670_, _08612_);
  not (_08739_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_08740_, _08670_, _08739_);
  nor (_08741_, _08740_, _08738_);
  nor (_08742_, _08741_, _08665_);
  and (_08743_, _08665_, word_in[13]);
  or (_08744_, _08743_, _08742_);
  and (_08745_, _08744_, _08663_);
  and (_08746_, _08016_, word_in[21]);
  and (_08747_, _08662_, _08746_);
  or (_08748_, _08747_, _08745_);
  and (_08749_, _08748_, _08660_);
  and (_08750_, _08659_, word_in[29]);
  or (_07573_, _08750_, _08749_);
  and (_08751_, _08670_, _08628_);
  not (_08752_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_08753_, _08670_, _08752_);
  nor (_08754_, _08753_, _08751_);
  nor (_08755_, _08754_, _08665_);
  and (_08756_, _08665_, word_in[14]);
  or (_08757_, _08756_, _08755_);
  and (_08758_, _08757_, _08663_);
  and (_08759_, _08016_, word_in[22]);
  and (_08760_, _08662_, _08759_);
  or (_08761_, _08760_, _08758_);
  and (_08762_, _08761_, _08660_);
  and (_08763_, _08659_, word_in[30]);
  or (_07575_, _08763_, _08762_);
  nor (_08764_, _08670_, _07746_);
  and (_08765_, _08670_, _08029_);
  or (_08766_, _08765_, _08764_);
  or (_08767_, _08766_, _08665_);
  nand (_08768_, _08665_, _08642_);
  and (_08769_, _08768_, _08767_);
  or (_08771_, _08769_, _08662_);
  or (_08772_, _08663_, _08037_);
  and (_08773_, _08772_, _08660_);
  and (_08774_, _08773_, _08771_);
  and (_08776_, _08659_, word_in[31]);
  or (_07578_, _08776_, _08774_);
  and (_08778_, _08016_, _07761_);
  and (_08779_, _08778_, _07891_);
  not (_08780_, _08779_);
  and (_08782_, _08021_, _07788_);
  and (_08783_, _08782_, _07781_);
  not (_08784_, _08024_);
  and (_08786_, _08530_, _08784_);
  and (_08787_, _08786_, _08081_);
  and (_08789_, _08787_, _08666_);
  not (_08790_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor (_08791_, _08787_, _08790_);
  nor (_08793_, _08791_, _08789_);
  nor (_08794_, _08793_, _08783_);
  and (_08795_, _08783_, word_in[8]);
  or (_08797_, _08795_, _08794_);
  and (_08798_, _08797_, _08780_);
  and (_08799_, _08010_, _07765_);
  and (_08800_, _08799_, _07947_);
  and (_08801_, _08779_, _08544_);
  or (_08802_, _08801_, _08800_);
  or (_08803_, _08802_, _08798_);
  not (_08804_, _08800_);
  or (_08805_, _08804_, word_in[24]);
  and (_07655_, _08805_, _08803_);
  and (_08806_, _05563_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_08807_, _06004_, _05523_);
  or (_08808_, _08807_, _08806_);
  and (_07658_, _08808_, _05141_);
  and (_08809_, _08787_, _08556_);
  not (_08810_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_08811_, _08787_, _08810_);
  nor (_08812_, _08811_, _08809_);
  nor (_08813_, _08812_, _08783_);
  and (_08814_, _08783_, word_in[9]);
  or (_08815_, _08814_, _08813_);
  and (_08816_, _08815_, _08780_);
  and (_08817_, _08779_, _08694_);
  or (_08818_, _08817_, _08800_);
  or (_08819_, _08818_, _08816_);
  or (_08820_, _08804_, word_in[25]);
  and (_07660_, _08820_, _08819_);
  and (_08822_, _08787_, _08572_);
  not (_08823_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_08824_, _08787_, _08823_);
  nor (_08825_, _08824_, _08822_);
  nor (_08826_, _08825_, _08783_);
  and (_08827_, _08783_, word_in[10]);
  or (_08828_, _08827_, _08826_);
  and (_08829_, _08828_, _08780_);
  and (_08830_, _08779_, word_in[18]);
  or (_08831_, _08830_, _08800_);
  or (_08832_, _08831_, _08829_);
  or (_08833_, _08804_, word_in[26]);
  and (_07664_, _08833_, _08832_);
  and (_08834_, _08779_, word_in[19]);
  and (_08835_, _08787_, _08586_);
  not (_08836_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_08837_, _08787_, _08836_);
  nor (_08838_, _08837_, _08835_);
  nor (_08839_, _08838_, _08783_);
  and (_08840_, _08783_, word_in[11]);
  or (_08841_, _08840_, _08839_);
  and (_08842_, _08841_, _08780_);
  or (_08843_, _08842_, _08834_);
  and (_08844_, _08843_, _08804_);
  and (_08845_, _08800_, word_in[27]);
  or (_07667_, _08845_, _08844_);
  and (_08846_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_08847_, _06004_, _05617_);
  or (_08848_, _08847_, _08846_);
  and (_07670_, _08848_, _05141_);
  and (_08849_, _08787_, _08598_);
  not (_08850_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_08851_, _08787_, _08850_);
  nor (_08852_, _08851_, _08849_);
  nor (_08853_, _08852_, _08783_);
  and (_08854_, _08783_, word_in[12]);
  or (_08855_, _08854_, _08853_);
  and (_08856_, _08855_, _08780_);
  and (_08857_, _08779_, word_in[20]);
  or (_08858_, _08857_, _08800_);
  or (_08860_, _08858_, _08856_);
  or (_08861_, _08804_, word_in[28]);
  and (_07672_, _08861_, _08860_);
  not (_08862_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_08863_, _08787_, _08862_);
  and (_08864_, _08787_, _08612_);
  or (_08865_, _08864_, _08863_);
  or (_08866_, _08865_, _08783_);
  not (_08868_, _08783_);
  or (_08869_, _08868_, word_in[13]);
  and (_08871_, _08869_, _08866_);
  or (_08872_, _08871_, _08779_);
  or (_08874_, _08780_, word_in[21]);
  and (_08875_, _08874_, _08804_);
  and (_08876_, _08875_, _08872_);
  and (_08878_, _08800_, word_in[29]);
  or (_07677_, _08878_, _08876_);
  and (_08880_, _05614_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nand (_08881_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_08883_, _08881_, _05609_);
  and (_08884_, _05605_, _05283_);
  or (_08885_, _08884_, _08883_);
  or (_08886_, _08885_, _08880_);
  and (_07680_, _08886_, _05141_);
  and (_08888_, _08787_, _08628_);
  not (_08890_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_08891_, _08787_, _08890_);
  nor (_08892_, _08891_, _08888_);
  nor (_08893_, _08892_, _08783_);
  and (_08894_, _08783_, word_in[14]);
  or (_08895_, _08894_, _08893_);
  and (_08896_, _08895_, _08780_);
  and (_08897_, _08779_, _08759_);
  or (_08898_, _08897_, _08800_);
  or (_08899_, _08898_, _08896_);
  or (_08900_, _08804_, word_in[30]);
  and (_07682_, _08900_, _08899_);
  and (_08901_, _08787_, _08029_);
  nor (_08902_, _08787_, _07834_);
  or (_08903_, _08902_, _08901_);
  or (_08904_, _08903_, _08783_);
  nand (_08905_, _08783_, _08642_);
  and (_08906_, _08905_, _08780_);
  and (_08907_, _08906_, _08904_);
  and (_08908_, _08779_, _08037_);
  or (_08909_, _08908_, _08800_);
  or (_08910_, _08909_, _08907_);
  or (_08911_, _08804_, word_in[31]);
  and (_07687_, _08911_, _08910_);
  or (_08912_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand (_08913_, _07619_, _06399_);
  and (_08914_, _08913_, _05141_);
  and (_07749_, _08914_, _08912_);
  and (_08915_, _08010_, _08071_);
  not (_08916_, _08915_);
  and (_08917_, _08016_, _07788_);
  and (_08918_, _08917_, _07891_);
  not (_08919_, _08918_);
  and (_08920_, _08022_, _07781_);
  not (_08921_, _08025_);
  nor (_08922_, _08667_, _08921_);
  and (_08923_, _08922_, _08666_);
  not (_08924_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor (_08925_, _08922_, _08924_);
  nor (_08926_, _08925_, _08923_);
  nor (_08927_, _08926_, _08920_);
  and (_08928_, _08920_, word_in[8]);
  or (_08929_, _08928_, _08927_);
  and (_08930_, _08929_, _08919_);
  and (_08931_, _08918_, word_in[16]);
  or (_08932_, _08931_, _08930_);
  and (_08933_, _08932_, _08916_);
  and (_08934_, _08915_, word_in[24]);
  or (_07755_, _08934_, _08933_);
  and (_08935_, _08918_, word_in[17]);
  and (_08936_, _08922_, _08556_);
  not (_08937_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_08938_, _08922_, _08937_);
  nor (_08939_, _08938_, _08936_);
  nor (_08940_, _08939_, _08920_);
  and (_08941_, _08920_, word_in[9]);
  or (_08942_, _08941_, _08940_);
  and (_08943_, _08942_, _08919_);
  or (_08944_, _08943_, _08935_);
  and (_08945_, _08944_, _08916_);
  and (_08946_, _08915_, word_in[25]);
  or (_07760_, _08946_, _08945_);
  and (_08947_, _08915_, word_in[26]);
  and (_08948_, _08922_, _08572_);
  not (_08949_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_08950_, _08922_, _08949_);
  nor (_08951_, _08950_, _08948_);
  nor (_08952_, _08951_, _08920_);
  and (_08953_, _08920_, word_in[10]);
  or (_08954_, _08953_, _08952_);
  or (_08955_, _08954_, _08918_);
  or (_08956_, _08919_, _08707_);
  and (_08957_, _08956_, _08916_);
  and (_08958_, _08957_, _08955_);
  or (_07762_, _08958_, _08947_);
  and (_08959_, _08922_, _08586_);
  not (_08960_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_08961_, _08922_, _08960_);
  nor (_08962_, _08961_, _08959_);
  nor (_08963_, _08962_, _08920_);
  and (_08964_, _08920_, word_in[11]);
  or (_08965_, _08964_, _08963_);
  and (_08966_, _08965_, _08919_);
  and (_08967_, _08918_, word_in[19]);
  or (_08968_, _08967_, _08915_);
  or (_08969_, _08968_, _08966_);
  or (_08970_, _08916_, word_in[27]);
  and (_07764_, _08970_, _08969_);
  and (_08971_, _08922_, _08598_);
  not (_08972_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_08973_, _08922_, _08972_);
  nor (_08974_, _08973_, _08971_);
  nor (_08975_, _08974_, _08920_);
  and (_08976_, _08920_, word_in[12]);
  or (_08977_, _08976_, _08975_);
  and (_08978_, _08977_, _08919_);
  and (_08979_, _08918_, word_in[20]);
  or (_08980_, _08979_, _08915_);
  or (_08981_, _08980_, _08978_);
  or (_08982_, _08916_, word_in[28]);
  and (_07767_, _08982_, _08981_);
  and (_08983_, _08922_, _08612_);
  not (_08984_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_08985_, _08922_, _08984_);
  nor (_08986_, _08985_, _08983_);
  nor (_08987_, _08986_, _08920_);
  and (_08988_, _08920_, word_in[13]);
  or (_08989_, _08988_, _08987_);
  and (_08990_, _08989_, _08919_);
  and (_08992_, _08918_, _08746_);
  or (_08993_, _08992_, _08915_);
  or (_08994_, _08993_, _08990_);
  or (_08995_, _08916_, word_in[29]);
  and (_07770_, _08995_, _08994_);
  and (_08996_, _08915_, word_in[30]);
  and (_08997_, _08922_, _08628_);
  not (_08998_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_08999_, _08922_, _08998_);
  nor (_09000_, _08999_, _08997_);
  nor (_09001_, _09000_, _08920_);
  and (_09002_, _08920_, word_in[14]);
  or (_09003_, _09002_, _09001_);
  or (_09004_, _09003_, _08918_);
  or (_09005_, _08919_, _08759_);
  and (_09006_, _09005_, _08916_);
  and (_09007_, _09006_, _09004_);
  or (_07775_, _09007_, _08996_);
  nor (_09008_, _08922_, _07730_);
  and (_09009_, _08922_, _08029_);
  or (_09010_, _09009_, _09008_);
  or (_09011_, _09010_, _08920_);
  nand (_09012_, _08920_, _08642_);
  and (_09013_, _09012_, _09011_);
  or (_09014_, _09013_, _08918_);
  or (_09015_, _08919_, _08037_);
  and (_09016_, _09015_, _08916_);
  and (_09017_, _09016_, _09014_);
  and (_09018_, _08915_, word_in[31]);
  or (_07778_, _09018_, _09017_);
  and (_09019_, _08017_, _07927_);
  and (_09020_, _09019_, _07798_);
  not (_09021_, _09020_);
  and (_09022_, _08021_, _08064_);
  not (_09023_, _09022_);
  or (_09024_, _09023_, word_in[8]);
  not (_09025_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_09026_, _08026_, _07777_);
  and (_09027_, _09026_, _08531_);
  nor (_09028_, _09027_, _09025_);
  and (_09029_, _09027_, word_in[0]);
  or (_09030_, _09029_, _09028_);
  or (_09031_, _09030_, _09022_);
  and (_09032_, _09031_, _09024_);
  and (_09033_, _09032_, _09021_);
  and (_09034_, _08010_, _07941_);
  and (_09035_, _09034_, _07946_);
  and (_09036_, _09035_, _07788_);
  and (_09037_, _09020_, _08544_);
  or (_09038_, _09037_, _09036_);
  or (_09039_, _09038_, _09033_);
  and (_09040_, _08010_, word_in[24]);
  not (_09041_, _09036_);
  or (_09042_, _09041_, _09040_);
  and (_07863_, _09042_, _09039_);
  not (_09043_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_09044_, _09027_, _09043_);
  and (_09045_, _09027_, word_in[1]);
  or (_09046_, _09045_, _09044_);
  and (_09047_, _09046_, _09023_);
  and (_09048_, _09022_, word_in[9]);
  or (_09049_, _09048_, _09047_);
  and (_09050_, _09049_, _09021_);
  and (_09051_, _09020_, _08694_);
  or (_09052_, _09051_, _09036_);
  or (_09053_, _09052_, _09050_);
  or (_09054_, _09041_, _08566_);
  and (_07866_, _09054_, _09053_);
  not (_09055_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_09056_, _09027_, _09055_);
  and (_09057_, _09027_, word_in[2]);
  or (_09058_, _09057_, _09056_);
  or (_09059_, _09058_, _09022_);
  or (_09060_, _09023_, word_in[10]);
  and (_09061_, _09060_, _09059_);
  and (_09062_, _09061_, _09021_);
  and (_09063_, _09020_, _08707_);
  or (_09064_, _09063_, _09036_);
  or (_09065_, _09064_, _09062_);
  or (_09066_, _09041_, _08568_);
  and (_07869_, _09066_, _09065_);
  not (_09067_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_09068_, _09027_, _09067_);
  and (_09069_, _09027_, word_in[3]);
  or (_09070_, _09069_, _09068_);
  and (_09071_, _09070_, _09023_);
  and (_09072_, _09022_, word_in[11]);
  or (_09073_, _09072_, _09071_);
  and (_09074_, _09073_, _09021_);
  and (_09075_, _09020_, _08712_);
  or (_09076_, _09075_, _09036_);
  or (_09077_, _09076_, _09074_);
  or (_09078_, _09041_, _08582_);
  and (_07873_, _09078_, _09077_);
  not (_09079_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_09080_, _09027_, _09079_);
  and (_09081_, _09027_, word_in[4]);
  or (_09082_, _09081_, _09080_);
  or (_09083_, _09082_, _09022_);
  or (_09084_, _09023_, word_in[12]);
  and (_09085_, _09084_, _09083_);
  and (_09086_, _09085_, _09021_);
  and (_09087_, _09020_, _08733_);
  or (_09088_, _09087_, _09036_);
  or (_09089_, _09088_, _09086_);
  or (_09090_, _09041_, _08608_);
  and (_07876_, _09090_, _09089_);
  not (_09091_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_09092_, _09027_, _09091_);
  and (_09093_, _09027_, word_in[5]);
  or (_09094_, _09093_, _09092_);
  and (_09095_, _09094_, _09023_);
  and (_09096_, _09022_, word_in[13]);
  or (_09097_, _09096_, _09095_);
  and (_09098_, _09097_, _09021_);
  and (_09099_, _09020_, _08746_);
  or (_09100_, _09099_, _09036_);
  or (_09101_, _09100_, _09098_);
  or (_09102_, _09041_, _08622_);
  and (_07879_, _09102_, _09101_);
  not (_09103_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_09104_, _09027_, _09103_);
  and (_09105_, _09027_, word_in[6]);
  or (_09106_, _09105_, _09104_);
  and (_09107_, _09106_, _09023_);
  and (_09108_, _09022_, word_in[14]);
  or (_09110_, _09108_, _09107_);
  and (_09111_, _09110_, _09021_);
  and (_09112_, _09020_, _08759_);
  or (_09113_, _09112_, _09036_);
  or (_09114_, _09113_, _09111_);
  or (_09115_, _09041_, _08624_);
  and (_07881_, _09115_, _09114_);
  nor (_09116_, _09027_, _07851_);
  and (_09117_, _09027_, word_in[7]);
  or (_09118_, _09117_, _09116_);
  and (_09120_, _09118_, _09023_);
  and (_09121_, _09022_, word_in[15]);
  or (_09122_, _09121_, _09120_);
  and (_09123_, _09122_, _09021_);
  and (_09124_, _09020_, _08037_);
  or (_09125_, _09124_, _09036_);
  or (_09126_, _09125_, _09123_);
  or (_09127_, _09041_, _08011_);
  and (_07885_, _09127_, _09126_);
  and (_09128_, _08664_, _07807_);
  not (_09129_, _09128_);
  or (_09130_, _09129_, word_in[8]);
  and (_09131_, _09019_, _07765_);
  not (_09132_, _09131_);
  not (_09133_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_09134_, _09026_, _08668_);
  nor (_09135_, _09134_, _09133_);
  and (_09136_, _09134_, word_in[0]);
  or (_09137_, _09136_, _09135_);
  or (_09138_, _09137_, _09128_);
  and (_09139_, _09138_, _09132_);
  and (_09140_, _09139_, _09130_);
  and (_09141_, _09035_, _07798_);
  and (_09142_, _09131_, _08544_);
  or (_09144_, _09142_, _09141_);
  or (_09145_, _09144_, _09140_);
  not (_09146_, _09141_);
  or (_09147_, _09146_, word_in[24]);
  and (_07953_, _09147_, _09145_);
  and (_09148_, _09131_, _08694_);
  and (_09149_, _09134_, word_in[1]);
  not (_09150_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_09151_, _09134_, _09150_);
  nor (_09152_, _09151_, _09149_);
  nor (_09153_, _09152_, _09128_);
  and (_09154_, _09128_, word_in[9]);
  or (_09155_, _09154_, _09153_);
  and (_09156_, _09155_, _09132_);
  or (_09157_, _09156_, _09148_);
  and (_09158_, _09157_, _09146_);
  and (_09159_, _09141_, word_in[25]);
  or (_07957_, _09159_, _09158_);
  or (_09160_, _09132_, _08707_);
  not (_09161_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_09162_, _09134_, _09161_);
  and (_09163_, _09134_, word_in[2]);
  or (_09164_, _09163_, _09162_);
  or (_09165_, _09164_, _09128_);
  or (_09166_, _09129_, word_in[10]);
  and (_09167_, _09166_, _09165_);
  or (_09168_, _09167_, _09131_);
  and (_09169_, _09168_, _09160_);
  and (_09171_, _09169_, _09146_);
  and (_09172_, _09141_, word_in[26]);
  or (_07961_, _09172_, _09171_);
  or (_09174_, _09132_, _08712_);
  not (_09175_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_09176_, _09134_, _09175_);
  and (_09177_, _09134_, word_in[3]);
  or (_09178_, _09177_, _09176_);
  or (_09179_, _09178_, _09128_);
  or (_09180_, _09129_, word_in[11]);
  and (_09181_, _09180_, _09179_);
  or (_09182_, _09181_, _09131_);
  and (_09183_, _09182_, _09174_);
  or (_09184_, _09183_, _09141_);
  or (_09185_, _09146_, word_in[27]);
  and (_07965_, _09185_, _09184_);
  not (_09186_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_09187_, _09134_, _09186_);
  and (_09188_, _09134_, word_in[4]);
  nor (_09189_, _09188_, _09187_);
  nor (_09190_, _09189_, _09128_);
  and (_09191_, _09128_, word_in[12]);
  or (_09192_, _09191_, _09190_);
  and (_09193_, _09192_, _09132_);
  and (_09194_, _09131_, _08733_);
  or (_09195_, _09194_, _09141_);
  or (_09196_, _09195_, _09193_);
  or (_09197_, _09146_, word_in[28]);
  and (_07969_, _09197_, _09196_);
  not (_09198_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_09199_, _09134_, _09198_);
  and (_09200_, _09134_, word_in[5]);
  nor (_09201_, _09200_, _09199_);
  nor (_09202_, _09201_, _09128_);
  and (_09203_, _09128_, word_in[13]);
  or (_09204_, _09203_, _09202_);
  and (_09205_, _09204_, _09132_);
  and (_09206_, _09131_, _08746_);
  or (_09207_, _09206_, _09141_);
  or (_09208_, _09207_, _09205_);
  or (_09209_, _09146_, word_in[29]);
  and (_07971_, _09209_, _09208_);
  or (_09210_, _09132_, _08759_);
  not (_09211_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_09212_, _09134_, _09211_);
  and (_09213_, _09134_, word_in[6]);
  or (_09214_, _09213_, _09212_);
  or (_09215_, _09214_, _09128_);
  or (_09216_, _09129_, word_in[14]);
  and (_09217_, _09216_, _09215_);
  or (_09218_, _09217_, _09131_);
  and (_09219_, _09218_, _09210_);
  and (_09220_, _09219_, _09146_);
  and (_09221_, _09141_, word_in[30]);
  or (_07974_, _09221_, _09220_);
  or (_09222_, _09132_, _08037_);
  nor (_09223_, _09134_, _07741_);
  and (_09224_, _09134_, word_in[7]);
  or (_09225_, _09224_, _09223_);
  or (_09226_, _09225_, _09128_);
  nand (_09227_, _09128_, _08642_);
  and (_09228_, _09227_, _09226_);
  or (_09229_, _09228_, _09131_);
  and (_09230_, _09229_, _09222_);
  and (_09231_, _09230_, _09146_);
  and (_09232_, _09141_, word_in[31]);
  or (_07976_, _09232_, _09231_);
  and (_09233_, _09035_, _07765_);
  and (_09234_, _09019_, _07761_);
  and (_09235_, _08782_, _07807_);
  not (_09236_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_09237_, _08786_, _07777_);
  nor (_09238_, _09237_, _09236_);
  and (_09239_, _09237_, _08666_);
  or (_09240_, _09239_, _09238_);
  or (_09241_, _09240_, _09235_);
  not (_09242_, _09235_);
  or (_09243_, _09242_, word_in[8]);
  and (_09244_, _09243_, _09241_);
  or (_09245_, _09244_, _09234_);
  not (_09246_, _09234_);
  or (_09247_, _09246_, _08544_);
  and (_09248_, _09247_, _09245_);
  or (_09249_, _09248_, _09233_);
  not (_09250_, _09233_);
  or (_09251_, _09250_, word_in[24]);
  and (_08042_, _09251_, _09249_);
  and (_09252_, _09237_, _08556_);
  not (_09253_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_09254_, _09237_, _09253_);
  nor (_09255_, _09254_, _09252_);
  nor (_09256_, _09255_, _09235_);
  and (_09257_, _09235_, word_in[9]);
  or (_09258_, _09257_, _09256_);
  and (_09259_, _09258_, _09246_);
  and (_09260_, _09234_, _08694_);
  or (_09261_, _09260_, _09233_);
  or (_09262_, _09261_, _09259_);
  or (_09263_, _09250_, word_in[25]);
  and (_08045_, _09263_, _09262_);
  not (_09264_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_09265_, _09237_, _09264_);
  and (_09266_, _09237_, _08572_);
  or (_09267_, _09266_, _09265_);
  or (_09268_, _09267_, _09235_);
  or (_09269_, _09242_, word_in[10]);
  and (_09270_, _09269_, _09268_);
  or (_09271_, _09270_, _09234_);
  or (_09272_, _09246_, _08707_);
  and (_09273_, _09272_, _09271_);
  and (_09274_, _09273_, _09250_);
  and (_09275_, _09233_, word_in[26]);
  or (_08048_, _09275_, _09274_);
  not (_09276_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_09277_, _09237_, _09276_);
  and (_09278_, _09237_, _08586_);
  or (_09279_, _09278_, _09277_);
  or (_09280_, _09279_, _09235_);
  or (_09281_, _09242_, word_in[11]);
  and (_09282_, _09281_, _09280_);
  or (_09283_, _09282_, _09234_);
  or (_09284_, _09246_, _08712_);
  and (_09285_, _09284_, _09283_);
  or (_09286_, _09285_, _09233_);
  or (_09287_, _09250_, word_in[27]);
  and (_08051_, _09287_, _09286_);
  or (_09288_, _09246_, _08733_);
  not (_09289_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_09290_, _09237_, _09289_);
  and (_09291_, _09237_, _08598_);
  or (_09292_, _09291_, _09290_);
  or (_09293_, _09292_, _09235_);
  or (_09294_, _09242_, word_in[12]);
  and (_09295_, _09294_, _09293_);
  or (_09296_, _09295_, _09234_);
  and (_09297_, _09296_, _09288_);
  or (_09298_, _09297_, _09233_);
  or (_09299_, _09250_, word_in[28]);
  and (_08053_, _09299_, _09298_);
  and (_09300_, _09237_, _08612_);
  not (_09301_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_09302_, _09237_, _09301_);
  nor (_09303_, _09302_, _09300_);
  nor (_09304_, _09303_, _09235_);
  and (_09305_, _09235_, word_in[13]);
  or (_09306_, _09305_, _09304_);
  and (_09307_, _09306_, _09246_);
  and (_09308_, _09234_, _08746_);
  or (_09309_, _09308_, _09307_);
  and (_09310_, _09309_, _09250_);
  and (_09311_, _09233_, word_in[29]);
  or (_08056_, _09311_, _09310_);
  and (_09312_, _09237_, _08628_);
  not (_09313_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_09314_, _09237_, _09313_);
  nor (_09315_, _09314_, _09312_);
  nor (_09316_, _09315_, _09235_);
  and (_09317_, _09235_, word_in[14]);
  or (_09318_, _09317_, _09316_);
  and (_09319_, _09318_, _09246_);
  and (_09320_, _09234_, _08759_);
  or (_09321_, _09320_, _09233_);
  or (_09322_, _09321_, _09319_);
  or (_09323_, _09250_, word_in[30]);
  and (_08058_, _09323_, _09322_);
  nor (_09324_, _09237_, _07846_);
  and (_09325_, _09237_, _08029_);
  or (_09326_, _09325_, _09324_);
  or (_09327_, _09326_, _09235_);
  nand (_09328_, _09235_, _08642_);
  and (_09329_, _09328_, _09327_);
  or (_09330_, _09329_, _09234_);
  or (_09331_, _09246_, _08037_);
  and (_09332_, _09331_, _09330_);
  or (_09333_, _09332_, _09233_);
  or (_09334_, _09250_, word_in[31]);
  and (_08060_, _09334_, _09333_);
  and (_09335_, _08010_, _08065_);
  and (_09336_, _09335_, _09040_);
  not (_09337_, _09335_);
  and (_09338_, _09019_, _07788_);
  not (_09339_, _09338_);
  and (_09340_, _08022_, _07807_);
  and (_09341_, _09026_, _08025_);
  and (_09342_, _09341_, word_in[0]);
  not (_09343_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor (_09344_, _09341_, _09343_);
  nor (_09345_, _09344_, _09342_);
  nor (_09346_, _09345_, _09340_);
  and (_09347_, _09340_, word_in[8]);
  or (_09348_, _09347_, _09346_);
  and (_09349_, _09348_, _09339_);
  and (_09350_, _09338_, _08544_);
  or (_09351_, _09350_, _09349_);
  and (_09352_, _09351_, _09337_);
  or (_08120_, _09352_, _09336_);
  and (_09353_, _09338_, _08694_);
  not (_09354_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_09355_, _09341_, _09354_);
  and (_09356_, _09341_, word_in[1]);
  nor (_09357_, _09356_, _09355_);
  nor (_09358_, _09357_, _09340_);
  and (_09359_, _09340_, word_in[9]);
  or (_09360_, _09359_, _09358_);
  and (_09361_, _09360_, _09339_);
  or (_09362_, _09361_, _09353_);
  and (_09363_, _09362_, _09337_);
  and (_09364_, _09335_, word_in[25]);
  or (_08123_, _09364_, _09363_);
  and (_09365_, _09338_, _08707_);
  not (_09366_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_09367_, _09341_, _09366_);
  and (_09368_, _09341_, word_in[2]);
  nor (_09369_, _09368_, _09367_);
  nor (_09370_, _09369_, _09340_);
  and (_09371_, _09340_, word_in[10]);
  or (_09372_, _09371_, _09370_);
  and (_09373_, _09372_, _09339_);
  or (_09374_, _09373_, _09365_);
  and (_09375_, _09374_, _09337_);
  and (_09376_, _09335_, word_in[26]);
  or (_13490_, _09376_, _09375_);
  and (_09377_, _09338_, _08712_);
  not (_09378_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_09379_, _09341_, _09378_);
  and (_09380_, _09341_, word_in[3]);
  nor (_09381_, _09380_, _09379_);
  nor (_09382_, _09381_, _09340_);
  and (_09383_, _09340_, word_in[11]);
  or (_09384_, _09383_, _09382_);
  and (_09385_, _09384_, _09339_);
  or (_09386_, _09385_, _09377_);
  and (_09387_, _09386_, _09337_);
  and (_09388_, _09335_, word_in[27]);
  or (_13491_, _09388_, _09387_);
  and (_09389_, _09338_, _08733_);
  not (_09390_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_09391_, _09341_, _09390_);
  and (_09392_, _09341_, word_in[4]);
  nor (_09393_, _09392_, _09391_);
  nor (_09394_, _09393_, _09340_);
  and (_09395_, _09340_, word_in[12]);
  or (_09396_, _09395_, _09394_);
  and (_09397_, _09396_, _09339_);
  or (_09398_, _09397_, _09389_);
  and (_09399_, _09398_, _09337_);
  and (_09400_, _09335_, word_in[28]);
  or (_13492_, _09400_, _09399_);
  and (_09401_, _09338_, _08746_);
  not (_09402_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_09403_, _09341_, _09402_);
  and (_09404_, _09341_, word_in[5]);
  nor (_09405_, _09404_, _09403_);
  nor (_09406_, _09405_, _09340_);
  and (_09407_, _09340_, word_in[13]);
  or (_09408_, _09407_, _09406_);
  and (_09409_, _09408_, _09339_);
  or (_09410_, _09409_, _09401_);
  and (_09411_, _09410_, _09337_);
  and (_09412_, _09335_, word_in[29]);
  or (_13493_, _09412_, _09411_);
  not (_09413_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_09414_, _09341_, _09413_);
  and (_09415_, _09341_, word_in[6]);
  or (_09416_, _09415_, _09414_);
  or (_09417_, _09416_, _09340_);
  not (_09418_, word_in[14]);
  nand (_09419_, _09340_, _09418_);
  and (_09420_, _09419_, _09417_);
  or (_09421_, _09420_, _09338_);
  or (_09422_, _09339_, _08759_);
  and (_09423_, _09422_, _09337_);
  and (_09424_, _09423_, _09421_);
  and (_09425_, _09335_, word_in[30]);
  or (_13494_, _09425_, _09424_);
  nor (_09426_, _09341_, _07735_);
  and (_09427_, _09341_, word_in[7]);
  or (_09428_, _09427_, _09426_);
  or (_09429_, _09428_, _09340_);
  nand (_09430_, _09340_, _08642_);
  and (_09431_, _09430_, _09429_);
  or (_09432_, _09431_, _09338_);
  or (_09433_, _09339_, _08037_);
  and (_09434_, _09433_, _09432_);
  or (_09435_, _09434_, _09335_);
  or (_09436_, _09337_, word_in[31]);
  and (_08141_, _09436_, _09435_);
  not (_09437_, _08385_);
  not (_09438_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_09439_, _08389_, _09438_);
  and (_09440_, _08389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_09441_, _09440_, _09439_);
  and (_09442_, _09441_, _09437_);
  nor (_09443_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_09444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_09445_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_09446_, _09445_, _09444_);
  nor (_09447_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_09448_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_09449_, _09448_, _09447_);
  and (_09450_, _09449_, _09446_);
  and (_09451_, _09450_, _09443_);
  and (_09452_, _09451_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_09453_, _09452_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_09454_, _09453_, _08385_);
  nor (_09455_, _09454_, _09442_);
  nor (_09456_, _09455_, _08243_);
  nor (_09457_, _06691_, _05604_);
  and (_09458_, _09457_, _08243_);
  or (_09459_, _09458_, _09456_);
  and (_08210_, _09459_, _05141_);
  and (_09460_, _08010_, _07949_);
  and (_09461_, _09460_, _07788_);
  not (_09462_, _09461_);
  and (_09463_, _08016_, _08110_);
  and (_09464_, _09463_, word_in[16]);
  not (_09465_, _09463_);
  and (_09466_, _08021_, _07779_);
  not (_09467_, _09466_);
  not (_09468_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_09469_, _07776_, _07626_);
  and (_09470_, _08026_, _09469_);
  and (_09471_, _09470_, _08531_);
  nor (_09472_, _09471_, _09468_);
  and (_09473_, _09471_, word_in[0]);
  or (_09474_, _09473_, _09472_);
  and (_09475_, _09474_, _09467_);
  and (_09476_, _09466_, word_in[8]);
  or (_09477_, _09476_, _09475_);
  and (_09478_, _09477_, _09465_);
  or (_09479_, _09478_, _09464_);
  and (_09480_, _09479_, _09462_);
  and (_09481_, _09461_, word_in[24]);
  or (_13495_, _09481_, _09480_);
  and (_09482_, _09463_, word_in[17]);
  not (_09483_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_09484_, _09471_, _09483_);
  and (_09485_, _09471_, word_in[1]);
  or (_09486_, _09485_, _09484_);
  and (_09487_, _09486_, _09467_);
  and (_09488_, _09466_, word_in[9]);
  or (_09489_, _09488_, _09487_);
  and (_09490_, _09489_, _09465_);
  or (_09491_, _09490_, _09482_);
  and (_09492_, _09491_, _09462_);
  and (_09493_, _09461_, word_in[25]);
  or (_08219_, _09493_, _09492_);
  and (_09494_, _09463_, word_in[18]);
  not (_09495_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_09496_, _09471_, _09495_);
  and (_09497_, _09471_, word_in[2]);
  or (_09498_, _09497_, _09496_);
  and (_09499_, _09498_, _09467_);
  and (_09500_, _09466_, word_in[10]);
  or (_09501_, _09500_, _09499_);
  and (_09502_, _09501_, _09465_);
  or (_09503_, _09502_, _09494_);
  and (_09504_, _09503_, _09462_);
  and (_09505_, _09461_, word_in[26]);
  or (_08224_, _09505_, _09504_);
  and (_09506_, _09463_, word_in[19]);
  not (_09507_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_09508_, _09471_, _09507_);
  and (_09509_, _09471_, word_in[3]);
  or (_09510_, _09509_, _09508_);
  and (_09511_, _09510_, _09467_);
  and (_09512_, _09466_, word_in[11]);
  or (_09513_, _09512_, _09511_);
  and (_09514_, _09513_, _09465_);
  or (_09515_, _09514_, _09506_);
  and (_09516_, _09515_, _09462_);
  and (_09517_, _09461_, word_in[27]);
  or (_08229_, _09517_, _09516_);
  and (_09518_, _09463_, word_in[20]);
  not (_09519_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_09520_, _09471_, _09519_);
  and (_09521_, _09471_, word_in[4]);
  or (_09522_, _09521_, _09520_);
  and (_09523_, _09522_, _09467_);
  and (_09524_, _09466_, word_in[12]);
  or (_09525_, _09524_, _09523_);
  and (_09526_, _09525_, _09465_);
  or (_09527_, _09526_, _09518_);
  and (_09528_, _09527_, _09462_);
  and (_09529_, _09461_, word_in[28]);
  or (_08234_, _09529_, _09528_);
  and (_09530_, _09463_, word_in[21]);
  not (_09531_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_09532_, _09471_, _09531_);
  and (_09533_, _09471_, word_in[5]);
  or (_09534_, _09533_, _09532_);
  and (_09535_, _09534_, _09467_);
  and (_09536_, _09466_, word_in[13]);
  or (_09537_, _09536_, _09535_);
  and (_09538_, _09537_, _09465_);
  or (_09539_, _09538_, _09530_);
  and (_09540_, _09539_, _09462_);
  and (_09541_, _09461_, word_in[29]);
  or (_08236_, _09541_, _09540_);
  and (_09542_, _09463_, word_in[22]);
  not (_09543_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_09544_, _09471_, _09543_);
  and (_09545_, _09471_, word_in[6]);
  or (_09546_, _09545_, _09544_);
  and (_09547_, _09546_, _09467_);
  and (_09548_, _09466_, word_in[14]);
  or (_09549_, _09548_, _09547_);
  and (_09550_, _09549_, _09465_);
  or (_09551_, _09550_, _09542_);
  and (_09552_, _09551_, _09462_);
  and (_09553_, _09461_, word_in[30]);
  or (_08240_, _09553_, _09552_);
  and (_09554_, _09463_, word_in[23]);
  nor (_09555_, _09471_, _07827_);
  and (_09556_, _09471_, word_in[7]);
  or (_09557_, _09556_, _09555_);
  and (_09558_, _09557_, _09467_);
  and (_09559_, _09466_, word_in[15]);
  or (_09560_, _09559_, _09558_);
  and (_09561_, _09560_, _09465_);
  or (_09562_, _09561_, _09554_);
  and (_09563_, _09562_, _09462_);
  and (_09565_, _09461_, word_in[31]);
  or (_08244_, _09565_, _09563_);
  and (_09566_, _08010_, _08110_);
  not (_09567_, _09566_);
  and (_09568_, _08661_, _07889_);
  and (_09570_, _09568_, _08544_);
  not (_09571_, _09568_);
  and (_09573_, _08664_, _07783_);
  and (_09574_, _09470_, _08668_);
  and (_09575_, _09574_, _08666_);
  not (_09576_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_09577_, _09574_, _09576_);
  nor (_09578_, _09577_, _09575_);
  nor (_09579_, _09578_, _09573_);
  and (_09580_, _09573_, word_in[8]);
  or (_09581_, _09580_, _09579_);
  and (_09582_, _09581_, _09571_);
  or (_09583_, _09582_, _09570_);
  and (_09584_, _09583_, _09567_);
  and (_09585_, _09566_, word_in[24]);
  or (_08310_, _09585_, _09584_);
  and (_09586_, _06695_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_09587_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_09588_, _09587_, _06687_);
  and (_09589_, _09588_, _06697_);
  or (_09590_, _09589_, _09586_);
  and (_08312_, _09590_, _05141_);
  and (_09591_, _09574_, _08556_);
  not (_09592_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_09593_, _09574_, _09592_);
  nor (_09594_, _09593_, _09591_);
  nor (_09595_, _09594_, _09573_);
  and (_09596_, _09573_, word_in[9]);
  or (_09597_, _09596_, _09595_);
  or (_09598_, _09597_, _09568_);
  or (_09599_, _09571_, _08694_);
  and (_09600_, _09599_, _09567_);
  and (_09601_, _09600_, _09598_);
  and (_09602_, _09566_, word_in[25]);
  or (_08314_, _09602_, _09601_);
  or (_09603_, _09571_, _08707_);
  not (_09604_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_09605_, _09574_, _09604_);
  and (_09606_, _09574_, _08572_);
  or (_09607_, _09606_, _09605_);
  or (_09608_, _09607_, _09573_);
  not (_09609_, _09573_);
  or (_09610_, _09609_, word_in[10]);
  and (_09611_, _09610_, _09608_);
  or (_09612_, _09611_, _09568_);
  and (_09613_, _09612_, _09603_);
  or (_09614_, _09613_, _09566_);
  or (_09615_, _09567_, word_in[26]);
  and (_08317_, _09615_, _09614_);
  and (_09616_, _09574_, _08586_);
  not (_09617_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_09618_, _09574_, _09617_);
  nor (_09619_, _09618_, _09616_);
  nor (_09620_, _09619_, _09573_);
  and (_09621_, _09573_, word_in[11]);
  or (_09622_, _09621_, _09620_);
  and (_09623_, _09622_, _09571_);
  and (_09624_, _09568_, _08712_);
  or (_09625_, _09624_, _09566_);
  or (_09626_, _09625_, _09623_);
  or (_09627_, _09567_, word_in[27]);
  and (_08321_, _09627_, _09626_);
  not (_09628_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_09629_, _09574_, _09628_);
  and (_09630_, _09574_, _08598_);
  or (_09631_, _09630_, _09629_);
  or (_09632_, _09631_, _09573_);
  or (_09633_, _09609_, word_in[12]);
  and (_09634_, _09633_, _09632_);
  or (_09635_, _09634_, _09568_);
  or (_09636_, _09571_, _08733_);
  and (_09637_, _09636_, _09567_);
  and (_09638_, _09637_, _09635_);
  and (_09639_, _09566_, word_in[28]);
  or (_08325_, _09639_, _09638_);
  not (_09640_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_09641_, _09574_, _09640_);
  and (_09642_, _09574_, _08612_);
  or (_09643_, _09642_, _09641_);
  or (_09644_, _09643_, _09573_);
  or (_09645_, _09609_, word_in[13]);
  and (_09646_, _09645_, _09644_);
  or (_09647_, _09646_, _09568_);
  or (_09648_, _09571_, _08746_);
  and (_09649_, _09648_, _09567_);
  and (_09650_, _09649_, _09647_);
  and (_09651_, _09566_, word_in[29]);
  or (_08329_, _09651_, _09650_);
  not (_09652_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_09653_, _09574_, _09652_);
  and (_09654_, _09574_, _08628_);
  or (_09655_, _09654_, _09653_);
  or (_09656_, _09655_, _09573_);
  nand (_09657_, _09573_, _09418_);
  and (_09658_, _09657_, _09656_);
  or (_09659_, _09658_, _09568_);
  or (_09660_, _09571_, _08759_);
  and (_09661_, _09660_, _09659_);
  or (_09662_, _09661_, _09566_);
  or (_09663_, _09567_, word_in[30]);
  and (_08331_, _09663_, _09662_);
  or (_09664_, _09571_, _08037_);
  nor (_09665_, _09574_, _07722_);
  and (_09666_, _09574_, _08029_);
  or (_09667_, _09666_, _09665_);
  or (_09668_, _09667_, _09573_);
  nand (_09669_, _09573_, _08642_);
  and (_09670_, _09669_, _09668_);
  or (_09671_, _09670_, _09568_);
  and (_09672_, _09671_, _09664_);
  or (_09673_, _09672_, _09566_);
  or (_09674_, _09567_, word_in[31]);
  and (_08335_, _09674_, _09673_);
  and (_09675_, _09460_, _07765_);
  and (_09676_, _08778_, _07889_);
  not (_09677_, _09676_);
  or (_09678_, _09677_, _08544_);
  and (_09679_, _08782_, _07783_);
  not (_09680_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_09681_, _09470_, _08786_);
  nor (_09682_, _09681_, _09680_);
  and (_09683_, _09681_, _08666_);
  or (_09684_, _09683_, _09682_);
  or (_09685_, _09684_, _09679_);
  not (_09686_, _09679_);
  or (_09687_, _09686_, word_in[8]);
  and (_09688_, _09687_, _09685_);
  or (_09690_, _09688_, _09676_);
  and (_09691_, _09690_, _09678_);
  or (_09692_, _09691_, _09675_);
  not (_09693_, _09675_);
  or (_09694_, _09693_, word_in[24]);
  and (_08400_, _09694_, _09692_);
  not (_09695_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_09696_, _09681_, _09695_);
  and (_09697_, _09681_, _08556_);
  or (_09698_, _09697_, _09696_);
  or (_09699_, _09698_, _09679_);
  or (_09700_, _09686_, word_in[9]);
  and (_09701_, _09700_, _09699_);
  or (_09702_, _09701_, _09676_);
  or (_09703_, _09677_, _08694_);
  and (_09704_, _09703_, _09693_);
  and (_09705_, _09704_, _09702_);
  and (_09706_, _09675_, word_in[25]);
  or (_08403_, _09706_, _09705_);
  or (_09707_, _09677_, _08707_);
  not (_09708_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_09709_, _09681_, _09708_);
  and (_09710_, _09681_, _08572_);
  or (_09711_, _09710_, _09709_);
  or (_09712_, _09711_, _09679_);
  or (_09713_, _09686_, word_in[10]);
  and (_09714_, _09713_, _09712_);
  or (_09715_, _09714_, _09676_);
  and (_09716_, _09715_, _09707_);
  or (_09717_, _09716_, _09675_);
  or (_09718_, _09693_, word_in[26]);
  and (_08407_, _09718_, _09717_);
  or (_09719_, _09677_, _08712_);
  not (_09720_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_09721_, _09681_, _09720_);
  and (_09722_, _09681_, _08586_);
  or (_09723_, _09722_, _09721_);
  or (_09724_, _09723_, _09679_);
  or (_09725_, _09686_, word_in[11]);
  and (_09726_, _09725_, _09724_);
  or (_09727_, _09726_, _09676_);
  and (_09728_, _09727_, _09719_);
  or (_09729_, _09728_, _09675_);
  or (_09730_, _09693_, word_in[27]);
  and (_08410_, _09730_, _09729_);
  not (_09731_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_09732_, _09681_, _09731_);
  and (_09733_, _09681_, _08598_);
  or (_09734_, _09733_, _09732_);
  or (_09735_, _09734_, _09679_);
  or (_09736_, _09686_, word_in[12]);
  and (_09737_, _09736_, _09735_);
  or (_09738_, _09737_, _09676_);
  or (_09739_, _09677_, _08733_);
  and (_09740_, _09739_, _09693_);
  and (_09741_, _09740_, _09738_);
  and (_09742_, _09675_, word_in[28]);
  or (_08413_, _09742_, _09741_);
  or (_09743_, _09677_, _08746_);
  not (_09744_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_09745_, _09681_, _09744_);
  and (_09746_, _09681_, _08612_);
  or (_09747_, _09746_, _09745_);
  or (_09748_, _09747_, _09679_);
  or (_09749_, _09686_, word_in[13]);
  and (_09750_, _09749_, _09748_);
  or (_09751_, _09750_, _09676_);
  and (_09752_, _09751_, _09743_);
  or (_09753_, _09752_, _09675_);
  or (_09754_, _09693_, word_in[29]);
  and (_08416_, _09754_, _09753_);
  or (_09755_, _09677_, _08759_);
  not (_09756_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_09757_, _09681_, _09756_);
  and (_09758_, _09681_, _08628_);
  or (_09759_, _09758_, _09757_);
  or (_09760_, _09759_, _09679_);
  nand (_09761_, _09679_, _09418_);
  and (_09762_, _09761_, _09760_);
  or (_09763_, _09762_, _09676_);
  and (_09764_, _09763_, _09755_);
  and (_09765_, _09764_, _09693_);
  and (_09766_, _09675_, word_in[30]);
  or (_08419_, _09766_, _09765_);
  nor (_09767_, _09681_, _07822_);
  and (_09768_, _09681_, _08029_);
  or (_09769_, _09768_, _09767_);
  or (_09770_, _09769_, _09679_);
  nand (_09771_, _09679_, _08642_);
  and (_09772_, _09771_, _09770_);
  or (_09773_, _09772_, _09676_);
  or (_09774_, _09677_, _08037_);
  and (_09775_, _09774_, _09693_);
  and (_09776_, _09775_, _09773_);
  and (_09777_, _09675_, word_in[31]);
  or (_08421_, _09777_, _09776_);
  and (_09778_, _06703_, _05277_);
  not (_09779_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_09780_, _05277_, _09779_);
  or (_09781_, _09780_, _05572_);
  or (_09782_, _09781_, _09778_);
  or (_09783_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_09784_, _09783_, _05141_);
  and (_08473_, _09784_, _09782_);
  not (_09785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  or (_09786_, _06695_, _09785_);
  or (_09787_, _06697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_09788_, _09787_, _05141_);
  and (_08477_, _09788_, _09786_);
  and (_09789_, _08917_, _07889_);
  and (_09790_, _08022_, _07783_);
  and (_09791_, _09790_, word_in[8]);
  and (_09792_, _09470_, _08025_);
  and (_09793_, _09792_, _08666_);
  not (_09794_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor (_09795_, _09792_, _09794_);
  nor (_09796_, _09795_, _09793_);
  nor (_09797_, _09796_, _09790_);
  or (_09798_, _09797_, _09791_);
  or (_09799_, _09798_, _09789_);
  and (_09800_, _09460_, _07761_);
  not (_09801_, _09789_);
  nor (_09802_, _09801_, _08544_);
  nor (_09803_, _09802_, _09800_);
  and (_09804_, _09803_, _09799_);
  and (_09805_, _09800_, word_in[24]);
  or (_08486_, _09805_, _09804_);
  not (_09806_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_09807_, _09792_, _09806_);
  and (_09808_, _09792_, _08556_);
  or (_09809_, _09808_, _09807_);
  or (_09810_, _09809_, _09790_);
  not (_09811_, _09790_);
  or (_09812_, _09811_, word_in[9]);
  and (_09813_, _09812_, _09810_);
  or (_09814_, _09813_, _09789_);
  not (_09815_, _09800_);
  or (_09816_, _09801_, _08694_);
  and (_09817_, _09816_, _09815_);
  and (_09818_, _09817_, _09814_);
  and (_09819_, _09800_, _08566_);
  or (_08490_, _09819_, _09818_);
  not (_09820_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_09821_, _09792_, _09820_);
  and (_09822_, _09792_, _08572_);
  or (_09823_, _09822_, _09821_);
  or (_09824_, _09823_, _09790_);
  or (_09825_, _09811_, word_in[10]);
  and (_09826_, _09825_, _09824_);
  or (_09827_, _09826_, _09789_);
  or (_09828_, _09801_, _08707_);
  and (_09829_, _09828_, _09815_);
  and (_09830_, _09829_, _09827_);
  and (_09831_, _09800_, _08568_);
  or (_08493_, _09831_, _09830_);
  not (_09832_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_09834_, _09792_, _09832_);
  and (_09835_, _09792_, _08586_);
  or (_09836_, _09835_, _09834_);
  or (_09837_, _09836_, _09790_);
  or (_09838_, _09811_, word_in[11]);
  and (_09839_, _09838_, _09837_);
  or (_09840_, _09839_, _09789_);
  or (_09841_, _09801_, _08712_);
  and (_09842_, _09841_, _09815_);
  and (_09843_, _09842_, _09840_);
  and (_09844_, _09800_, _08582_);
  or (_08495_, _09844_, _09843_);
  not (_09845_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_09846_, _09792_, _09845_);
  and (_09847_, _09792_, _08598_);
  or (_09848_, _09847_, _09846_);
  or (_09849_, _09848_, _09790_);
  or (_09850_, _09811_, word_in[12]);
  and (_09851_, _09850_, _09849_);
  or (_09852_, _09851_, _09789_);
  or (_09853_, _09801_, _08733_);
  and (_09854_, _09853_, _09815_);
  and (_09856_, _09854_, _09852_);
  and (_09857_, _09800_, _08608_);
  or (_08498_, _09857_, _09856_);
  not (_09858_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_09860_, _09792_, _09858_);
  and (_09861_, _09792_, _08612_);
  or (_09863_, _09861_, _09860_);
  or (_09864_, _09863_, _09790_);
  or (_09865_, _09811_, word_in[13]);
  and (_09866_, _09865_, _09864_);
  or (_09867_, _09866_, _09789_);
  or (_09868_, _09801_, _08746_);
  and (_09869_, _09868_, _09815_);
  and (_09870_, _09869_, _09867_);
  and (_09871_, _09800_, _08622_);
  or (_08502_, _09871_, _09870_);
  not (_09872_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_09873_, _09792_, _09872_);
  and (_09874_, _09792_, _08628_);
  or (_09875_, _09874_, _09873_);
  or (_09876_, _09875_, _09790_);
  nand (_09877_, _09790_, _09418_);
  and (_09878_, _09877_, _09876_);
  or (_09879_, _09878_, _09789_);
  or (_09880_, _09801_, _08759_);
  and (_09881_, _09880_, _09815_);
  and (_09882_, _09881_, _09879_);
  and (_09883_, _09800_, _08624_);
  or (_08506_, _09883_, _09882_);
  nor (_09884_, _09792_, _07711_);
  and (_09885_, _09792_, _08029_);
  or (_09886_, _09885_, _09884_);
  or (_09887_, _09886_, _09790_);
  nand (_09888_, _09790_, _08642_);
  and (_09889_, _09888_, _09887_);
  or (_09890_, _09889_, _09789_);
  or (_09891_, _09801_, _08037_);
  and (_09892_, _09891_, _09815_);
  and (_09893_, _09892_, _09890_);
  and (_09894_, _09800_, _08011_);
  or (_08510_, _09894_, _09893_);
  and (_09895_, _08382_, _05522_);
  and (_09896_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_09897_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_09898_, _09897_, _09896_);
  nor (_09899_, _09898_, _08243_);
  and (_09900_, _08396_, _06290_);
  or (_09901_, _09900_, _09899_);
  or (_09902_, _09901_, _09895_);
  and (_08517_, _09902_, _05141_);
  and (_09903_, _08018_, _07798_);
  not (_09904_, _09903_);
  and (_09905_, _08021_, _08254_);
  not (_09906_, _09905_);
  or (_09907_, _09906_, word_in[8]);
  not (_09908_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_09909_, _08531_, _08027_);
  nor (_09910_, _09909_, _09908_);
  and (_09911_, _09909_, word_in[0]);
  or (_09912_, _09911_, _09910_);
  or (_09913_, _09912_, _09905_);
  and (_09914_, _09913_, _09907_);
  and (_09915_, _09914_, _09904_);
  not (_09916_, _07946_);
  and (_09917_, _09034_, _09916_);
  and (_09918_, _09917_, _07788_);
  and (_09919_, _09903_, _08544_);
  or (_09920_, _09919_, _09918_);
  or (_09921_, _09920_, _09915_);
  not (_09922_, _09918_);
  or (_09923_, _09922_, _09040_);
  and (_13475_, _09923_, _09921_);
  not (_09924_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_09925_, _09909_, _09924_);
  and (_09926_, _09909_, word_in[1]);
  or (_09927_, _09926_, _09925_);
  and (_09928_, _09927_, _09906_);
  and (_09929_, _09905_, word_in[9]);
  or (_09930_, _09929_, _09928_);
  and (_09931_, _09930_, _09904_);
  and (_09932_, _09903_, _08694_);
  or (_09933_, _09932_, _09918_);
  or (_09934_, _09933_, _09931_);
  or (_09935_, _09922_, _08566_);
  and (_13476_, _09935_, _09934_);
  not (_09936_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_09937_, _09909_, _09936_);
  and (_09938_, _09909_, word_in[2]);
  or (_09939_, _09938_, _09937_);
  and (_09940_, _09939_, _09906_);
  and (_09941_, _09905_, word_in[10]);
  or (_09942_, _09941_, _09940_);
  and (_09943_, _09942_, _09904_);
  and (_09944_, _09903_, _08707_);
  or (_09945_, _09944_, _09918_);
  or (_09946_, _09945_, _09943_);
  or (_09947_, _09922_, _08568_);
  and (_13477_, _09947_, _09946_);
  not (_09948_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_09949_, _09909_, _09948_);
  and (_09950_, _09909_, word_in[3]);
  or (_09951_, _09950_, _09949_);
  and (_09952_, _09951_, _09906_);
  and (_09953_, _09905_, word_in[11]);
  or (_09954_, _09953_, _09952_);
  and (_09955_, _09954_, _09904_);
  and (_09956_, _09903_, _08712_);
  or (_09957_, _09956_, _09918_);
  or (_09958_, _09957_, _09955_);
  or (_09959_, _09922_, _08582_);
  and (_13478_, _09959_, _09958_);
  not (_09960_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_09961_, _09909_, _09960_);
  and (_09962_, _09909_, word_in[4]);
  or (_09963_, _09962_, _09961_);
  and (_09964_, _09963_, _09906_);
  and (_09965_, _09905_, word_in[12]);
  or (_09966_, _09965_, _09964_);
  and (_09967_, _09966_, _09904_);
  and (_09968_, _09903_, _08733_);
  or (_09969_, _09968_, _09918_);
  or (_09970_, _09969_, _09967_);
  or (_09971_, _09922_, _08608_);
  and (_13479_, _09971_, _09970_);
  not (_09972_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_09973_, _09909_, _09972_);
  and (_09974_, _09909_, word_in[5]);
  or (_09975_, _09974_, _09973_);
  or (_09976_, _09975_, _09905_);
  or (_09977_, _09906_, word_in[13]);
  and (_09978_, _09977_, _09976_);
  and (_09979_, _09978_, _09904_);
  and (_09980_, _09903_, _08746_);
  or (_09981_, _09980_, _09918_);
  or (_09982_, _09981_, _09979_);
  or (_09983_, _09922_, _08622_);
  and (_13480_, _09983_, _09982_);
  not (_09984_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_09985_, _09909_, _09984_);
  and (_09986_, _09909_, word_in[6]);
  or (_09987_, _09986_, _09985_);
  and (_09988_, _09987_, _09906_);
  and (_09989_, _09905_, word_in[14]);
  or (_09990_, _09989_, _09988_);
  and (_09991_, _09990_, _09904_);
  and (_09992_, _09903_, _08759_);
  or (_09993_, _09992_, _09918_);
  or (_09994_, _09993_, _09991_);
  or (_09995_, _09922_, _08624_);
  and (_13481_, _09995_, _09994_);
  nor (_09996_, _09909_, _07864_);
  and (_09997_, _09909_, word_in[7]);
  or (_09998_, _09997_, _09996_);
  and (_09999_, _09998_, _09906_);
  and (_10000_, _09905_, word_in[15]);
  or (_10001_, _10000_, _09999_);
  and (_10002_, _10001_, _09904_);
  and (_10003_, _09903_, _08037_);
  or (_10004_, _10003_, _09918_);
  or (_10005_, _10004_, _10002_);
  or (_10006_, _09922_, _08011_);
  and (_13482_, _10006_, _10005_);
  and (_10007_, _09917_, _07798_);
  and (_10008_, _08018_, _07765_);
  and (_10009_, _08664_, _07811_);
  not (_10010_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_10011_, _08668_, _08027_);
  nor (_10012_, _10011_, _10010_);
  and (_10013_, _10011_, _08666_);
  or (_10014_, _10013_, _10012_);
  or (_10015_, _10014_, _10009_);
  not (_10016_, word_in[8]);
  nand (_10017_, _10009_, _10016_);
  and (_10018_, _10017_, _10015_);
  or (_10019_, _10018_, _10008_);
  not (_10020_, _10008_);
  or (_10021_, _10020_, _08544_);
  and (_10022_, _10021_, _10019_);
  or (_10023_, _10022_, _10007_);
  not (_10024_, _10007_);
  or (_10025_, _10024_, word_in[24]);
  and (_13483_, _10025_, _10023_);
  not (_10026_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_10027_, _10011_, _10026_);
  and (_10028_, _10011_, _08556_);
  nor (_10029_, _10028_, _10027_);
  nor (_10030_, _10029_, _10009_);
  and (_10031_, _10009_, word_in[9]);
  or (_10032_, _10031_, _10030_);
  and (_10033_, _10032_, _10020_);
  and (_10034_, _10008_, _08694_);
  or (_10035_, _10034_, _10007_);
  or (_10036_, _10035_, _10033_);
  or (_10037_, _10024_, word_in[25]);
  and (_13484_, _10037_, _10036_);
  not (_10038_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_10039_, _10011_, _10038_);
  and (_10040_, _10011_, _08572_);
  nor (_10041_, _10040_, _10039_);
  nor (_10042_, _10041_, _10009_);
  and (_10043_, _10009_, word_in[10]);
  or (_10044_, _10043_, _10042_);
  and (_10045_, _10044_, _10020_);
  and (_10046_, _10008_, _08707_);
  or (_10047_, _10046_, _10007_);
  or (_10048_, _10047_, _10045_);
  or (_10049_, _10024_, word_in[26]);
  and (_13485_, _10049_, _10048_);
  not (_10050_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_10051_, _10011_, _10050_);
  and (_10052_, _10011_, _08586_);
  nor (_10053_, _10052_, _10051_);
  nor (_10054_, _10053_, _10009_);
  and (_10055_, _10009_, word_in[11]);
  or (_10056_, _10055_, _10054_);
  and (_10057_, _10056_, _10020_);
  and (_10058_, _10008_, _08712_);
  or (_10059_, _10058_, _10007_);
  or (_10060_, _10059_, _10057_);
  or (_10061_, _10024_, word_in[27]);
  and (_08679_, _10061_, _10060_);
  and (_10062_, _08382_, _06290_);
  and (_10063_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_10064_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_10065_, _10064_, _10063_);
  nor (_10066_, _10065_, _08243_);
  and (_10067_, _08396_, _05561_);
  or (_10069_, _10067_, _10066_);
  or (_10070_, _10069_, _10062_);
  and (_08682_, _10070_, _05141_);
  not (_10071_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_10073_, _10011_, _10071_);
  and (_10074_, _10011_, _08598_);
  nor (_10075_, _10074_, _10073_);
  nor (_10076_, _10075_, _10009_);
  and (_10077_, _10009_, word_in[12]);
  or (_10078_, _10077_, _10076_);
  and (_10079_, _10078_, _10020_);
  and (_10080_, _10008_, _08733_);
  or (_10081_, _10080_, _10007_);
  or (_10082_, _10081_, _10079_);
  or (_10083_, _10024_, word_in[28]);
  and (_13486_, _10083_, _10082_);
  not (_10084_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_10085_, _10011_, _10084_);
  and (_10086_, _10011_, _08612_);
  nor (_10087_, _10086_, _10085_);
  nor (_10088_, _10087_, _10009_);
  and (_10089_, _10009_, word_in[13]);
  or (_10090_, _10089_, _10088_);
  and (_10091_, _10090_, _10020_);
  and (_10092_, _10008_, _08746_);
  or (_10093_, _10092_, _10007_);
  or (_10094_, _10093_, _10091_);
  or (_10095_, _10024_, word_in[29]);
  and (_13487_, _10095_, _10094_);
  not (_10096_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_10097_, _10011_, _10096_);
  and (_10098_, _10011_, _08628_);
  nor (_10099_, _10098_, _10097_);
  nor (_10100_, _10099_, _10009_);
  and (_10101_, _10009_, word_in[14]);
  or (_10102_, _10101_, _10100_);
  and (_10103_, _10102_, _10020_);
  and (_10104_, _10008_, _08759_);
  or (_10105_, _10104_, _10007_);
  or (_10106_, _10105_, _10103_);
  or (_10107_, _10024_, word_in[30]);
  and (_13488_, _10107_, _10106_);
  and (_10108_, _08382_, _06283_);
  and (_10109_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_10110_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_10111_, _10110_, _10109_);
  nor (_10112_, _10111_, _08243_);
  and (_10113_, _08396_, _06004_);
  or (_10114_, _10113_, _10112_);
  or (_10116_, _10114_, _10108_);
  and (_08691_, _10116_, _05141_);
  nor (_10117_, _10011_, _07717_);
  and (_10118_, _10011_, _08029_);
  nor (_10119_, _10118_, _10117_);
  nor (_10120_, _10119_, _10009_);
  and (_10121_, _10009_, word_in[15]);
  or (_10122_, _10121_, _10120_);
  and (_10123_, _10122_, _10020_);
  and (_10124_, _10008_, _08037_);
  or (_10125_, _10124_, _10007_);
  or (_10126_, _10125_, _10123_);
  or (_10127_, _10024_, word_in[31]);
  and (_13489_, _10127_, _10126_);
  and (_10128_, _09917_, _07765_);
  and (_10129_, _08018_, _07761_);
  and (_10130_, _08782_, _07811_);
  not (_10131_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_10132_, _08786_, _08008_);
  nor (_10133_, _10132_, _10131_);
  and (_10134_, _10132_, _08666_);
  or (_10135_, _10134_, _10133_);
  or (_10136_, _10135_, _10130_);
  nand (_10137_, _10130_, _10016_);
  and (_10138_, _10137_, _10136_);
  or (_10139_, _10138_, _10129_);
  not (_10140_, _10129_);
  or (_10141_, _10140_, _08544_);
  and (_10142_, _10141_, _10139_);
  or (_10143_, _10142_, _10128_);
  not (_10144_, _10128_);
  or (_10145_, _10144_, word_in[24]);
  and (_08770_, _10145_, _10143_);
  not (_10146_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_10147_, _10132_, _10146_);
  and (_10148_, _10132_, _08556_);
  nor (_10149_, _10148_, _10147_);
  nor (_10150_, _10149_, _10130_);
  and (_10151_, _10130_, word_in[9]);
  or (_10152_, _10151_, _10150_);
  and (_10154_, _10152_, _10140_);
  and (_10155_, _10129_, _08694_);
  or (_10156_, _10155_, _10128_);
  or (_10157_, _10156_, _10154_);
  or (_10158_, _10144_, word_in[25]);
  and (_08775_, _10158_, _10157_);
  not (_10159_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_10160_, _10132_, _10159_);
  and (_10161_, _10132_, _08572_);
  or (_10162_, _10161_, _10160_);
  or (_10163_, _10162_, _10130_);
  not (_10164_, _10130_);
  or (_10165_, _10164_, word_in[10]);
  and (_10166_, _10165_, _10163_);
  or (_10167_, _10166_, _10129_);
  or (_10168_, _10140_, _08707_);
  and (_10169_, _10168_, _10144_);
  and (_10170_, _10169_, _10167_);
  and (_10171_, _10128_, word_in[26]);
  or (_08777_, _10171_, _10170_);
  not (_10172_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_10173_, _10132_, _10172_);
  and (_10174_, _10132_, _08586_);
  nor (_10175_, _10174_, _10173_);
  nor (_10176_, _10175_, _10130_);
  and (_10177_, _10130_, word_in[11]);
  or (_10178_, _10177_, _10176_);
  and (_10179_, _10178_, _10140_);
  and (_10180_, _10129_, _08712_);
  or (_10181_, _10180_, _10128_);
  or (_10182_, _10181_, _10179_);
  or (_10183_, _10144_, word_in[27]);
  and (_08781_, _10183_, _10182_);
  not (_10184_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_10185_, _10132_, _10184_);
  and (_10186_, _10132_, _08598_);
  nor (_10187_, _10186_, _10185_);
  nor (_10188_, _10187_, _10130_);
  and (_10189_, _10130_, word_in[12]);
  or (_10190_, _10189_, _10188_);
  and (_10192_, _10190_, _10140_);
  and (_10193_, _10129_, _08733_);
  or (_10194_, _10193_, _10128_);
  or (_10195_, _10194_, _10192_);
  or (_10196_, _10144_, word_in[28]);
  and (_08785_, _10196_, _10195_);
  not (_10197_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_10198_, _10132_, _10197_);
  and (_10199_, _10132_, _08612_);
  nor (_10200_, _10199_, _10198_);
  nor (_10201_, _10200_, _10130_);
  and (_10202_, _10130_, word_in[13]);
  or (_10203_, _10202_, _10201_);
  and (_10204_, _10203_, _10140_);
  and (_10205_, _10129_, _08746_);
  or (_10206_, _10205_, _10128_);
  or (_10207_, _10206_, _10204_);
  or (_10208_, _10144_, word_in[29]);
  and (_08788_, _10208_, _10207_);
  not (_10209_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_10210_, _10132_, _10209_);
  and (_10211_, _10132_, _08628_);
  nor (_10212_, _10211_, _10210_);
  nor (_10213_, _10212_, _10130_);
  and (_10214_, _10130_, word_in[14]);
  or (_10215_, _10214_, _10213_);
  and (_10216_, _10215_, _10140_);
  and (_10217_, _10129_, _08759_);
  or (_10218_, _10217_, _10128_);
  or (_10219_, _10218_, _10216_);
  or (_10220_, _10144_, word_in[30]);
  and (_08792_, _10220_, _10219_);
  nor (_10221_, _10132_, _07858_);
  and (_10222_, _10132_, _08029_);
  nor (_10223_, _10222_, _10221_);
  nor (_10224_, _10223_, _10130_);
  and (_10225_, _10130_, word_in[15]);
  or (_10226_, _10225_, _10224_);
  and (_10227_, _10226_, _10140_);
  and (_10228_, _10129_, _08037_);
  or (_10229_, _10228_, _10128_);
  or (_10230_, _10229_, _10227_);
  or (_10231_, _10144_, word_in[31]);
  and (_08796_, _10231_, _10230_);
  and (_10232_, _09040_, _08013_);
  and (_10233_, _08028_, word_in[0]);
  not (_10234_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_10235_, _08028_, _10234_);
  nor (_10237_, _10235_, _10233_);
  nor (_10238_, _10237_, _08023_);
  and (_10240_, _08023_, word_in[8]);
  or (_10241_, _10240_, _10238_);
  and (_10242_, _10241_, _08020_);
  and (_10243_, _08544_, _08019_);
  or (_10244_, _10243_, _10242_);
  and (_10246_, _10244_, _08015_);
  or (_08867_, _10246_, _10232_);
  and (_10247_, _08566_, _08013_);
  not (_10248_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_10249_, _08028_, _10248_);
  and (_10250_, _08028_, word_in[1]);
  nor (_10252_, _10250_, _10249_);
  nor (_10253_, _10252_, _08023_);
  and (_10254_, _08023_, word_in[9]);
  or (_10255_, _10254_, _10253_);
  and (_10256_, _10255_, _08020_);
  and (_10257_, _08694_, _08019_);
  or (_10258_, _10257_, _10256_);
  and (_10259_, _10258_, _08015_);
  or (_08870_, _10259_, _10247_);
  not (_10260_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_10261_, _08028_, _10260_);
  and (_10262_, _08028_, word_in[2]);
  nor (_10263_, _10262_, _10261_);
  nor (_10264_, _10263_, _08023_);
  and (_10265_, _08023_, word_in[10]);
  or (_10266_, _10265_, _10264_);
  and (_10267_, _10266_, _08020_);
  and (_10268_, _08707_, _08019_);
  or (_10269_, _10268_, _08013_);
  or (_10270_, _10269_, _10267_);
  or (_10271_, _08015_, word_in[26]);
  and (_08873_, _10271_, _10270_);
  not (_10272_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_10273_, _08028_, _10272_);
  and (_10274_, _08028_, word_in[3]);
  nor (_10275_, _10274_, _10273_);
  nor (_10276_, _10275_, _08023_);
  and (_10277_, _08023_, word_in[11]);
  or (_10278_, _10277_, _10276_);
  and (_10279_, _10278_, _08020_);
  and (_10280_, _08712_, _08019_);
  or (_10281_, _10280_, _08013_);
  or (_10282_, _10281_, _10279_);
  or (_10283_, _08015_, word_in[27]);
  and (_08877_, _10283_, _10282_);
  and (_10284_, _08608_, _08013_);
  and (_10285_, _08028_, word_in[4]);
  not (_10286_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_10287_, _08028_, _10286_);
  nor (_10288_, _10287_, _10285_);
  nor (_10289_, _10288_, _08023_);
  and (_10290_, _08023_, word_in[12]);
  or (_10291_, _10290_, _10289_);
  and (_10292_, _10291_, _08020_);
  and (_10293_, _08733_, _08019_);
  or (_10294_, _10293_, _10292_);
  and (_10295_, _10294_, _08015_);
  or (_08879_, _10295_, _10284_);
  and (_10296_, _08622_, _08013_);
  and (_10297_, _08028_, word_in[5]);
  not (_10298_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_10299_, _08028_, _10298_);
  nor (_10300_, _10299_, _10297_);
  nor (_10301_, _10300_, _08023_);
  and (_10302_, _08023_, word_in[13]);
  or (_10303_, _10302_, _10301_);
  and (_10304_, _10303_, _08020_);
  and (_10305_, _08746_, _08019_);
  or (_10306_, _10305_, _10304_);
  and (_10307_, _10306_, _08015_);
  or (_08882_, _10307_, _10296_);
  and (_10308_, _08624_, _08013_);
  not (_10309_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_10310_, _08028_, _10309_);
  and (_10311_, _08028_, word_in[6]);
  nor (_10312_, _10311_, _10310_);
  nor (_10313_, _10312_, _08023_);
  and (_10314_, _08023_, word_in[14]);
  or (_10315_, _10314_, _10313_);
  and (_10316_, _10315_, _08020_);
  and (_10317_, _08759_, _08019_);
  or (_10318_, _10317_, _10316_);
  and (_10320_, _10318_, _08015_);
  or (_08887_, _10320_, _10308_);
  or (_08889_, _06811_, _06831_);
  or (_10321_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand (_10322_, _07619_, _06324_);
  and (_10323_, _10322_, _05141_);
  and (_08991_, _10323_, _10321_);
  and (_10324_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_10325_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_09143_, _10325_, _10324_);
  or (_10326_, _05842_, _05840_);
  not (_10327_, _05686_);
  nand (_10328_, _05840_, _10327_);
  and (_10329_, _10328_, _05656_);
  and (_10330_, _10329_, _10326_);
  and (_10331_, _06600_, ABINPUT000000[0]);
  and (_10332_, _06606_, ABINPUT000[0]);
  or (_10333_, _10332_, _10331_);
  nand (_10334_, _05879_, _05846_);
  and (_10335_, _05880_, _05844_);
  and (_10336_, _10335_, _10334_);
  or (_10337_, _10336_, _10333_);
  or (_10338_, _10337_, _10330_);
  and (_10339_, _10338_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_10341_, _05256_);
  and (_10342_, _06877_, _10341_);
  and (_10343_, _05266_, _05228_);
  and (_10345_, _10343_, _05647_);
  and (_10346_, _10345_, _10342_);
  not (_10348_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_10349_, _10348_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_10350_, _10349_, _10346_);
  or (_10351_, _10350_, _10339_);
  and (_10352_, _06018_, _05210_);
  and (_10353_, _06733_, _05281_);
  and (_10354_, _10353_, _10352_);
  not (_10355_, _10354_);
  and (_10356_, _05922_, _06620_);
  not (_10357_, _06620_);
  nand (_10358_, _10357_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand (_10359_, _10358_, _10346_);
  or (_10360_, _10359_, _10356_);
  and (_10361_, _10360_, _10355_);
  and (_10362_, _10361_, _10351_);
  nor (_10363_, _10355_, _05560_);
  or (_10364_, _10363_, _10362_);
  and (_09170_, _10364_, _05141_);
  and (_10365_, _10352_, _06733_);
  and (_10366_, _10365_, _05281_);
  and (_10367_, _10346_, _05288_);
  nand (_10368_, _10367_, _05963_);
  or (_10369_, _10367_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_10370_, _10369_, _10368_);
  or (_10371_, _10370_, _10366_);
  nand (_10372_, _10354_, _06178_);
  and (_10373_, _10372_, _05141_);
  and (_09173_, _10373_, _10371_);
  nor (_10374_, _05209_, _06007_);
  nor (_10375_, _10374_, _08469_);
  not (_10376_, _10346_);
  or (_10378_, _10376_, _10375_);
  and (_10379_, _10378_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_10380_, _05922_, _08469_);
  and (_10381_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_10383_, _10381_, _10380_);
  and (_10384_, _10383_, _10346_);
  or (_10385_, _10384_, _10379_);
  and (_10386_, _10385_, _10355_);
  and (_10387_, _10354_, _05522_);
  or (_10389_, _10387_, _10386_);
  and (_09564_, _10389_, _05141_);
  and (_10390_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_10391_, _05864_, _05844_);
  and (_10392_, _05835_, _05656_);
  or (_10393_, _10392_, _10391_);
  and (_10394_, _10393_, _10390_);
  nand (_10395_, _10390_, _06598_);
  and (_10396_, _10395_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_10397_, _10396_, _10346_);
  or (_10398_, _10397_, _10394_);
  or (_10399_, _06207_, _07328_);
  nand (_10400_, _10399_, _10346_);
  or (_10401_, _10400_, _06208_);
  and (_10402_, _10401_, _10398_);
  or (_10403_, _10402_, _10354_);
  nand (_10404_, _10354_, _06244_);
  and (_10405_, _10404_, _05141_);
  and (_09569_, _10405_, _10403_);
  and (_10407_, _05275_, _06007_);
  and (_10408_, _10346_, _10407_);
  nand (_10410_, _10408_, _05963_);
  or (_10411_, _10408_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_10413_, _10411_, _10410_);
  or (_10414_, _10413_, _10366_);
  or (_10415_, _10355_, _06004_);
  and (_10416_, _10415_, _05141_);
  and (_09572_, _10416_, _10414_);
  or (_10418_, _06389_, _07117_);
  or (_10419_, _06270_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_10420_, _10419_, _05141_);
  and (_09689_, _10420_, _10418_);
  and (_10421_, _07758_, word_in[0]);
  nand (_10422_, _07613_, _09576_);
  or (_10423_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_10424_, _10423_, _10422_);
  and (_10425_, _10424_, _07666_);
  nand (_10426_, _07613_, _09794_);
  or (_10427_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_10428_, _10427_, _10426_);
  and (_10429_, _10428_, _07643_);
  nand (_10430_, _07613_, _10010_);
  or (_10431_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_10432_, _10431_, _10430_);
  and (_10433_, _10432_, _07640_);
  or (_10434_, _10433_, _10429_);
  or (_10435_, _10434_, _10425_);
  nand (_10436_, _07613_, _10234_);
  or (_10438_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_10439_, _10438_, _10436_);
  and (_10440_, _10439_, _07650_);
  or (_10441_, _10440_, _07676_);
  or (_10442_, _10441_, _10435_);
  nand (_10443_, _07613_, _08672_);
  or (_10444_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_10445_, _10444_, _10443_);
  and (_10446_, _10445_, _07666_);
  nand (_10447_, _07613_, _08924_);
  or (_10448_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_10449_, _10448_, _10447_);
  and (_10450_, _10449_, _07643_);
  nand (_10451_, _07613_, _09133_);
  or (_10452_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_10453_, _10452_, _10451_);
  and (_10454_, _10453_, _07640_);
  or (_10455_, _10454_, _10450_);
  or (_10456_, _10455_, _10446_);
  nand (_10457_, _07613_, _09343_);
  or (_10459_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_10460_, _10459_, _10457_);
  and (_10462_, _10460_, _07650_);
  or (_10463_, _10462_, _07626_);
  or (_10464_, _10463_, _10456_);
  and (_10465_, _10464_, _10442_);
  and (_10466_, _10465_, _07705_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _10466_, _10421_);
  and (_10467_, _07758_, word_in[1]);
  nand (_10468_, _07613_, _09592_);
  or (_10469_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_10470_, _10469_, _10468_);
  and (_10471_, _10470_, _07666_);
  nand (_10472_, _07613_, _09806_);
  or (_10473_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_10474_, _10473_, _10472_);
  and (_10475_, _10474_, _07643_);
  nand (_10477_, _07613_, _10026_);
  or (_10478_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_10479_, _10478_, _10477_);
  and (_10480_, _10479_, _07640_);
  or (_10481_, _10480_, _10475_);
  or (_10482_, _10481_, _10471_);
  nand (_10483_, _07613_, _10248_);
  or (_10484_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_10485_, _10484_, _10483_);
  and (_10486_, _10485_, _07650_);
  or (_10487_, _10486_, _07676_);
  or (_10488_, _10487_, _10482_);
  nand (_10490_, _07613_, _08685_);
  or (_10491_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_10493_, _10491_, _10490_);
  and (_10495_, _10493_, _07666_);
  nand (_10496_, _07613_, _08937_);
  or (_10497_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_10498_, _10497_, _10496_);
  and (_10500_, _10498_, _07643_);
  nand (_10501_, _07613_, _09150_);
  or (_10502_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_10504_, _10502_, _10501_);
  and (_10505_, _10504_, _07640_);
  or (_10506_, _10505_, _10500_);
  or (_10507_, _10506_, _10495_);
  nand (_10508_, _07613_, _09354_);
  or (_10509_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_10511_, _10509_, _10508_);
  and (_10512_, _10511_, _07650_);
  or (_10513_, _10512_, _07626_);
  or (_10514_, _10513_, _10507_);
  and (_10515_, _10514_, _10488_);
  and (_10516_, _10515_, _07705_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _10516_, _10467_);
  and (_10517_, _07758_, word_in[2]);
  nand (_10518_, _07613_, _09604_);
  or (_10519_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_10520_, _10519_, _10518_);
  and (_10521_, _10520_, _07666_);
  nand (_10522_, _07613_, _10038_);
  or (_10523_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_10524_, _10523_, _10522_);
  and (_10525_, _10524_, _07640_);
  nand (_10526_, _07613_, _09820_);
  or (_10527_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_10528_, _10527_, _10526_);
  and (_10530_, _10528_, _07643_);
  or (_10531_, _10530_, _10525_);
  or (_10532_, _10531_, _10521_);
  nand (_10533_, _07613_, _10260_);
  or (_10534_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_10535_, _10534_, _10533_);
  and (_10536_, _10535_, _07650_);
  or (_10537_, _10536_, _07676_);
  or (_10538_, _10537_, _10532_);
  nand (_10539_, _07613_, _08700_);
  or (_10541_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_10542_, _10541_, _10539_);
  and (_10543_, _10542_, _07666_);
  nand (_10544_, _07613_, _08949_);
  or (_10545_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_10546_, _10545_, _10544_);
  and (_10547_, _10546_, _07643_);
  nand (_10548_, _07613_, _09161_);
  or (_10549_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_10550_, _10549_, _10548_);
  and (_10551_, _10550_, _07640_);
  or (_10552_, _10551_, _10547_);
  or (_10553_, _10552_, _10543_);
  nand (_10554_, _07613_, _09366_);
  or (_10556_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_10558_, _10556_, _10554_);
  and (_10559_, _10558_, _07650_);
  or (_10560_, _10559_, _07626_);
  or (_10561_, _10560_, _10553_);
  and (_10562_, _10561_, _10538_);
  and (_10563_, _10562_, _07705_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _10563_, _10517_);
  and (_10564_, _07758_, word_in[3]);
  nand (_10565_, _07613_, _09617_);
  or (_10566_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_10567_, _10566_, _10565_);
  and (_10568_, _10567_, _07666_);
  nand (_10569_, _07613_, _10050_);
  or (_10571_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_10572_, _10571_, _10569_);
  and (_10573_, _10572_, _07640_);
  nand (_10574_, _07613_, _09832_);
  or (_10576_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_10577_, _10576_, _10574_);
  and (_10578_, _10577_, _07643_);
  or (_10579_, _10578_, _10573_);
  or (_10580_, _10579_, _10568_);
  nand (_10581_, _07613_, _10272_);
  or (_10582_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_10584_, _10582_, _10581_);
  and (_10585_, _10584_, _07650_);
  or (_10586_, _10585_, _07676_);
  or (_10587_, _10586_, _10580_);
  nand (_10588_, _07613_, _08714_);
  or (_10589_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_10590_, _10589_, _10588_);
  and (_10591_, _10590_, _07666_);
  nand (_10592_, _07613_, _08960_);
  or (_10593_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_10594_, _10593_, _10592_);
  and (_10595_, _10594_, _07643_);
  nand (_10596_, _07613_, _09175_);
  or (_10597_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_10598_, _10597_, _10596_);
  and (_10599_, _10598_, _07640_);
  or (_10600_, _10599_, _10595_);
  or (_10601_, _10600_, _10591_);
  nand (_10602_, _07613_, _09378_);
  or (_10603_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_10604_, _10603_, _10602_);
  and (_10605_, _10604_, _07650_);
  or (_10606_, _10605_, _07626_);
  or (_10607_, _10606_, _10601_);
  and (_10608_, _10607_, _10587_);
  and (_10609_, _10608_, _07705_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _10609_, _10564_);
  and (_10611_, _07758_, word_in[4]);
  nand (_10612_, _07613_, _09628_);
  or (_10613_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_10614_, _10613_, _10612_);
  and (_10615_, _10614_, _07666_);
  nand (_10616_, _07613_, _09845_);
  or (_10617_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_10618_, _10617_, _10616_);
  and (_10619_, _10618_, _07643_);
  nand (_10620_, _07613_, _10071_);
  or (_10621_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_10622_, _10621_, _10620_);
  and (_10623_, _10622_, _07640_);
  or (_10624_, _10623_, _10619_);
  or (_10625_, _10624_, _10615_);
  nand (_10626_, _07613_, _10286_);
  or (_10627_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_10628_, _10627_, _10626_);
  and (_10629_, _10628_, _07650_);
  or (_10630_, _10629_, _07676_);
  or (_10631_, _10630_, _10625_);
  nand (_10632_, _07613_, _08726_);
  or (_10633_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_10634_, _10633_, _10632_);
  and (_10635_, _10634_, _07666_);
  nand (_10636_, _07613_, _08972_);
  or (_10637_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_10638_, _10637_, _10636_);
  and (_10639_, _10638_, _07643_);
  nand (_10641_, _07613_, _09186_);
  or (_10642_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_10643_, _10642_, _10641_);
  and (_10644_, _10643_, _07640_);
  or (_10645_, _10644_, _10639_);
  or (_10646_, _10645_, _10635_);
  nand (_10648_, _07613_, _09390_);
  or (_10649_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_10650_, _10649_, _10648_);
  and (_10651_, _10650_, _07650_);
  or (_10652_, _10651_, _07626_);
  or (_10653_, _10652_, _10646_);
  and (_10654_, _10653_, _10631_);
  and (_10655_, _10654_, _07705_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _10655_, _10611_);
  and (_10657_, _07758_, word_in[5]);
  nand (_10658_, _07613_, _09858_);
  or (_10659_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_10660_, _10659_, _10658_);
  and (_10661_, _10660_, _07643_);
  nand (_10662_, _07613_, _10084_);
  or (_10663_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_10664_, _10663_, _10662_);
  and (_10665_, _10664_, _07640_);
  nand (_10666_, _07613_, _09640_);
  or (_10667_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_10668_, _10667_, _10666_);
  and (_10669_, _10668_, _07666_);
  or (_10670_, _10669_, _10665_);
  or (_10671_, _10670_, _10661_);
  nand (_10672_, _07613_, _10298_);
  or (_10673_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_10674_, _10673_, _10672_);
  and (_10675_, _10674_, _07650_);
  or (_10676_, _10675_, _07676_);
  or (_10677_, _10676_, _10671_);
  nand (_10678_, _07613_, _08984_);
  or (_10679_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_10680_, _10679_, _10678_);
  and (_10681_, _10680_, _07643_);
  nand (_10682_, _07613_, _08739_);
  or (_10683_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_10684_, _10683_, _10682_);
  and (_10685_, _10684_, _07666_);
  nand (_10686_, _07613_, _09198_);
  or (_10687_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_10688_, _10687_, _10686_);
  and (_10689_, _10688_, _07640_);
  or (_10690_, _10689_, _10685_);
  or (_10691_, _10690_, _10681_);
  nand (_10692_, _07613_, _09402_);
  or (_10693_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_10694_, _10693_, _10692_);
  and (_10695_, _10694_, _07650_);
  or (_10696_, _10695_, _07626_);
  or (_10697_, _10696_, _10691_);
  and (_10699_, _10697_, _10677_);
  and (_10700_, _10699_, _07705_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _10700_, _10657_);
  and (_10701_, _07758_, word_in[6]);
  nand (_10702_, _07613_, _09872_);
  or (_10703_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_10704_, _10703_, _10702_);
  and (_10705_, _10704_, _07643_);
  nand (_10706_, _07613_, _10096_);
  or (_10707_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_10708_, _10707_, _10706_);
  and (_10709_, _10708_, _07640_);
  nand (_10710_, _07613_, _09652_);
  or (_10711_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_10712_, _10711_, _10710_);
  and (_10713_, _10712_, _07666_);
  or (_10714_, _10713_, _10709_);
  or (_10716_, _10714_, _10705_);
  nand (_10717_, _07613_, _10309_);
  or (_10719_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_10720_, _10719_, _10717_);
  and (_10721_, _10720_, _07650_);
  or (_10722_, _10721_, _07676_);
  or (_10723_, _10722_, _10716_);
  nand (_10724_, _07613_, _08998_);
  or (_10725_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_10726_, _10725_, _10724_);
  and (_10727_, _10726_, _07643_);
  nand (_10728_, _07613_, _08752_);
  or (_10729_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_10730_, _10729_, _10728_);
  and (_10731_, _10730_, _07666_);
  nand (_10732_, _07613_, _09211_);
  or (_10733_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_10734_, _10733_, _10732_);
  and (_10735_, _10734_, _07640_);
  or (_10736_, _10735_, _10731_);
  or (_10737_, _10736_, _10727_);
  nand (_10738_, _07613_, _09413_);
  or (_10739_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_10740_, _10739_, _10738_);
  and (_10741_, _10740_, _07650_);
  or (_10743_, _10741_, _07626_);
  or (_10744_, _10743_, _10737_);
  and (_10745_, _10744_, _10723_);
  and (_10746_, _10745_, _07705_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _10746_, _10701_);
  and (_10748_, _07819_, word_in[8]);
  nand (_10749_, _07613_, _08790_);
  or (_10751_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_10752_, _10751_, _10749_);
  and (_10753_, _10752_, _07821_);
  nand (_10754_, _07613_, _08535_);
  or (_10755_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_10756_, _10755_, _10754_);
  and (_10757_, _10756_, _07820_);
  or (_10758_, _10757_, _10753_);
  and (_10759_, _10758_, _07781_);
  nand (_10760_, _07613_, _09680_);
  or (_10761_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_10762_, _10761_, _10760_);
  and (_10763_, _10762_, _07821_);
  nand (_10764_, _07613_, _09468_);
  or (_10765_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_10766_, _10765_, _10764_);
  and (_10767_, _10766_, _07820_);
  or (_10768_, _10767_, _10763_);
  and (_10769_, _10768_, _07783_);
  nand (_10770_, _07613_, _09236_);
  or (_10771_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_10772_, _10771_, _10770_);
  and (_10773_, _10772_, _07821_);
  nand (_10774_, _07613_, _09025_);
  or (_10775_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_10776_, _10775_, _10774_);
  and (_10777_, _10776_, _07820_);
  or (_10778_, _10777_, _10773_);
  and (_10779_, _10778_, _07807_);
  nand (_10780_, _07613_, _10131_);
  or (_10781_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_10782_, _10781_, _10780_);
  and (_10783_, _10782_, _07821_);
  nand (_10784_, _07613_, _09908_);
  or (_10785_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_10786_, _10785_, _10784_);
  and (_10787_, _10786_, _07820_);
  or (_10788_, _10787_, _10783_);
  and (_10789_, _10788_, _07811_);
  or (_10790_, _10789_, _10779_);
  or (_10791_, _10790_, _10769_);
  nor (_10793_, _10791_, _10759_);
  nor (_10794_, _10793_, _07819_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _10794_, _10748_);
  and (_10795_, _07819_, word_in[9]);
  nand (_10796_, _07613_, _08810_);
  or (_10797_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_10798_, _10797_, _10796_);
  and (_10799_, _10798_, _07821_);
  nand (_10801_, _07613_, _08554_);
  or (_10802_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_10803_, _10802_, _10801_);
  and (_10804_, _10803_, _07820_);
  or (_10805_, _10804_, _10799_);
  and (_10806_, _10805_, _07781_);
  nand (_10807_, _07613_, _09695_);
  or (_10808_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_10809_, _10808_, _10807_);
  and (_10810_, _10809_, _07821_);
  nand (_10811_, _07613_, _09483_);
  or (_10812_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_10813_, _10812_, _10811_);
  and (_10814_, _10813_, _07820_);
  or (_10815_, _10814_, _10810_);
  and (_10816_, _10815_, _07783_);
  nand (_10817_, _07613_, _09253_);
  or (_10818_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_10819_, _10818_, _10817_);
  and (_10820_, _10819_, _07821_);
  nand (_10821_, _07613_, _09043_);
  or (_10822_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_10823_, _10822_, _10821_);
  and (_10824_, _10823_, _07820_);
  or (_10825_, _10824_, _10820_);
  and (_10826_, _10825_, _07807_);
  nand (_10827_, _07613_, _10146_);
  or (_10828_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_10829_, _10828_, _10827_);
  and (_10830_, _10829_, _07821_);
  nand (_10831_, _07613_, _09924_);
  or (_10832_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_10833_, _10832_, _10831_);
  and (_10834_, _10833_, _07820_);
  or (_10835_, _10834_, _10830_);
  and (_10836_, _10835_, _07811_);
  or (_10837_, _10836_, _10826_);
  or (_10838_, _10837_, _10816_);
  nor (_10839_, _10838_, _10806_);
  nor (_10840_, _10839_, _07819_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _10840_, _10795_);
  and (_10841_, _07819_, word_in[10]);
  nand (_10842_, _07613_, _08823_);
  or (_10843_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_10844_, _10843_, _10842_);
  and (_10845_, _10844_, _07821_);
  nand (_10846_, _07613_, _08570_);
  or (_10847_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_10848_, _10847_, _10846_);
  and (_10849_, _10848_, _07820_);
  or (_10850_, _10849_, _10845_);
  and (_10851_, _10850_, _07781_);
  nand (_10852_, _07613_, _09708_);
  or (_10853_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_10854_, _10853_, _10852_);
  and (_10855_, _10854_, _07821_);
  nand (_10856_, _07613_, _09495_);
  or (_10857_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_10858_, _10857_, _10856_);
  and (_10859_, _10858_, _07820_);
  or (_10860_, _10859_, _10855_);
  and (_10861_, _10860_, _07783_);
  nand (_10862_, _07613_, _09264_);
  or (_10863_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_10864_, _10863_, _10862_);
  and (_10865_, _10864_, _07821_);
  nand (_10866_, _07613_, _09055_);
  or (_10867_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_10868_, _10867_, _10866_);
  and (_10869_, _10868_, _07820_);
  or (_10870_, _10869_, _10865_);
  and (_10872_, _10870_, _07807_);
  nand (_10873_, _07613_, _10159_);
  or (_10874_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_10875_, _10874_, _10873_);
  and (_10876_, _10875_, _07821_);
  nand (_10877_, _07613_, _09936_);
  or (_10878_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_10879_, _10878_, _10877_);
  and (_10880_, _10879_, _07820_);
  or (_10881_, _10880_, _10876_);
  and (_10882_, _10881_, _07811_);
  or (_10883_, _10882_, _10872_);
  or (_10884_, _10883_, _10861_);
  nor (_10885_, _10884_, _10851_);
  nor (_10886_, _10885_, _07819_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _10886_, _10841_);
  and (_10888_, _07819_, word_in[11]);
  nand (_10889_, _07613_, _08836_);
  or (_10891_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_10892_, _10891_, _10889_);
  and (_10893_, _10892_, _07821_);
  nand (_10894_, _07613_, _08584_);
  or (_10895_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_10896_, _10895_, _10894_);
  and (_10897_, _10896_, _07820_);
  or (_10898_, _10897_, _10893_);
  and (_10899_, _10898_, _07781_);
  nand (_10900_, _07613_, _09720_);
  or (_10901_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_10902_, _10901_, _10900_);
  and (_10903_, _10902_, _07821_);
  nand (_10904_, _07613_, _09507_);
  or (_10905_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_10906_, _10905_, _10904_);
  and (_10907_, _10906_, _07820_);
  or (_10908_, _10907_, _10903_);
  and (_10909_, _10908_, _07783_);
  nand (_10910_, _07613_, _09276_);
  or (_10911_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_10912_, _10911_, _10910_);
  and (_10913_, _10912_, _07821_);
  nand (_10914_, _07613_, _09067_);
  or (_10915_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_10916_, _10915_, _10914_);
  and (_10917_, _10916_, _07820_);
  or (_10918_, _10917_, _10913_);
  and (_10919_, _10918_, _07807_);
  nand (_10920_, _07613_, _10172_);
  or (_10921_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_10922_, _10921_, _10920_);
  and (_10923_, _10922_, _07821_);
  nand (_10924_, _07613_, _09948_);
  or (_10925_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_10926_, _10925_, _10924_);
  and (_10927_, _10926_, _07820_);
  or (_10928_, _10927_, _10923_);
  and (_10929_, _10928_, _07811_);
  or (_10930_, _10929_, _10919_);
  or (_10931_, _10930_, _10909_);
  nor (_10932_, _10931_, _10899_);
  nor (_10933_, _10932_, _07819_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _10933_, _10888_);
  and (_10934_, _07819_, word_in[12]);
  nand (_10935_, _07613_, _08850_);
  or (_10937_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_10938_, _10937_, _10935_);
  and (_10939_, _10938_, _07821_);
  nand (_10941_, _07613_, _08596_);
  or (_10942_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_10944_, _10942_, _10941_);
  and (_10945_, _10944_, _07820_);
  or (_10946_, _10945_, _10939_);
  and (_10947_, _10946_, _07781_);
  nand (_10948_, _07613_, _09731_);
  or (_10949_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_10950_, _10949_, _10948_);
  and (_10951_, _10950_, _07821_);
  nand (_10952_, _07613_, _09519_);
  or (_10953_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_10954_, _10953_, _10952_);
  and (_10955_, _10954_, _07820_);
  or (_10956_, _10955_, _10951_);
  and (_10957_, _10956_, _07783_);
  nand (_10958_, _07613_, _09289_);
  or (_10959_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_10960_, _10959_, _10958_);
  and (_10961_, _10960_, _07821_);
  nand (_10962_, _07613_, _09079_);
  or (_10963_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_10964_, _10963_, _10962_);
  and (_10965_, _10964_, _07820_);
  or (_10966_, _10965_, _10961_);
  and (_10967_, _10966_, _07807_);
  nand (_10968_, _07613_, _10184_);
  or (_10969_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_10970_, _10969_, _10968_);
  and (_10971_, _10970_, _07821_);
  nand (_10972_, _07613_, _09960_);
  or (_10973_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_10974_, _10973_, _10972_);
  and (_10975_, _10974_, _07820_);
  or (_10976_, _10975_, _10971_);
  and (_10977_, _10976_, _07811_);
  or (_10978_, _10977_, _10967_);
  or (_10979_, _10978_, _10957_);
  nor (_10980_, _10979_, _10947_);
  nor (_10981_, _10980_, _07819_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _10981_, _10934_);
  and (_10982_, _07819_, word_in[13]);
  nand (_10983_, _07613_, _08862_);
  or (_10984_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_10985_, _10984_, _10983_);
  and (_10987_, _10985_, _07821_);
  nand (_10988_, _07613_, _08610_);
  or (_10989_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_10990_, _10989_, _10988_);
  and (_10991_, _10990_, _07820_);
  or (_10992_, _10991_, _10987_);
  and (_10993_, _10992_, _07781_);
  nand (_10994_, _07613_, _09744_);
  or (_10995_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_10996_, _10995_, _10994_);
  and (_10997_, _10996_, _07821_);
  nand (_10998_, _07613_, _09531_);
  or (_10999_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_11000_, _10999_, _10998_);
  and (_11001_, _11000_, _07820_);
  or (_11002_, _11001_, _10997_);
  and (_11003_, _11002_, _07783_);
  nand (_11004_, _07613_, _09301_);
  or (_11005_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_11006_, _11005_, _11004_);
  and (_11007_, _11006_, _07821_);
  nand (_11008_, _07613_, _09091_);
  or (_11009_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_11010_, _11009_, _11008_);
  and (_11011_, _11010_, _07820_);
  or (_11012_, _11011_, _11007_);
  and (_11013_, _11012_, _07807_);
  nand (_11014_, _07613_, _10197_);
  or (_11015_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_11016_, _11015_, _11014_);
  and (_11017_, _11016_, _07821_);
  nand (_11018_, _07613_, _09972_);
  or (_11019_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_11020_, _11019_, _11018_);
  and (_11021_, _11020_, _07820_);
  or (_11022_, _11021_, _11017_);
  and (_11023_, _11022_, _07811_);
  or (_11024_, _11023_, _11013_);
  or (_11025_, _11024_, _11003_);
  nor (_11026_, _11025_, _10993_);
  nor (_11027_, _11026_, _07819_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _11027_, _10982_);
  and (_11028_, _07819_, word_in[14]);
  nand (_11029_, _07613_, _08890_);
  or (_11031_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_11032_, _11031_, _11029_);
  and (_11033_, _11032_, _07821_);
  nand (_11035_, _07613_, _08626_);
  or (_11036_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_11037_, _11036_, _11035_);
  and (_11038_, _11037_, _07820_);
  or (_11039_, _11038_, _11033_);
  and (_11040_, _11039_, _07781_);
  nand (_11041_, _07613_, _09756_);
  or (_11042_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_11043_, _11042_, _11041_);
  and (_11044_, _11043_, _07821_);
  nand (_11045_, _07613_, _09543_);
  or (_11046_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_11047_, _11046_, _11045_);
  and (_11048_, _11047_, _07820_);
  or (_11049_, _11048_, _11044_);
  and (_11050_, _11049_, _07783_);
  nand (_11051_, _07613_, _09313_);
  or (_11052_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_11053_, _11052_, _11051_);
  and (_11054_, _11053_, _07821_);
  nand (_11055_, _07613_, _09103_);
  or (_11056_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_11057_, _11056_, _11055_);
  and (_11058_, _11057_, _07820_);
  or (_11059_, _11058_, _11054_);
  and (_11060_, _11059_, _07807_);
  nand (_11061_, _07613_, _10209_);
  or (_11062_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_11064_, _11062_, _11061_);
  and (_11065_, _11064_, _07821_);
  nand (_11066_, _07613_, _09984_);
  or (_11067_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_11069_, _11067_, _11066_);
  and (_11070_, _11069_, _07820_);
  or (_11071_, _11070_, _11065_);
  and (_11072_, _11071_, _07811_);
  or (_11073_, _11072_, _11060_);
  or (_11074_, _11073_, _11050_);
  nor (_11075_, _11074_, _11040_);
  nor (_11076_, _11075_, _07819_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _11076_, _11028_);
  and (_11078_, _07917_, word_in[16]);
  and (_11079_, _10453_, _07643_);
  and (_11080_, _10445_, _07650_);
  or (_11081_, _11080_, _11079_);
  and (_11082_, _10460_, _07640_);
  and (_11083_, _10449_, _07666_);
  or (_11084_, _11083_, _11082_);
  or (_11085_, _11084_, _11081_);
  or (_11086_, _11085_, _07888_);
  and (_11087_, _10424_, _07650_);
  and (_11088_, _10439_, _07640_);
  or (_11089_, _11088_, _11087_);
  and (_11090_, _10432_, _07643_);
  and (_11091_, _10428_, _07666_);
  or (_11092_, _11091_, _11090_);
  or (_11093_, _11092_, _11089_);
  or (_11095_, _11093_, _07927_);
  nand (_11096_, _11095_, _11086_);
  nor (_11097_, _11096_, _07917_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _11097_, _11078_);
  and (_11099_, _07917_, word_in[17]);
  and (_11101_, _10504_, _07643_);
  and (_11102_, _10493_, _07650_);
  or (_11103_, _11102_, _11101_);
  and (_11105_, _10511_, _07640_);
  and (_11106_, _10498_, _07666_);
  or (_11108_, _11106_, _11105_);
  or (_11109_, _11108_, _11103_);
  or (_11110_, _11109_, _07888_);
  and (_11111_, _10470_, _07650_);
  and (_11112_, _10485_, _07640_);
  or (_11113_, _11112_, _11111_);
  and (_11114_, _10479_, _07643_);
  and (_11115_, _10474_, _07666_);
  or (_11116_, _11115_, _11114_);
  or (_11117_, _11116_, _11113_);
  or (_11118_, _11117_, _07927_);
  nand (_11119_, _11118_, _11110_);
  nor (_11120_, _11119_, _07917_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _11120_, _11099_);
  and (_11121_, _07917_, word_in[18]);
  and (_11122_, _10542_, _07650_);
  and (_11123_, _10558_, _07640_);
  or (_11124_, _11123_, _11122_);
  and (_11125_, _10550_, _07643_);
  and (_11126_, _10546_, _07666_);
  or (_11127_, _11126_, _11125_);
  or (_11128_, _11127_, _11124_);
  or (_11129_, _11128_, _07888_);
  and (_11130_, _10524_, _07643_);
  and (_11131_, _10520_, _07650_);
  or (_11132_, _11131_, _11130_);
  and (_11133_, _10535_, _07640_);
  and (_11134_, _10528_, _07666_);
  or (_11135_, _11134_, _11133_);
  or (_11136_, _11135_, _11132_);
  or (_11137_, _11136_, _07927_);
  nand (_11138_, _11137_, _11129_);
  nor (_11139_, _11138_, _07917_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _11139_, _11121_);
  and (_11140_, _07917_, word_in[19]);
  and (_11141_, _10590_, _07650_);
  and (_11142_, _10604_, _07640_);
  or (_11143_, _11142_, _11141_);
  and (_11144_, _10598_, _07643_);
  and (_11145_, _10594_, _07666_);
  or (_11146_, _11145_, _11144_);
  or (_11147_, _11146_, _11143_);
  or (_11148_, _11147_, _07888_);
  and (_11149_, _10567_, _07650_);
  and (_11150_, _10584_, _07640_);
  or (_11151_, _11150_, _11149_);
  and (_11152_, _10572_, _07643_);
  and (_11153_, _10577_, _07666_);
  or (_11154_, _11153_, _11152_);
  or (_11155_, _11154_, _11151_);
  or (_11156_, _11155_, _07927_);
  nand (_11157_, _11156_, _11148_);
  nor (_11158_, _11157_, _07917_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _11158_, _11140_);
  and (_11159_, _07917_, word_in[20]);
  and (_11160_, _10643_, _07643_);
  and (_11162_, _10634_, _07650_);
  or (_11164_, _11162_, _11160_);
  and (_11165_, _10650_, _07640_);
  and (_11167_, _10638_, _07666_);
  or (_11168_, _11167_, _11165_);
  or (_11169_, _11168_, _11164_);
  or (_11170_, _11169_, _07888_);
  and (_11171_, _10614_, _07650_);
  and (_11172_, _10628_, _07640_);
  or (_11173_, _11172_, _11171_);
  and (_11174_, _10622_, _07643_);
  and (_11175_, _10618_, _07666_);
  or (_11176_, _11175_, _11174_);
  or (_11177_, _11176_, _11173_);
  or (_11178_, _11177_, _07927_);
  nand (_11179_, _11178_, _11170_);
  nor (_11181_, _11179_, _07917_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _11181_, _11159_);
  and (_11182_, _07917_, word_in[21]);
  and (_11183_, _10688_, _07643_);
  and (_11184_, _10684_, _07650_);
  or (_11185_, _11184_, _11183_);
  and (_11186_, _10694_, _07640_);
  and (_11187_, _10680_, _07666_);
  or (_11188_, _11187_, _11186_);
  or (_11189_, _11188_, _11185_);
  or (_11190_, _11189_, _07888_);
  and (_11191_, _10664_, _07643_);
  and (_11192_, _10668_, _07650_);
  or (_11193_, _11192_, _11191_);
  and (_11194_, _10674_, _07640_);
  and (_11195_, _10660_, _07666_);
  or (_11196_, _11195_, _11194_);
  or (_11197_, _11196_, _11193_);
  or (_11198_, _11197_, _07927_);
  nand (_11199_, _11198_, _11190_);
  nor (_11200_, _11199_, _07917_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _11200_, _11182_);
  and (_11201_, _07917_, word_in[22]);
  and (_11202_, _10734_, _07643_);
  and (_11203_, _10730_, _07650_);
  or (_11204_, _11203_, _11202_);
  and (_11205_, _10740_, _07640_);
  and (_11206_, _10726_, _07666_);
  or (_11207_, _11206_, _11205_);
  or (_11208_, _11207_, _11204_);
  or (_11209_, _11208_, _07888_);
  and (_11210_, _10712_, _07650_);
  and (_11211_, _10720_, _07640_);
  or (_11212_, _11211_, _11210_);
  and (_11213_, _10708_, _07643_);
  and (_11215_, _10704_, _07666_);
  or (_11216_, _11215_, _11213_);
  or (_11218_, _11216_, _11212_);
  or (_11219_, _11218_, _07927_);
  nand (_11220_, _11219_, _11209_);
  nor (_11222_, _11220_, _07917_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _11222_, _11201_);
  and (_11223_, _07984_, word_in[24]);
  and (_11224_, _10766_, _07821_);
  and (_11225_, _10762_, _07820_);
  or (_11226_, _11225_, _11224_);
  and (_11227_, _11226_, _07949_);
  and (_11228_, _10756_, _07821_);
  and (_11230_, _10752_, _07820_);
  or (_11231_, _11230_, _11228_);
  and (_11232_, _11231_, _07947_);
  and (_11233_, _10776_, _07821_);
  and (_11234_, _10772_, _07820_);
  or (_11235_, _11234_, _11233_);
  and (_11237_, _11235_, _07993_);
  and (_11238_, _10786_, _07821_);
  and (_11240_, _10782_, _07820_);
  or (_11241_, _11240_, _11238_);
  and (_11242_, _11241_, _08001_);
  or (_11243_, _11242_, _11237_);
  or (_11244_, _11243_, _11232_);
  nor (_11245_, _11244_, _11227_);
  nor (_11246_, _11245_, _07984_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _11246_, _11223_);
  and (_11247_, _07984_, word_in[25]);
  and (_11248_, _10813_, _07821_);
  and (_11249_, _10809_, _07820_);
  or (_11250_, _11249_, _11248_);
  and (_11251_, _11250_, _07949_);
  and (_11252_, _10803_, _07821_);
  and (_11253_, _10798_, _07820_);
  or (_11255_, _11253_, _11252_);
  and (_11256_, _11255_, _07947_);
  and (_11257_, _10823_, _07821_);
  and (_11258_, _10819_, _07820_);
  or (_11260_, _11258_, _11257_);
  and (_11261_, _11260_, _07993_);
  and (_11262_, _10833_, _07821_);
  and (_11264_, _10829_, _07820_);
  or (_11265_, _11264_, _11262_);
  and (_11266_, _11265_, _08001_);
  or (_11267_, _11266_, _11261_);
  or (_11268_, _11267_, _11256_);
  nor (_11269_, _11268_, _11251_);
  nor (_11270_, _11269_, _07984_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _11270_, _11247_);
  and (_11271_, _07984_, word_in[26]);
  and (_11272_, _10848_, _07821_);
  and (_11273_, _10844_, _07820_);
  or (_11274_, _11273_, _11272_);
  and (_11275_, _11274_, _07947_);
  and (_11276_, _10858_, _07821_);
  and (_11277_, _10854_, _07820_);
  or (_11278_, _11277_, _11276_);
  and (_11279_, _11278_, _07949_);
  and (_11280_, _10868_, _07821_);
  and (_11282_, _10864_, _07820_);
  or (_11283_, _11282_, _11280_);
  and (_11284_, _11283_, _07993_);
  and (_11285_, _10879_, _07821_);
  and (_11286_, _10875_, _07820_);
  or (_11287_, _11286_, _11285_);
  and (_11288_, _11287_, _08001_);
  or (_11289_, _11288_, _11284_);
  or (_11290_, _11289_, _11279_);
  nor (_11291_, _11290_, _11275_);
  nor (_11292_, _11291_, _07984_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _11292_, _11271_);
  and (_11293_, _07984_, word_in[27]);
  and (_11294_, _10906_, _07821_);
  and (_11295_, _10902_, _07820_);
  or (_11296_, _11295_, _11294_);
  and (_11297_, _11296_, _07949_);
  and (_11298_, _10896_, _07821_);
  and (_11299_, _10892_, _07820_);
  or (_11301_, _11299_, _11298_);
  and (_11302_, _11301_, _07947_);
  and (_11303_, _10916_, _07821_);
  and (_11304_, _10912_, _07820_);
  or (_11305_, _11304_, _11303_);
  and (_11306_, _11305_, _07993_);
  and (_11307_, _10926_, _07821_);
  and (_11308_, _10922_, _07820_);
  or (_11309_, _11308_, _11307_);
  and (_11311_, _11309_, _08001_);
  or (_11312_, _11311_, _11306_);
  or (_11313_, _11312_, _11302_);
  nor (_11314_, _11313_, _11297_);
  nor (_11315_, _11314_, _07984_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _11315_, _11293_);
  and (_11316_, _07984_, word_in[28]);
  and (_11317_, _10954_, _07821_);
  and (_11318_, _10950_, _07820_);
  or (_11320_, _11318_, _11317_);
  and (_11321_, _11320_, _07949_);
  and (_11322_, _10944_, _07821_);
  and (_11324_, _10938_, _07820_);
  or (_11325_, _11324_, _11322_);
  and (_11326_, _11325_, _07947_);
  and (_11327_, _10964_, _07821_);
  and (_11328_, _10960_, _07820_);
  or (_11329_, _11328_, _11327_);
  and (_11330_, _11329_, _07993_);
  and (_11331_, _10974_, _07821_);
  and (_11332_, _10970_, _07820_);
  or (_11333_, _11332_, _11331_);
  and (_11334_, _11333_, _08001_);
  or (_11336_, _11334_, _11330_);
  or (_11337_, _11336_, _11326_);
  nor (_11338_, _11337_, _11321_);
  nor (_11339_, _11338_, _07984_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _11339_, _11316_);
  and (_11340_, _07984_, word_in[29]);
  and (_11341_, _11000_, _07821_);
  and (_11342_, _10996_, _07820_);
  or (_11343_, _11342_, _11341_);
  and (_11344_, _11343_, _07949_);
  and (_11345_, _10990_, _07821_);
  and (_11347_, _10985_, _07820_);
  or (_11348_, _11347_, _11345_);
  and (_11349_, _11348_, _07947_);
  and (_11350_, _11010_, _07821_);
  and (_11351_, _11006_, _07820_);
  or (_11352_, _11351_, _11350_);
  and (_11353_, _11352_, _07993_);
  and (_11354_, _11020_, _07821_);
  and (_11355_, _11016_, _07820_);
  or (_11357_, _11355_, _11354_);
  and (_11358_, _11357_, _08001_);
  or (_11359_, _11358_, _11353_);
  or (_11361_, _11359_, _11349_);
  nor (_11362_, _11361_, _11344_);
  nor (_11364_, _11362_, _07984_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _11364_, _11340_);
  and (_11365_, _07984_, word_in[30]);
  and (_11366_, _11037_, _07821_);
  and (_11367_, _11032_, _07820_);
  or (_11368_, _11367_, _11366_);
  and (_11369_, _11368_, _07947_);
  and (_11370_, _11047_, _07821_);
  and (_11371_, _11043_, _07820_);
  or (_11372_, _11371_, _11370_);
  and (_11373_, _11372_, _07949_);
  and (_11374_, _11057_, _07821_);
  and (_11375_, _11053_, _07820_);
  or (_11377_, _11375_, _11374_);
  and (_11378_, _11377_, _07993_);
  and (_11379_, _11069_, _07821_);
  and (_11380_, _11064_, _07820_);
  or (_11381_, _11380_, _11379_);
  and (_11382_, _11381_, _08001_);
  or (_11383_, _11382_, _11378_);
  or (_11384_, _11383_, _11373_);
  nor (_11385_, _11384_, _11369_);
  nor (_11386_, _11385_, _07984_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _11386_, _11365_);
  nand (_11387_, _06415_, _06270_);
  or (_11388_, _06270_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_11390_, _11388_, _05141_);
  and (_09833_, _11390_, _11387_);
  or (_11391_, _06497_, _07117_);
  or (_11392_, _06270_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_11393_, _11392_, _05141_);
  and (_09855_, _11393_, _11391_);
  or (_11394_, _06447_, _07117_);
  or (_11395_, _06270_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_11396_, _11395_, _05141_);
  and (_09859_, _11396_, _11394_);
  or (_11397_, _06524_, _07117_);
  or (_11398_, _06270_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_11399_, _11398_, _05141_);
  and (_09862_, _11399_, _11397_);
  and (_11400_, _08382_, _06004_);
  and (_11401_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_11402_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_11403_, _11402_, _11401_);
  nor (_11404_, _11403_, _08243_);
  and (_11405_, _08396_, _05522_);
  or (_11406_, _11405_, _11404_);
  or (_11407_, _11406_, _11400_);
  and (_10068_, _11407_, _05141_);
  nor (_11408_, _08656_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_11410_, _11408_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_11411_, _11408_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_11412_, _11411_, _05141_);
  and (_10072_, _11412_, _11410_);
  nand (_11413_, _07350_, _06624_);
  or (_11414_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_11415_, _11414_, _05141_);
  and (_10236_, _11415_, _11413_);
  nor (_11417_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_11418_, _11417_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_03037_, _11418_, _05141_);
  and (_10494_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _05141_);
  and (_11419_, _10494_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_10245_, _11419_, _03037_);
  not (_11420_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_11421_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , _11420_);
  and (_10251_, _11421_, _05141_);
  and (_11422_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_11423_, _11422_);
  nand (_11424_, _08344_, _05143_);
  and (_11425_, _11424_, _11423_);
  and (_11426_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_11427_, _11426_);
  or (_11428_, _06564_, _06556_);
  and (_11429_, _11428_, _06771_);
  and (_11430_, _06771_, _06563_);
  and (_11431_, _11430_, _06450_);
  nor (_11432_, _11431_, _11429_);
  or (_11433_, _07053_, _06529_);
  nand (_11434_, _11433_, _06771_);
  nand (_11435_, _07044_, _06449_);
  and (_11436_, _11435_, _11434_);
  and (_11437_, _11436_, _11432_);
  nand (_11438_, _06556_, _06544_);
  not (_11439_, _11438_);
  nor (_11440_, _11439_, _07076_);
  and (_11441_, _07069_, _06766_);
  nor (_11442_, _11441_, _06772_);
  and (_11443_, _06771_, _06765_);
  nor (_11444_, _11443_, _06979_);
  and (_11445_, _11444_, _11442_);
  and (_11446_, _11445_, _11440_);
  and (_11447_, _11446_, _11437_);
  nand (_11448_, _11447_, _08337_);
  nand (_11449_, _11448_, _06821_);
  and (_11450_, _11439_, _07087_);
  and (_11451_, _11450_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_11452_, _07088_, _06575_);
  nor (_11453_, _11452_, _11451_);
  nand (_11454_, _11453_, _11449_);
  nand (_11455_, _11454_, _05143_);
  nand (_11456_, _11455_, _11427_);
  and (_11457_, _11456_, _11425_);
  and (_10319_, _11457_, _05141_);
  and (_10340_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _05141_);
  and (_11458_, _10343_, _06204_);
  and (_11459_, _11458_, _05288_);
  nand (_11460_, _11459_, _05963_);
  or (_11461_, _11459_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_11462_, _06734_, _05926_);
  not (_11463_, _11462_);
  and (_11464_, _11463_, _11461_);
  and (_11465_, _11464_, _11460_);
  nor (_11466_, _11463_, _06178_);
  or (_11467_, _11466_, _11465_);
  and (_10344_, _11467_, _05141_);
  and (_11468_, _11458_, _05210_);
  and (_11469_, _11468_, _05963_);
  nor (_11470_, _11468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_11471_, _11470_, _11469_);
  nand (_11472_, _11471_, _11463_);
  nand (_11473_, _11462_, _05604_);
  and (_11474_, _11473_, _05141_);
  and (_10347_, _11474_, _11472_);
  nor (_11475_, _07619_, _07516_);
  nor (_11476_, _06363_, _06337_);
  and (_11477_, _11476_, _07010_);
  not (_11478_, _11477_);
  and (_11479_, _06497_, _07023_);
  and (_11480_, _11479_, _07007_);
  and (_11481_, _06524_, _07006_);
  and (_11482_, _11481_, _07014_);
  nor (_11483_, _11482_, _11480_);
  nor (_11484_, _11483_, _11478_);
  not (_11485_, _11484_);
  and (_11486_, _06497_, _06447_);
  nor (_11487_, _06497_, _06447_);
  nor (_11488_, _11487_, _11486_);
  and (_11489_, _11488_, _07007_);
  and (_11490_, _11489_, _07018_);
  not (_11491_, _07021_);
  and (_11492_, _06524_, _06472_);
  and (_11493_, _11492_, _11479_);
  and (_11494_, _07006_, _06447_);
  and (_11495_, _11494_, _07007_);
  nor (_11496_, _11495_, _11493_);
  nor (_11497_, _11496_, _11491_);
  nor (_11498_, _11497_, _11490_);
  and (_11499_, _11498_, _11485_);
  and (_11500_, _11494_, _11492_);
  and (_11501_, _11500_, _11477_);
  not (_11502_, _11501_);
  nor (_11503_, _07017_, _06337_);
  and (_11504_, _11503_, _07010_);
  and (_11505_, _07023_, _06415_);
  and (_11506_, _06389_, _06337_);
  and (_11507_, _11506_, _11505_);
  and (_11508_, _11507_, _07007_);
  nor (_11509_, _11508_, _11504_);
  and (_11510_, _11509_, _11502_);
  and (_11511_, _11492_, _11486_);
  and (_11512_, _11511_, _07022_);
  and (_11513_, _11493_, _07011_);
  nor (_11514_, _11513_, _11512_);
  and (_11516_, _11514_, _11510_);
  and (_11517_, _06524_, _07014_);
  and (_11518_, _11517_, _11479_);
  and (_11519_, _07021_, _06363_);
  and (_11520_, _11519_, _11518_);
  not (_11521_, _11519_);
  and (_11522_, _11517_, _11487_);
  nor (_11524_, _11522_, _07015_);
  nor (_11525_, _11524_, _11521_);
  nor (_11527_, _11525_, _11520_);
  and (_11528_, _11527_, _11516_);
  and (_11529_, _11528_, _11499_);
  nor (_11530_, _07021_, _07018_);
  and (_11531_, _11492_, _11487_);
  and (_11532_, _11517_, _11486_);
  and (_11533_, _11519_, _11532_);
  nor (_11534_, _11533_, _11531_);
  nor (_11535_, _11534_, _11530_);
  not (_11536_, _11535_);
  and (_11537_, _07015_, _07006_);
  and (_11538_, _11537_, _07018_);
  not (_11539_, _11538_);
  and (_11540_, _11477_, _07015_);
  nand (_11541_, _11540_, _11488_);
  not (_11542_, _11541_);
  and (_11543_, _11517_, _11494_);
  and (_11544_, _11543_, _11519_);
  nor (_11545_, _11544_, _11542_);
  and (_11546_, _11545_, _11539_);
  and (_11547_, _11486_, _07007_);
  and (_11548_, _11547_, _07022_);
  and (_11549_, _11487_, _07007_);
  nor (_11550_, _11511_, _11549_);
  nor (_11551_, _11550_, _11521_);
  nor (_11552_, _11551_, _11548_);
  and (_11553_, _11552_, _11546_);
  and (_11554_, _11553_, _11536_);
  and (_11555_, _11554_, _11529_);
  and (_11556_, _07007_, _06497_);
  not (_11557_, _11556_);
  nor (_11558_, _11543_, _11511_);
  and (_11559_, _11558_, _11557_);
  nor (_11560_, _11559_, _06415_);
  not (_11561_, _11500_);
  nor (_11562_, _11530_, _11561_);
  nor (_11563_, _11562_, _11560_);
  and (_11564_, _11547_, _11519_);
  and (_11565_, _11500_, _07012_);
  nor (_11566_, _11565_, _11564_);
  not (_11567_, _11566_);
  not (_11568_, _07018_);
  nor (_11569_, _11522_, _11547_);
  and (_11570_, _11569_, _11558_);
  nor (_11571_, _11570_, _11568_);
  nor (_11572_, _11571_, _11567_);
  and (_11573_, _11572_, _11563_);
  not (_11574_, _11549_);
  nor (_11575_, _11477_, _07009_);
  and (_11576_, _11575_, _11568_);
  or (_11577_, _11576_, _11574_);
  and (_11578_, _06447_, _06415_);
  and (_11579_, _11506_, _11578_);
  and (_11580_, _11492_, _06497_);
  or (_11581_, _11556_, _11580_);
  and (_11582_, _11581_, _11579_);
  not (_11583_, _11582_);
  nand (_11584_, _11580_, _11477_);
  not (_11585_, _11584_);
  and (_11586_, _07022_, _07016_);
  nor (_11587_, _11586_, _11585_);
  and (_11588_, _11587_, _11583_);
  and (_11589_, _11588_, _11577_);
  and (_11590_, _11531_, _07012_);
  and (_11591_, _11495_, _11477_);
  nor (_11592_, _11591_, _11590_);
  not (_11593_, _11592_);
  not (_11594_, _11547_);
  and (_11595_, _11486_, _07015_);
  nor (_11596_, _11531_, _11595_);
  and (_11597_, _11596_, _11594_);
  nor (_11598_, _11597_, _11478_);
  nor (_11599_, _11598_, _11593_);
  and (_11600_, _11599_, _11589_);
  and (_11601_, _11600_, _11573_);
  and (_11602_, _11601_, _11555_);
  nor (_11603_, _11602_, _06318_);
  not (_11604_, _11602_);
  and (_11605_, _11513_, _06363_);
  not (_11606_, _11605_);
  and (_11607_, _11477_, _11595_);
  or (_11608_, _11506_, _07009_);
  and (_11609_, _11608_, _11547_);
  nor (_11610_, _11609_, _11607_);
  and (_11611_, _11610_, _11606_);
  and (_11612_, _11611_, _11592_);
  and (_11613_, _11612_, _11566_);
  and (_11614_, _11613_, _11553_);
  nand (_11615_, _11614_, _11604_);
  and (_11617_, _11615_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_11618_, _11602_, _06318_);
  nor (_11619_, _11618_, _11603_);
  and (_11620_, _11619_, _11617_);
  nor (_11621_, _11620_, _11603_);
  nor (_11622_, _11621_, _07516_);
  and (_11623_, _11622_, _06302_);
  nor (_11624_, _11622_, _06302_);
  nor (_11625_, _11624_, _11623_);
  nor (_11626_, _11625_, _11475_);
  and (_11627_, _06319_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_11628_, _11627_, _11475_);
  nor (_11629_, _11628_, _11614_);
  or (_11630_, _11629_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_11631_, _11630_, _11626_);
  and (_10377_, _11631_, _05141_);
  and (_11633_, _05141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  not (_11634_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor (_11635_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_11636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_11637_, _11636_, _11635_);
  not (_11639_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_11640_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_11642_, _11640_, _11639_);
  and (_11643_, _11642_, _11637_);
  and (_11644_, _11643_, _11634_);
  and (_11646_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _05141_);
  and (_11647_, _11646_, _11644_);
  or (_10382_, _11647_, _11633_);
  nor (_11648_, _11644_, rst);
  or (_11649_, _07516_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_11650_, _11649_, _10340_);
  or (_10388_, _11650_, _11648_);
  not (_11651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_11652_, _06725_, _11651_);
  or (_11653_, _11652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_11654_, _11653_, _11458_);
  not (_11655_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_11656_, _06207_, _11655_);
  nand (_11657_, _11656_, _11458_);
  or (_11659_, _11657_, _06208_);
  and (_11660_, _11659_, _11654_);
  or (_11661_, _11660_, _11462_);
  nand (_11662_, _11462_, _06244_);
  and (_11663_, _11662_, _05141_);
  and (_10406_, _11663_, _11661_);
  and (_11665_, _05922_, _10407_);
  or (_11667_, _05209_, _05186_);
  nor (_11668_, _05287_, _08651_);
  and (_11669_, _11668_, _11667_);
  or (_11671_, _11669_, _11665_);
  and (_11672_, _11671_, _11458_);
  nor (_11673_, _06209_, _05287_);
  nand (_11674_, _11458_, _11673_);
  and (_11676_, _11674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_11678_, _11676_, _11462_);
  or (_11680_, _11678_, _11672_);
  or (_11681_, _11463_, _06004_);
  and (_11683_, _11681_, _05141_);
  and (_10409_, _11683_, _11680_);
  and (_11684_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_11685_, _11684_, _10380_);
  and (_11686_, _11685_, _11458_);
  not (_11687_, _11458_);
  or (_11689_, _11687_, _10375_);
  and (_11690_, _11689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_11691_, _11690_, _11462_);
  or (_11692_, _11691_, _11686_);
  or (_11693_, _11463_, _05522_);
  and (_11694_, _11693_, _05141_);
  and (_10412_, _11694_, _11692_);
  and (_11696_, _08283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_11698_, _11696_, _08281_);
  and (_11699_, _11698_, _11458_);
  nand (_11701_, _11458_, _05186_);
  and (_11702_, _11701_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_11704_, _11702_, _11462_);
  or (_11705_, _11704_, _11699_);
  nand (_11706_, _11462_, _06062_);
  and (_11707_, _11706_, _05141_);
  and (_10417_, _11707_, _11705_);
  and (_11708_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_11709_, _11708_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  or (_11710_, _11709_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_10458_, _11710_, _05141_);
  not (_11711_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_11712_, _08463_, _11711_);
  nor (_11713_, _06727_, _11711_);
  and (_11714_, _11713_, _08439_);
  and (_11715_, _11714_, _08457_);
  and (_11716_, _08453_, _08439_);
  and (_11718_, _11716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor (_11720_, _11716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor (_11721_, _11720_, _11718_);
  or (_11722_, _11721_, _08463_);
  or (_11723_, _11722_, _11715_);
  and (_11724_, _11723_, _11712_);
  and (_11725_, _06736_, _10407_);
  and (_11726_, _11725_, _06734_);
  nor (_11727_, _11726_, _08471_);
  and (_11728_, _11727_, _11724_);
  and (_11729_, _08478_, _06703_);
  and (_11730_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_11731_, _11730_, _11729_);
  or (_11732_, _11731_, _11728_);
  and (_10461_, _11732_, _05141_);
  not (_11733_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_11734_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor (_11735_, _11734_, _11733_);
  and (_11736_, _11734_, _11733_);
  nor (_11737_, _11736_, _11735_);
  not (_11738_, _11737_);
  and (_11739_, _11738_, _10458_);
  nor (_11740_, _11735_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_11741_, _11735_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_11742_, _11741_, _11740_);
  nor (_11743_, _11708_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_11744_, _11743_, _11709_);
  or (_11745_, _11744_, _11734_);
  and (_11746_, _11745_, _11742_);
  and (_10476_, _11746_, _11739_);
  nor (_11747_, _08478_, _08471_);
  and (_11748_, _11718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_11749_, _11748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand (_11750_, _11749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_11751_, _11749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_11752_, _11751_, _11750_);
  not (_11753_, _06727_);
  and (_11754_, _08439_, _11753_);
  and (_11755_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_11756_, _11755_, _08457_);
  or (_11757_, _11756_, _08463_);
  or (_11758_, _11757_, _11752_);
  or (_11759_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_11760_, _11759_, _11758_);
  and (_11761_, _11760_, _11747_);
  nor (_11762_, _08479_, _06062_);
  and (_11763_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_11764_, _11763_, _11762_);
  or (_11765_, _11764_, _11761_);
  and (_10489_, _11765_, _05141_);
  nor (_11766_, _11748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_11767_, _11766_, _11749_);
  or (_11768_, _11767_, _08463_);
  and (_11769_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_11770_, _11769_, _08457_);
  or (_11771_, _11770_, _11768_);
  or (_11772_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_11773_, _11772_, _11771_);
  and (_11774_, _11773_, _11747_);
  and (_11775_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_11776_, _11775_, _11774_);
  nor (_11777_, _08479_, _05560_);
  or (_11778_, _11777_, _11776_);
  and (_10492_, _11778_, _05141_);
  and (_11779_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_11780_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_11781_, _11718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_11782_, _11781_, _11748_);
  or (_11783_, _11782_, _08463_);
  and (_11784_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_11785_, _11784_, _08457_);
  or (_11786_, _11785_, _11783_);
  and (_11787_, _11786_, _11780_);
  and (_11788_, _11787_, _11727_);
  not (_11789_, _11726_);
  nor (_11790_, _11789_, _06178_);
  or (_11791_, _11790_, _11788_);
  or (_11792_, _11791_, _11779_);
  and (_10499_, _11792_, _05141_);
  and (_11793_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _07611_);
  and (_11794_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_11795_, _11794_, _11793_);
  and (_10503_, _11795_, _05141_);
  and (_11796_, _06520_, _06468_);
  and (_11797_, _11796_, _06442_);
  and (_11798_, _06269_, _06317_);
  and (_11799_, _11798_, _06296_);
  and (_11800_, _11799_, _06332_);
  and (_11801_, _06493_, _06410_);
  and (_11802_, _11801_, _11800_);
  and (_11803_, _06385_, _06358_);
  and (_11804_, _11803_, _11802_);
  and (_10510_, _11804_, _11797_);
  and (_11805_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_11806_, _08478_, _06004_);
  or (_11807_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_11808_, _08453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_11809_, _11808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_11810_, _11809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_11811_, _11810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_11812_, _11811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_11813_, _11812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_11814_, _11813_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_11815_, _11814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_11816_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_11817_, _11816_, _11815_);
  and (_11818_, _08455_, _08439_);
  or (_11819_, _11818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand (_11820_, _11818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_11821_, _11820_, _11819_);
  or (_11822_, _11821_, _08463_);
  or (_11823_, _11822_, _11817_);
  and (_11824_, _11823_, _11807_);
  and (_11825_, _11824_, _11747_);
  or (_11826_, _11825_, _11806_);
  or (_11827_, _11826_, _11805_);
  and (_10529_, _11827_, _05141_);
  nand (_11828_, _11726_, _06244_);
  and (_11829_, _08456_, _08439_);
  and (_11830_, _11829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_11831_, _11829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_11832_, _11831_, _11830_);
  and (_11833_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_11834_, _11833_, _08439_);
  and (_11835_, _11834_, _08457_);
  or (_11836_, _11835_, _08463_);
  or (_11837_, _11836_, _11832_);
  nor (_11838_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_11839_, _11838_, _08471_);
  and (_11840_, _11839_, _11837_);
  and (_11841_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_11842_, _11841_, _08478_);
  or (_11843_, _11842_, _11840_);
  and (_11844_, _11843_, _05141_);
  and (_10540_, _11844_, _11828_);
  not (_11845_, _05522_);
  and (_11846_, _05256_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_11847_, _10355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_11848_, _11847_, _10387_);
  and (_11849_, _11848_, _10341_);
  nor (_11850_, _11849_, _11846_);
  and (_11851_, _06531_, _05197_);
  not (_11852_, _11851_);
  and (_11853_, _06365_, _05286_);
  nand (_11854_, _05266_, _05287_);
  nor (_11855_, _11854_, _11853_);
  and (_11856_, _11855_, _11852_);
  and (_11857_, _11856_, _05242_);
  and (_11858_, _11857_, _05297_);
  nand (_11859_, _10355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_11860_, _10355_, _06062_);
  nand (_11861_, _11860_, _11859_);
  or (_11862_, _11861_, _05172_);
  and (_11863_, _11860_, _11859_);
  or (_11864_, _11863_, _05173_);
  and (_11865_, _11864_, _11862_);
  and (_11866_, _11865_, _11858_);
  and (_11867_, _11866_, _11850_);
  nand (_11868_, _11867_, _05960_);
  not (_11869_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or (_11870_, _11847_, _10387_);
  and (_11871_, _11863_, _06365_);
  nand (_11872_, _11871_, _11870_);
  or (_11873_, _11872_, _11869_);
  and (_11874_, _11861_, _06365_);
  and (_11875_, _11874_, _11848_);
  nand (_11876_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_11877_, _11876_, _11873_);
  and (_11878_, _11863_, _06531_);
  and (_11879_, _11878_, _11870_);
  nand (_11880_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_11881_, _11878_, _11848_);
  nand (_11882_, _11881_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_11883_, _11882_, _11880_);
  and (_11884_, _11883_, _11877_);
  not (_11885_, _11867_);
  and (_11886_, _11861_, _06531_);
  and (_11887_, _11886_, _11870_);
  nand (_11888_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_11889_, _11874_, _11870_);
  nand (_11891_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_11892_, _11891_, _11888_);
  and (_11893_, _11886_, _11848_);
  nand (_11894_, _11893_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_11895_, _11871_, _11848_);
  nand (_11896_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_11897_, _11896_, _11894_);
  and (_11898_, _11897_, _11892_);
  and (_11899_, _11898_, _11885_);
  nand (_11900_, _11899_, _11884_);
  and (_11901_, _11900_, _11868_);
  and (_10555_, _11901_, _05141_);
  and (_10557_, _11870_, _05141_);
  not (_11902_, _08471_);
  or (_11903_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_11904_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_11905_, _11904_, _08439_);
  and (_11906_, _11905_, _08457_);
  nand (_11907_, _08448_, _08439_);
  nor (_11908_, _11907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_11909_, _11907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_11910_, _11909_, _08463_);
  or (_11911_, _11910_, _11908_);
  or (_11912_, _11911_, _11906_);
  nand (_11913_, _11912_, _11903_);
  nand (_11914_, _11913_, _11902_);
  nand (_11915_, _08471_, _06062_);
  and (_11916_, _11915_, _11914_);
  or (_11917_, _11916_, _11726_);
  or (_11918_, _11789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_11919_, _11918_, _05141_);
  and (_10570_, _11919_, _11917_);
  nor (_11920_, _11902_, _06244_);
  and (_11922_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_11923_, _11922_, _08439_);
  and (_11924_, _11923_, _08457_);
  nand (_11925_, _08451_, _08439_);
  nor (_11926_, _11925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_11927_, _11925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_11928_, _11927_, _08463_);
  or (_11929_, _11928_, _11926_);
  or (_11930_, _11929_, _11924_);
  nor (_11931_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_11932_, _11931_, _08471_);
  and (_11933_, _11932_, _11930_);
  or (_11934_, _11933_, _11726_);
  or (_11935_, _11934_, _11920_);
  or (_11936_, _11789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_11937_, _11936_, _05141_);
  and (_10575_, _11937_, _11935_);
  and (_11938_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_11939_, _11938_, _08439_);
  and (_11940_, _11939_, _08457_);
  and (_11941_, _08450_, _08439_);
  or (_11942_, _11941_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_11943_, _11942_, _11925_);
  or (_11944_, _11943_, _08463_);
  or (_11945_, _11944_, _11940_);
  nor (_11946_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor (_11948_, _11946_, _08471_);
  and (_11949_, _11948_, _11945_);
  and (_11950_, _08471_, _06004_);
  or (_11951_, _11950_, _08478_);
  or (_11952_, _11951_, _11949_);
  or (_11953_, _08479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_11954_, _11953_, _05141_);
  and (_10583_, _11954_, _11952_);
  and (_11955_, _05651_, _05209_);
  and (_11956_, _11955_, _06734_);
  and (_11957_, _11956_, _05925_);
  or (_11958_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_11959_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_11960_, _11959_, _08439_);
  and (_11961_, _11960_, _08457_);
  and (_11962_, _08449_, _08439_);
  nor (_11963_, _11962_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_11964_, _11963_, _11941_);
  or (_11965_, _11964_, _08463_);
  or (_11966_, _11965_, _11961_);
  nand (_11967_, _11966_, _11958_);
  nor (_11969_, _11967_, _11957_);
  and (_11970_, _11957_, _05522_);
  or (_11971_, _11970_, _11969_);
  or (_11972_, _11971_, _11726_);
  or (_11973_, _11789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_11974_, _11973_, _05141_);
  and (_10610_, _11974_, _11972_);
  and (_11976_, _05141_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_11977_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_11978_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_11980_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_11981_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_11982_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_11983_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_11984_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_11986_, _11985_, _11983_);
  and (_11988_, _11986_, _11984_);
  nor (_11989_, _11988_, _11983_);
  nor (_11990_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_11991_, _11990_, _11982_);
  not (_11992_, _11991_);
  nor (_11994_, _11992_, _11989_);
  nor (_11996_, _11994_, _11982_);
  not (_11997_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_11998_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_11999_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_12000_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_12001_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_12003_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_12004_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_12005_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_12006_, _12005_, _12004_);
  and (_12007_, _12006_, _12003_);
  and (_12009_, _12007_, _12001_);
  and (_12010_, _12009_, _12000_);
  and (_12011_, _12010_, _11999_);
  and (_12012_, _12011_, _11998_);
  and (_12014_, _12012_, _11997_);
  and (_12015_, _12014_, _11996_);
  and (_12017_, _12015_, _11981_);
  and (_12019_, _12017_, _11980_);
  and (_12020_, _12019_, _11978_);
  and (_12021_, _12020_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_12022_, _12020_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_12023_, _12022_, _12021_);
  nor (_12024_, _12019_, _11978_);
  nor (_12025_, _12024_, _12020_);
  nor (_12026_, _12017_, _11980_);
  nor (_12027_, _12026_, _12019_);
  nor (_12028_, _12015_, _11981_);
  nor (_12029_, _12028_, _12017_);
  not (_12030_, _12029_);
  and (_12031_, _12012_, _11996_);
  nor (_12032_, _12031_, _11997_);
  nor (_12033_, _12032_, _12015_);
  not (_12034_, _12033_);
  and (_12035_, _12011_, _11996_);
  nor (_12036_, _12035_, _11998_);
  nor (_12037_, _12036_, _12031_);
  not (_12038_, _12037_);
  and (_12039_, _12010_, _11996_);
  nor (_12040_, _12039_, _11999_);
  nor (_12041_, _12040_, _12035_);
  not (_12042_, _12041_);
  and (_12043_, _11996_, _12009_);
  nor (_12044_, _12043_, _12000_);
  nor (_12045_, _12044_, _12039_);
  not (_12046_, _12045_);
  and (_12047_, _11996_, _12007_);
  nor (_12048_, _12047_, _12001_);
  nor (_12049_, _12048_, _12043_);
  not (_12050_, _12049_);
  and (_12051_, _11996_, _12006_);
  nor (_12052_, _12051_, _12003_);
  or (_12053_, _12052_, _12047_);
  not (_12054_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  not (_12055_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_12056_, _11996_, _12055_);
  and (_12057_, _12056_, _12054_);
  nor (_12059_, _12057_, _12004_);
  or (_12060_, _12059_, _12051_);
  nor (_12061_, _11996_, _12055_);
  nor (_12062_, _12061_, _12056_);
  not (_12063_, _12062_);
  nor (_12064_, _11986_, _11984_);
  nor (_12065_, _12064_, _11988_);
  nand (_12066_, _12065_, _11604_);
  not (_12068_, _12066_);
  nor (_12069_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_12071_, _12069_, _11984_);
  and (_12072_, _12071_, _11615_);
  or (_12074_, _12065_, _11604_);
  and (_12075_, _12074_, _12066_);
  and (_12077_, _12075_, _12072_);
  or (_12078_, _12077_, _12068_);
  and (_12079_, _11992_, _11989_);
  nor (_12081_, _12079_, _11994_);
  and (_12083_, _12081_, _12078_);
  and (_12084_, _12083_, _12063_);
  nor (_12086_, _12056_, _12054_);
  or (_12087_, _12086_, _12057_);
  and (_12088_, _12087_, _12084_);
  and (_12089_, _12088_, _12060_);
  and (_12091_, _12089_, _12053_);
  and (_12092_, _12091_, _12050_);
  and (_12093_, _12092_, _12046_);
  and (_12094_, _12093_, _12042_);
  and (_12095_, _12094_, _12038_);
  and (_12096_, _12095_, _12034_);
  nand (_12097_, _12096_, _12030_);
  or (_12099_, _12097_, _12027_);
  or (_12100_, _12099_, _12025_);
  or (_12101_, _12100_, _12023_);
  nand (_12103_, _12100_, _12023_);
  and (_12105_, _12103_, _12101_);
  or (_12106_, _12105_, _07135_);
  or (_12107_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_12108_, rst, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_12110_, _12108_, _12107_);
  and (_12111_, _12110_, _12106_);
  or (_10640_, _12111_, _11977_);
  and (_12112_, _06782_, _06550_);
  and (_12114_, _08333_, _06544_);
  nor (_12115_, _12114_, _12112_);
  and (_12117_, _06760_, _06565_);
  and (_12118_, _06767_, _06550_);
  nor (_12120_, _12118_, _12117_);
  nand (_12121_, _12120_, _12115_);
  nor (_12123_, _12121_, _07040_);
  and (_12124_, _06566_, _06550_);
  or (_12126_, _12124_, _06559_);
  nor (_12127_, _12126_, _07056_);
  or (_12129_, _07047_, _06990_);
  and (_12130_, _06544_, _06572_);
  or (_12131_, _12130_, _07073_);
  nor (_12132_, _12131_, _12129_);
  and (_12133_, _12132_, _12127_);
  nand (_12135_, _06768_, _06760_);
  and (_12136_, _06760_, _07053_);
  or (_12138_, _12136_, _06994_);
  and (_12139_, _11428_, _06760_);
  nor (_12141_, _12139_, _12138_);
  and (_12142_, _12141_, _12135_);
  and (_12144_, _06760_, _06529_);
  or (_12145_, _07067_, _07044_);
  nor (_12147_, _12145_, _12144_);
  nor (_12148_, _07063_, _06799_);
  and (_12149_, _12148_, _11438_);
  and (_12150_, _12149_, _12147_);
  and (_12151_, _12150_, _12142_);
  and (_12152_, _12151_, _12133_);
  nand (_12153_, _12152_, _12123_);
  nand (_12155_, _12153_, _06821_);
  nor (_12156_, _11451_, _08341_);
  nand (_12158_, _12156_, _12155_);
  nand (_12159_, _12158_, _05143_);
  and (_12161_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_12162_, _12161_);
  nand (_12164_, _12162_, _12159_);
  not (_12165_, _11425_);
  or (_12166_, _11456_, _12165_);
  or (_12167_, _12166_, _12164_);
  or (_12168_, _12167_, _11848_);
  and (_12169_, _12162_, _12159_);
  or (_12170_, _12166_, _12169_);
  nor (_12171_, _06271_, _05312_);
  nor (_12172_, _06308_, _06427_);
  nor (_12173_, _06314_, _06429_);
  nor (_12174_, _12173_, _12172_);
  and (_12175_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_12176_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_12177_, _12176_, _12175_);
  and (_12178_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_12179_, _06320_, _06438_);
  nor (_12181_, _12179_, _12178_);
  and (_12182_, _12181_, _12177_);
  and (_12184_, _12182_, _12174_);
  nor (_12185_, _12184_, _07135_);
  nor (_12186_, _12185_, _12171_);
  or (_12188_, _12186_, _12170_);
  and (_12189_, _12188_, _12168_);
  and (_12191_, _12169_, _11456_);
  and (_12192_, _12191_, _11425_);
  and (_12193_, _11867_, _11845_);
  not (_12194_, _11872_);
  nand (_12195_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nand (_12196_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_12197_, _12196_, _12195_);
  nand (_12199_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nand (_12200_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_12201_, _12200_, _12199_);
  and (_12202_, _12201_, _12197_);
  or (_12204_, _11863_, _06365_);
  or (_12205_, _12204_, _11870_);
  or (_12207_, _12205_, _08129_);
  nand (_12208_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_12209_, _12208_, _12207_);
  nand (_12211_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nand (_12213_, _11878_, _11848_);
  or (_12214_, _12213_, _06719_);
  and (_12215_, _12214_, _12211_);
  and (_12216_, _12215_, _12209_);
  and (_12217_, _12216_, _11885_);
  and (_12219_, _12217_, _12202_);
  nor (_12220_, _12219_, _12193_);
  nand (_12221_, _12220_, _12192_);
  or (_12222_, _11456_, _11425_);
  nand (_12223_, _12164_, _11456_);
  nor (_12224_, _12223_, _12165_);
  and (_12225_, _06621_, _05288_);
  and (_12226_, _12225_, _05522_);
  nand (_12228_, _06621_, _05288_);
  or (_12229_, _12228_, _06062_);
  or (_12230_, _12225_, _05152_);
  nand (_12231_, _12230_, _12229_);
  or (_12232_, _12225_, _05153_);
  or (_12233_, _12228_, _05560_);
  nand (_12234_, _12233_, _12232_);
  nand (_12235_, _12228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  or (_12236_, _12228_, _06178_);
  and (_12237_, _12236_, _12235_);
  not (_12238_, _12237_);
  not (_12239_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  or (_12240_, _12225_, _05192_);
  or (_12241_, _12228_, _05604_);
  nand (_12243_, _12241_, _12240_);
  or (_12244_, _12243_, _12239_);
  or (_12245_, _12244_, _12238_);
  or (_12247_, _12245_, _12234_);
  nor (_12248_, _12247_, _12231_);
  and (_12249_, _12228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_12250_, _12249_, _12226_);
  and (_12251_, _12250_, _12248_);
  nor (_12252_, _12250_, _12248_);
  or (_12253_, _12252_, _12251_);
  nand (_12254_, _12253_, _05243_);
  nand (_12255_, _12254_, _05246_);
  and (_12256_, _12255_, _12228_);
  or (_12257_, _12256_, _12226_);
  nand (_12258_, _12257_, _12224_);
  and (_12259_, _12258_, _12222_);
  and (_12260_, _12259_, _12221_);
  and (_12261_, _12260_, _12189_);
  or (_12262_, _12261_, _10341_);
  nand (_12263_, _12260_, _12189_);
  or (_12264_, _12263_, _05256_);
  and (_12265_, _12264_, _12262_);
  and (_12266_, _11456_, _12165_);
  nand (_12267_, _12266_, _12164_);
  or (_12268_, _12170_, _07514_);
  nor (_12269_, _11885_, _06004_);
  nand (_12270_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nand (_12271_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_12272_, _12271_, _12270_);
  nand (_12273_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_12274_, _12205_, _08237_);
  and (_12275_, _12274_, _12273_);
  and (_12276_, _12275_, _12272_);
  or (_12277_, _11872_, _07096_);
  nand (_12278_, _11881_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_12279_, _12278_, _12277_);
  nand (_12280_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nand (_12281_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_12282_, _12281_, _12280_);
  and (_12283_, _12282_, _12279_);
  and (_12285_, _12283_, _11885_);
  and (_12286_, _12285_, _12276_);
  or (_12287_, _12286_, _12269_);
  not (_12288_, _12287_);
  nand (_12289_, _12288_, _12192_);
  and (_12290_, _12289_, _12268_);
  or (_12291_, _12223_, _12165_);
  and (_12292_, _12225_, _06004_);
  not (_12293_, _12292_);
  and (_12294_, _12228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_12296_, _12294_, _12292_);
  nand (_12297_, _12296_, _12251_);
  or (_12299_, _12296_, _12251_);
  and (_12300_, _12299_, _12297_);
  or (_12301_, _12300_, _05159_);
  and (_12302_, _12301_, _05259_);
  or (_12303_, _12302_, _12225_);
  and (_12304_, _12303_, _12293_);
  or (_12305_, _12304_, _12291_);
  or (_12306_, _12222_, _12164_);
  and (_12308_, _12306_, _12305_);
  and (_12309_, _12308_, _12290_);
  and (_12310_, _12309_, _12267_);
  and (_12312_, _12310_, _05280_);
  nand (_12313_, _12309_, _12267_);
  and (_12314_, _12313_, _05266_);
  nor (_12315_, _12314_, _12312_);
  and (_12317_, _12315_, _12265_);
  and (_12318_, _12247_, _12231_);
  nor (_12319_, _12318_, _12248_);
  nor (_12320_, _12319_, _05159_);
  not (_12321_, _12320_);
  nand (_12322_, _12321_, _05162_);
  nand (_12323_, _12322_, _12228_);
  nand (_12325_, _12323_, _12229_);
  nand (_12326_, _12325_, _12224_);
  or (_12327_, _12167_, _11863_);
  nand (_12329_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nand (_12330_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_12331_, _12330_, _12329_);
  nand (_12332_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nand (_12333_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_12335_, _12333_, _12332_);
  and (_12336_, _12335_, _12331_);
  or (_12338_, _12205_, _08076_);
  or (_12339_, _12213_, _08487_);
  and (_12340_, _12339_, _12338_);
  nand (_12341_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nand (_12343_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_12344_, _12343_, _12341_);
  and (_12346_, _12344_, _12340_);
  and (_12347_, _12346_, _11885_);
  nand (_12349_, _12347_, _12336_);
  nand (_12350_, _11867_, _06062_);
  and (_12351_, _12350_, _12349_);
  nand (_12352_, _12351_, _12192_);
  nor (_12354_, _06271_, _05385_);
  nor (_12355_, _06308_, _06403_);
  nor (_12356_, _06314_, _06395_);
  nor (_12357_, _12356_, _12355_);
  and (_12358_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_12359_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_12361_, _12359_, _12358_);
  nor (_12362_, _06304_, _06399_);
  nor (_12363_, _06320_, _06406_);
  nor (_12364_, _12363_, _12362_);
  and (_12365_, _12364_, _12361_);
  and (_12366_, _12365_, _12357_);
  nor (_12367_, _12366_, _07135_);
  nor (_12368_, _12367_, _12354_);
  or (_12369_, _12368_, _12170_);
  and (_12370_, _12369_, _12352_);
  and (_12371_, _12370_, _12327_);
  and (_12372_, _12371_, _12326_);
  or (_12373_, _12372_, _05173_);
  nand (_12374_, _12371_, _12326_);
  or (_12375_, _12374_, _05172_);
  and (_12376_, _12375_, _12373_);
  and (_12377_, _12225_, _05960_);
  not (_12378_, _12297_);
  nor (_12379_, _12228_, _06244_);
  and (_12380_, _12228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_12381_, _12380_, _12379_);
  and (_12382_, _12381_, _12378_);
  and (_12383_, _12228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand (_12384_, _12383_, _12382_);
  or (_12385_, _12383_, _12382_);
  and (_12386_, _12385_, _05243_);
  nand (_12387_, _12386_, _12384_);
  and (_12388_, _12228_, _05232_);
  and (_12389_, _12388_, _12387_);
  nor (_12390_, _12389_, _12377_);
  nand (_12391_, _12390_, _12224_);
  and (_12392_, _11901_, _12192_);
  and (_12393_, _12223_, _12165_);
  nor (_12394_, _12393_, _12392_);
  or (_12395_, _12170_, _07137_);
  and (_12396_, _12395_, _12267_);
  and (_12397_, _12396_, _12394_);
  and (_12398_, _12397_, _12391_);
  nand (_12399_, _12398_, _05241_);
  or (_12400_, _12398_, _05241_);
  and (_12401_, _12400_, _12399_);
  nand (_12402_, _12381_, _12378_);
  or (_12403_, _12381_, _12378_);
  nand (_12404_, _12403_, _12402_);
  nand (_12405_, _12404_, _05243_);
  nand (_12407_, _12405_, _05218_);
  and (_12408_, _12407_, _12228_);
  or (_12409_, _12408_, _12379_);
  nand (_12410_, _12409_, _12224_);
  and (_12411_, _12267_, _12222_);
  nor (_12412_, _06271_, _05692_);
  nor (_12413_, _06308_, _06514_);
  nor (_12414_, _06314_, _06510_);
  nor (_12415_, _12414_, _12413_);
  and (_12416_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_12417_, _06320_, _06516_);
  nor (_12418_, _12417_, _12416_);
  and (_12419_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_12420_, _06304_, _06508_);
  nor (_12421_, _12420_, _12419_);
  and (_12422_, _12421_, _12418_);
  and (_12423_, _12422_, _12415_);
  nor (_12424_, _12423_, _07135_);
  nor (_12425_, _12424_, _12412_);
  or (_12426_, _12425_, _12170_);
  nand (_12427_, _11867_, _06244_);
  nand (_12428_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nand (_12429_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_12430_, _12429_, _12428_);
  nand (_12431_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nand (_12432_, _11881_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_12433_, _12432_, _12431_);
  and (_12434_, _12433_, _12430_);
  nand (_12435_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nand (_12436_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_12437_, _12436_, _12435_);
  nand (_12438_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nand (_12439_, _11893_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_12440_, _12439_, _12438_);
  and (_12441_, _12440_, _12437_);
  and (_12442_, _12441_, _11885_);
  nand (_12443_, _12442_, _12434_);
  and (_12444_, _12443_, _12427_);
  nand (_12445_, _12444_, _12192_);
  and (_12446_, _12445_, _12426_);
  and (_12447_, _12446_, _12411_);
  nand (_12448_, _12447_, _12410_);
  and (_12449_, _12448_, _05227_);
  and (_12450_, _12447_, _12410_);
  and (_12451_, _12450_, _05228_);
  nor (_12452_, _12451_, _12449_);
  and (_12453_, _12452_, _12401_);
  and (_12454_, _12453_, _12376_);
  and (_12455_, _12454_, _12317_);
  nor (_12456_, _12243_, _12239_);
  and (_12457_, _12243_, _12239_);
  nor (_12458_, _12457_, _12456_);
  nor (_12459_, _12458_, _05159_);
  nor (_12460_, _12459_, _05193_);
  nor (_12461_, _12460_, _12225_);
  not (_12462_, _12461_);
  and (_12463_, _12462_, _12241_);
  or (_12464_, _12463_, _12291_);
  or (_12465_, _12167_, _06365_);
  nand (_12466_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  or (_12467_, _12213_, _09779_);
  and (_12468_, _12467_, _12466_);
  nand (_12469_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or (_12470_, _12205_, _05621_);
  and (_12471_, _12470_, _12469_);
  and (_12472_, _12471_, _12468_);
  nand (_12473_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nand (_12474_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_12475_, _12474_, _12473_);
  nand (_12476_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nand (_12477_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_12478_, _12477_, _12476_);
  and (_12479_, _12478_, _12475_);
  and (_12480_, _12479_, _11885_);
  nand (_12481_, _12480_, _12472_);
  nand (_12482_, _11867_, _05604_);
  and (_12483_, _12482_, _12481_);
  nand (_12484_, _12483_, _12192_);
  nor (_12485_, _06271_, _05406_);
  nor (_12486_, _06308_, _06351_);
  nor (_12487_, _06314_, _06343_);
  nor (_12488_, _12487_, _12486_);
  and (_12489_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_12490_, _06320_, _06353_);
  nor (_12491_, _12490_, _12489_);
  and (_12492_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_12493_, _06304_, _06347_);
  nor (_12494_, _12493_, _12492_);
  and (_12495_, _12494_, _12491_);
  and (_12496_, _12495_, _12488_);
  nor (_12497_, _12496_, _07135_);
  nor (_12498_, _12497_, _12485_);
  or (_12499_, _12498_, _12170_);
  and (_12500_, _12499_, _12484_);
  and (_12501_, _12500_, _12465_);
  and (_12502_, _12501_, _12464_);
  or (_12503_, _12502_, _05197_);
  nand (_12504_, _12501_, _12464_);
  or (_12505_, _12504_, _05286_);
  nand (_12506_, _12505_, _12503_);
  and (_12507_, _12506_, _05646_);
  and (_12508_, _12244_, _12238_);
  not (_12509_, _12508_);
  and (_12510_, _12509_, _12245_);
  nor (_12511_, _12510_, _05159_);
  nor (_12512_, _12511_, _05200_);
  nor (_12513_, _12512_, _12225_);
  not (_12514_, _12513_);
  and (_12515_, _12514_, _12236_);
  or (_12516_, _12515_, _12291_);
  nand (_12517_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nand (_12518_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_12519_, _12518_, _12517_);
  nand (_12520_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nand (_12521_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_12522_, _12521_, _12520_);
  and (_12523_, _12522_, _12519_);
  nand (_12524_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nand (_12525_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_12526_, _12525_, _12524_);
  or (_12527_, _12205_, _08155_);
  nand (_12528_, _11881_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_12529_, _12528_, _12527_);
  and (_12530_, _12529_, _12526_);
  and (_12531_, _12530_, _11885_);
  nand (_12532_, _12531_, _12523_);
  nand (_12533_, _11867_, _06178_);
  and (_12534_, _12533_, _12532_);
  nand (_12535_, _12534_, _12192_);
  nor (_12537_, _06271_, _05430_);
  nor (_12538_, _06308_, _06301_);
  nor (_12539_, _06314_, _06306_);
  nor (_12540_, _12539_, _12538_);
  and (_12541_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_12542_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_12543_, _12542_, _12541_);
  nor (_12544_, _06304_, _06324_);
  nor (_12545_, _06320_, _06311_);
  nor (_12546_, _12545_, _12544_);
  and (_12547_, _12546_, _12543_);
  and (_12548_, _12547_, _12540_);
  nor (_12549_, _12548_, _07135_);
  nor (_12550_, _12549_, _12537_);
  or (_12551_, _12550_, _12170_);
  and (_12552_, _12551_, _12535_);
  nand (_12553_, _12266_, _12169_);
  or (_12554_, _12167_, _06339_);
  and (_12555_, _12554_, _12553_);
  and (_12556_, _12555_, _12552_);
  and (_12557_, _12556_, _12516_);
  and (_12558_, _12557_, _05274_);
  nand (_12559_, _12556_, _12516_);
  and (_12560_, _12559_, _05208_);
  nor (_12561_, _12560_, _12558_);
  and (_12562_, _12245_, _12234_);
  not (_12563_, _12562_);
  and (_12564_, _12563_, _12247_);
  nor (_12565_, _12564_, _05159_);
  nor (_12566_, _12565_, _05178_);
  nor (_12567_, _12566_, _12225_);
  not (_12568_, _12567_);
  and (_12569_, _12568_, _12233_);
  or (_12570_, _12569_, _12291_);
  nand (_12571_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nand (_12572_, _11881_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_12573_, _12572_, _12571_);
  nand (_12574_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_12575_, _12205_, _08132_);
  and (_12576_, _12575_, _12574_);
  and (_12577_, _12576_, _12573_);
  nand (_12578_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nand (_12579_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_12580_, _12579_, _12578_);
  nand (_12581_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nand (_12582_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_12583_, _12582_, _12581_);
  and (_12584_, _12583_, _12580_);
  and (_12585_, _12584_, _11885_);
  and (_12586_, _12585_, _12577_);
  and (_12587_, _11867_, _05560_);
  nor (_12588_, _12587_, _12586_);
  nand (_12589_, _12588_, _12192_);
  or (_12590_, _12167_, _06533_);
  nor (_12591_, _06271_, _05447_);
  nor (_12592_, _06308_, _06376_);
  nor (_12593_, _06314_, _06374_);
  nor (_12594_, _12593_, _12592_);
  and (_12595_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_12596_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_12597_, _12596_, _12595_);
  nor (_12598_, _06304_, _06379_);
  nor (_12599_, _06320_, _06370_);
  nor (_12600_, _12599_, _12598_);
  and (_12601_, _12600_, _12597_);
  and (_12602_, _12601_, _12594_);
  nor (_12603_, _12602_, _07135_);
  nor (_12604_, _12603_, _12591_);
  or (_12605_, _12604_, _12170_);
  and (_12606_, _12605_, _12590_);
  and (_12607_, _12606_, _12589_);
  and (_12608_, _12607_, _12570_);
  or (_12609_, _12608_, _05186_);
  nand (_12610_, _12607_, _12570_);
  or (_12611_, _12610_, _06007_);
  nand (_12612_, _12611_, _12609_);
  and (_12613_, _12612_, _12561_);
  and (_12614_, _12613_, _12507_);
  and (_12615_, _12614_, _12455_);
  and (_12616_, _05241_, _05295_);
  nand (_12617_, _12616_, _12615_);
  not (_12618_, _08171_);
  and (_12619_, _11452_, _12618_);
  not (_12621_, _06846_);
  and (_12622_, _06563_, _06550_);
  nor (_12624_, _12622_, _06575_);
  not (_12625_, _12624_);
  and (_12626_, _12625_, _07088_);
  not (_12627_, _06558_);
  nor (_12628_, _12124_, _06554_);
  and (_12629_, _12628_, _12627_);
  and (_12631_, _12622_, _07088_);
  not (_12632_, _12631_);
  and (_12633_, _12632_, _12629_);
  nor (_12634_, _12633_, _06791_);
  nor (_12635_, _12634_, _12626_);
  and (_12636_, _06588_, _05824_);
  nand (_12637_, _12636_, _07322_);
  nor (_12638_, _12637_, _07233_);
  and (_12639_, _12638_, _07171_);
  and (_12640_, _12639_, _06662_);
  and (_12642_, _12640_, _07487_);
  and (_12643_, _12642_, _12635_);
  and (_12644_, _12643_, _12621_);
  and (_12645_, _07088_, _06563_);
  and (_12646_, _12645_, _06550_);
  not (_12647_, _12646_);
  nor (_12649_, _12646_, _12126_);
  nor (_12650_, _12649_, _06791_);
  and (_12651_, _12650_, _12647_);
  and (_12652_, _12651_, _05379_);
  nor (_12653_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_12654_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_12655_, _12654_, _12653_);
  nor (_12657_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_12658_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_12659_, _12658_, _12657_);
  and (_12660_, _12659_, _12655_);
  and (_12662_, _12660_, _11452_);
  and (_12663_, _12646_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_12664_, _12663_, _12662_);
  or (_12665_, _12664_, _12652_);
  nor (_12666_, _12665_, _12644_);
  and (_12667_, _08340_, _06450_);
  nor (_12668_, _12667_, _06559_);
  nor (_12669_, _12668_, _12666_);
  or (_12670_, _08334_, _06573_);
  and (_12671_, _06767_, _06755_);
  nor (_12672_, _12671_, _06981_);
  nor (_12673_, _06774_, _12124_);
  nand (_12674_, _12673_, _12672_);
  and (_12675_, _06570_, _06417_);
  and (_12676_, _08340_, _06449_);
  or (_12677_, _12676_, _12675_);
  or (_12678_, _12677_, _12674_);
  and (_12679_, _12678_, _12666_);
  or (_12680_, _12679_, _12670_);
  or (_12681_, _12680_, _12669_);
  and (_12682_, _12681_, _07088_);
  and (_12683_, _06552_, _06544_);
  nor (_12684_, _12683_, _06816_);
  nor (_12685_, _12684_, _08330_);
  nor (_12686_, _12685_, _11450_);
  not (_12687_, _12686_);
  nor (_12688_, _12687_, _12682_);
  nor (_12689_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_12690_, _12689_);
  nor (_12691_, _10354_, _12690_);
  and (_12692_, _12691_, _10376_);
  nor (_12693_, _12692_, _12632_);
  or (_12694_, _12693_, _12688_);
  nor (_12695_, _12694_, _12619_);
  nor (_12696_, _06735_, _06008_);
  and (_12697_, _12696_, _12455_);
  nand (_12698_, _12697_, _12651_);
  and (_12699_, _12698_, _12695_);
  and (_12700_, _12699_, _12617_);
  and (_12701_, _08334_, _07088_);
  and (_12702_, _12701_, _06975_);
  not (_12703_, _11451_);
  nor (_12704_, _12703_, _06875_);
  and (_12705_, _06821_, _06556_);
  and (_12706_, _12705_, _06550_);
  and (_12707_, _12683_, _06821_);
  or (_12708_, _12707_, _12706_);
  nor (_12709_, _12708_, _11451_);
  or (_12710_, _12674_, _06559_);
  nand (_12711_, _12710_, _07088_);
  and (_12712_, _12711_, _12709_);
  and (_12713_, _12712_, _12685_);
  nand (_12714_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_12715_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_12716_, _12715_, _12714_);
  nand (_12717_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand (_12718_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_12719_, \oc8051_top_1.oc8051_memory_interface1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_12720_, _12719_, _12718_);
  or (_12721_, _12720_, _12717_);
  or (_12723_, _12721_, _12716_);
  or (_12724_, _12723_, _05390_);
  or (_12725_, _12724_, _05317_);
  or (_12726_, _12725_, _05739_);
  or (_12727_, _12726_, _05699_);
  and (_12728_, _12727_, _05663_);
  nor (_12729_, _12727_, _05663_);
  nor (_12730_, _12729_, _12728_);
  and (_12731_, _12730_, _12713_);
  not (_12732_, _07137_);
  and (_12733_, _12707_, _12732_);
  nor (_12735_, _12701_, _12685_);
  nand (_12736_, _12735_, _12712_);
  or (_12737_, _08340_, _12675_);
  nor (_12739_, _12737_, _06774_);
  nand (_12740_, _12739_, _12672_);
  or (_12741_, _12670_, _12126_);
  or (_12742_, _12741_, _12740_);
  and (_12743_, _12742_, _07088_);
  or (_12744_, _12743_, _12706_);
  nor (_12745_, _12744_, _12736_);
  and (_12746_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_12747_, _12746_, _12733_);
  or (_12748_, _12747_, _12731_);
  or (_12749_, _12748_, _12704_);
  nor (_12750_, _12749_, _12702_);
  nand (_12751_, _12750_, _12700_);
  nand (_12752_, _12712_, _12732_);
  nor (_12753_, _06271_, _05658_);
  and (_12754_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12755_, _06308_, _06457_);
  nor (_12756_, _06320_, _06462_);
  nor (_12757_, _12756_, _12755_);
  and (_12758_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_12759_, _06314_, _06459_);
  nor (_12760_, _12759_, _12758_);
  and (_12761_, _12760_, _12757_);
  and (_12762_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_12763_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_12764_, _12763_, _12762_);
  and (_12765_, _12764_, _12761_);
  nor (_12766_, _12765_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12768_, _12766_, _12754_);
  nor (_12769_, _12768_, _07516_);
  nor (_12770_, _12769_, _12753_);
  or (_12771_, _12770_, _12712_);
  and (_12772_, _12771_, _12752_);
  not (_12773_, _12772_);
  nor (_12774_, \oc8051_top_1.oc8051_memory_interface1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_12775_, _12772_, _05665_);
  not (_12776_, _12425_);
  nand (_12777_, _12712_, _12776_);
  nor (_12778_, _06271_, _05694_);
  and (_12779_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12780_, _06308_, _06508_);
  nor (_12781_, _06320_, _06510_);
  nor (_12782_, _12781_, _12780_);
  and (_12783_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_12784_, _06314_, _06514_);
  nor (_12785_, _12784_, _12783_);
  and (_12786_, _12785_, _12782_);
  and (_12787_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_12789_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_12790_, _12789_, _12787_);
  and (_12792_, _12790_, _12786_);
  nor (_12793_, _12792_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12794_, _12793_, _12779_);
  nor (_12795_, _12794_, _07516_);
  nor (_12796_, _12795_, _12778_);
  or (_12797_, _12796_, _12712_);
  nand (_12798_, _12797_, _12777_);
  nand (_12799_, _12798_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_12800_, _12799_);
  nand (_12801_, _12772_, _05665_);
  and (_12802_, _12801_, _12775_);
  nand (_12803_, _12802_, _12800_);
  nand (_12804_, _12803_, _12775_);
  or (_12805_, _12798_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_12806_, _12805_, _12799_);
  and (_12807_, _12806_, _12802_);
  not (_12808_, _07514_);
  nand (_12809_, _12712_, _12808_);
  nor (_12810_, _06271_, _05734_);
  and (_12811_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12812_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor (_12813_, _06320_, _06484_);
  nor (_12814_, _12813_, _12812_);
  nor (_12816_, _06308_, _06482_);
  and (_12817_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_12818_, _12817_, _12816_);
  and (_12819_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_12820_, _06314_, _06487_);
  nor (_12821_, _12820_, _12819_);
  and (_12822_, _12821_, _12818_);
  and (_12823_, _12822_, _12814_);
  nor (_12824_, _12823_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12825_, _12824_, _12811_);
  nor (_12826_, _12825_, _07516_);
  nor (_12827_, _12826_, _12810_);
  or (_12828_, _12827_, _12712_);
  and (_12829_, _12828_, _12809_);
  or (_12830_, _12829_, _05742_);
  not (_12831_, _12186_);
  nand (_12832_, _12712_, _12831_);
  or (_12833_, _12712_, _07593_);
  nand (_12834_, _12833_, _12832_);
  nand (_12835_, _12834_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_12836_, _12829_, _05742_);
  and (_12837_, _12836_, _12830_);
  not (_12838_, _12837_);
  or (_12839_, _12838_, _12835_);
  nand (_12840_, _12839_, _12830_);
  and (_12841_, _12840_, _12807_);
  or (_12842_, _12841_, _12804_);
  not (_12843_, _12368_);
  and (_12844_, _12712_, _12843_);
  nor (_12845_, _12712_, _07572_);
  nor (_12846_, _12845_, _12844_);
  and (_12847_, _12846_, _05388_);
  nor (_12848_, _12846_, _05388_);
  not (_12849_, _12604_);
  nand (_12850_, _12712_, _12849_);
  or (_12851_, _12712_, _07550_);
  and (_12852_, _12851_, _12850_);
  nor (_12853_, _12852_, _05453_);
  not (_12855_, _12550_);
  nand (_12857_, _12712_, _12855_);
  nor (_12859_, _06271_, _05432_);
  and (_12860_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_12862_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor (_12863_, _06320_, _06306_);
  nor (_12864_, _12863_, _12862_);
  and (_12865_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nor (_12866_, _06314_, _06301_);
  nor (_12867_, _12866_, _12865_);
  and (_12868_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_12869_, _06308_, _06324_);
  nor (_12870_, _12869_, _12868_);
  and (_12871_, _12870_, _12867_);
  and (_12872_, _12871_, _12864_);
  nor (_12873_, _12872_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12874_, _12873_, _12860_);
  nor (_12875_, _12874_, _07516_);
  nor (_12876_, _12875_, _12859_);
  or (_12877_, _12876_, _12712_);
  and (_12878_, _12877_, _12857_);
  nor (_12879_, _12878_, _05438_);
  not (_12880_, _12498_);
  and (_12881_, _12712_, _12880_);
  nor (_12882_, _12712_, _07533_);
  or (_12883_, _12882_, _12881_);
  and (_12884_, _12883_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_12885_, _12879_);
  nand (_12886_, _12878_, _05438_);
  and (_12887_, _12886_, _12885_);
  and (_12888_, _12887_, _12884_);
  or (_12889_, _12888_, _12879_);
  not (_12890_, _12853_);
  nand (_12891_, _12852_, _05453_);
  and (_12892_, _12891_, _12890_);
  and (_12893_, _12892_, _12889_);
  or (_12894_, _12893_, _12853_);
  nor (_12895_, _12894_, _12848_);
  nor (_12896_, _12895_, _12847_);
  or (_12897_, _12834_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12898_, _12897_, _12835_);
  and (_12899_, _12837_, _12898_);
  and (_12900_, _12899_, _12807_);
  and (_12901_, _12900_, _12896_);
  or (_12902_, _12901_, _12842_);
  or (_12903_, _12902_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_12904_, _12903_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_12905_, _12904_, _12774_);
  and (_12906_, _12905_, _05317_);
  and (_12907_, _12906_, _05739_);
  nand (_12908_, _12907_, _05699_);
  nand (_12909_, _12908_, _12773_);
  and (_12910_, \oc8051_top_1.oc8051_memory_interface1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_12911_, _12910_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_12912_, _12902_, _12911_);
  nand (_12913_, _12912_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_12914_, _12913_, _05317_);
  nor (_12915_, _12914_, _05739_);
  nand (_12916_, _12915_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_12917_, _12916_, _12772_);
  nand (_12918_, _12917_, _12909_);
  nand (_12919_, _12918_, _05663_);
  or (_12920_, _12918_, _05663_);
  and (_12921_, _12920_, _12919_);
  not (_12922_, _12712_);
  or (_12923_, _12735_, _12922_);
  and (_12924_, _06821_, _06550_);
  and (_12926_, _12924_, _06556_);
  and (_12927_, _06778_, _06766_);
  nor (_12928_, _12927_, _11441_);
  nand (_12929_, _12928_, _12624_);
  or (_12930_, _12929_, _12670_);
  and (_12931_, _06767_, _06420_);
  and (_12932_, _06767_, _06760_);
  or (_12933_, _12932_, _12931_);
  or (_12934_, _12933_, _06981_);
  nor (_12935_, _12934_, _06988_);
  nand (_12936_, _12935_, _12629_);
  or (_12937_, _12936_, _12930_);
  and (_12938_, _12937_, _07088_);
  or (_12939_, _12938_, _12926_);
  and (_12940_, _12939_, _12923_);
  and (_12941_, _12940_, _12921_);
  or (_12942_, _12941_, _12751_);
  and (_12943_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_12944_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_12945_, _12944_, _12943_);
  and (_12946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_12947_, _12946_, _12945_);
  and (_12948_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_12949_, _12948_, _12947_);
  and (_12950_, _12949_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_12951_, _07619_);
  and (_12952_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_12953_, _12952_, _12951_);
  and (_12954_, _12953_, _12950_);
  and (_12955_, _12954_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_12956_, _12955_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_12957_, _12956_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_12958_, _12956_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_12959_, _12958_, _12957_);
  or (_12960_, _12959_, _12700_);
  and (_12961_, _12960_, _05141_);
  and (_10647_, _12961_, _12942_);
  and (_10656_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _05141_);
  nor (_12962_, _12089_, _12053_);
  nor (_12963_, _12962_, _12091_);
  or (_12964_, _12963_, _07135_);
  or (_12965_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_12966_, _12965_, _12108_);
  and (_12967_, _12966_, _12964_);
  and (_12968_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_10698_, _12968_, _12967_);
  or (_12969_, _12905_, _12772_);
  nand (_12970_, _12913_, _12772_);
  nand (_12971_, _12970_, _12969_);
  nand (_12972_, _12971_, _05317_);
  and (_12973_, _12744_, _12923_);
  or (_12974_, _12971_, _05317_);
  and (_12975_, _12974_, _12973_);
  and (_12976_, _12975_, _12972_);
  and (_12977_, _12701_, _07229_);
  and (_12978_, _12707_, _12831_);
  and (_12979_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12980_, \oc8051_top_1.oc8051_memory_interface1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_12981_, _12980_, _12979_);
  and (_12982_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_12983_, _12982_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_12984_, _12983_, _12911_);
  and (_12985_, _12984_, _12981_);
  and (_12986_, _12985_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_12987_, _12986_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_12988_, _12987_, _12725_);
  and (_12989_, _12988_, _12713_);
  or (_12990_, _12989_, _12978_);
  and (_12991_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_12992_, _12703_, _07259_);
  or (_12993_, _12992_, _12991_);
  or (_12995_, _12993_, _12990_);
  nor (_12996_, _12995_, _12977_);
  nand (_12997_, _12996_, _12700_);
  or (_12998_, _12997_, _12976_);
  and (_12999_, _12947_, _12951_);
  and (_13000_, _12999_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_13001_, _13000_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_13002_, _13001_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_13003_, _13002_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_13004_, _13003_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nand (_13005_, _13003_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_13006_, _13005_, _13004_);
  or (_13007_, _13006_, _12700_);
  and (_13008_, _13007_, _05141_);
  and (_10715_, _13008_, _12998_);
  nand (_13009_, _08396_, _05960_);
  and (_13010_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_13011_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_13012_, _13011_, _13010_);
  or (_13013_, _13012_, _08243_);
  and (_13014_, _13013_, _05141_);
  and (_10718_, _13014_, _13009_);
  and (_13015_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_13016_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or (_13017_, _13016_, _13015_);
  and (_10742_, _13017_, _05141_);
  or (_13018_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand (_13019_, _07619_, _06508_);
  and (_13020_, _13019_, _05141_);
  and (_10747_, _13020_, _13018_);
  or (_13022_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand (_13023_, _07619_, _06301_);
  and (_13024_, _13023_, _05141_);
  and (_10750_, _13024_, _13022_);
  and (_13025_, _08396_, _06283_);
  and (_13026_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_13027_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_13028_, _13027_, _13026_);
  nor (_13029_, _13028_, _08243_);
  not (_13031_, _05960_);
  and (_13032_, _08382_, _13031_);
  or (_13033_, _13032_, _13029_);
  or (_13034_, _13033_, _13025_);
  and (_10792_, _13034_, _05141_);
  and (_13035_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_13036_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_13037_, pc_log_change, _13036_);
  or (_13038_, _13037_, _13035_);
  and (_10800_, _13038_, _05141_);
  and (_13039_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_13040_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_13041_, _13040_, _13039_);
  nor (_13042_, _13041_, _08243_);
  or (_13043_, _08653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_13044_, _13043_, _08396_);
  or (_13045_, _13044_, _13042_);
  and (_10871_, _13045_, _05141_);
  and (_13046_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_13047_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  or (_13048_, _13047_, _13046_);
  and (_10887_, _13048_, _05141_);
  or (_13049_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand (_13050_, _07619_, _06376_);
  and (_13051_, _13050_, _05141_);
  and (_10890_, _13051_, _13049_);
  not (_13052_, _12700_);
  or (_13053_, _12883_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_13054_, _12884_);
  and (_13055_, _12973_, _13054_);
  and (_13056_, _13055_, _13053_);
  not (_13057_, _07496_);
  or (_13058_, _12745_, _12701_);
  and (_13059_, _13058_, _13057_);
  not (_13060_, _07533_);
  and (_13061_, _12707_, _13060_);
  and (_13062_, _12713_, _12880_);
  and (_13063_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_13064_, _13063_, _13062_);
  or (_13065_, _13064_, _13061_);
  or (_13066_, _13065_, _13059_);
  or (_13068_, _13066_, _13056_);
  or (_13069_, _13068_, _13052_);
  or (_13070_, _12700_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_13071_, _13070_, _05141_);
  and (_10936_, _13071_, _13069_);
  nor (_10940_, _12498_, rst);
  and (_13072_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_13073_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or (_13074_, _13073_, _13072_);
  and (_10943_, _13074_, _05141_);
  nor (_10986_, _12550_, rst);
  nand (_13075_, _11418_, _07434_);
  or (_13076_, _11418_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_13077_, _13076_, _05141_);
  and (_11030_, _13077_, _13075_);
  and (_13078_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_13079_, _12091_, _12050_);
  nor (_13080_, _13079_, _12092_);
  or (_13081_, _13080_, _07135_);
  or (_13082_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_13083_, _13082_, _12108_);
  and (_13084_, _13083_, _13081_);
  or (_11034_, _13084_, _13078_);
  and (_13085_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_13086_, _12094_, _12038_);
  nor (_13087_, _13086_, _12095_);
  or (_13088_, _13087_, _07135_);
  or (_13089_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_13090_, _13089_, _12108_);
  and (_13091_, _13090_, _13088_);
  or (_11063_, _13091_, _13085_);
  nor (_13092_, _12093_, _12042_);
  nor (_13093_, _13092_, _12094_);
  or (_13094_, _13093_, _07135_);
  or (_13095_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_13096_, _13095_, _12108_);
  and (_13097_, _13096_, _13094_);
  and (_13098_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_11068_, _13098_, _13097_);
  and (_13099_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_13100_, _12092_, _12046_);
  nor (_13101_, _13100_, _12093_);
  or (_13102_, _13101_, _07135_);
  or (_13103_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_13104_, _13103_, _12108_);
  and (_13105_, _13104_, _13102_);
  or (_11077_, _13105_, _13099_);
  or (_13106_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_13107_, _07619_, _06353_);
  and (_13108_, _13107_, _05141_);
  and (_11094_, _13108_, _13106_);
  and (_13109_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_13110_, _07619_, _06379_);
  or (_13111_, _13110_, _13109_);
  and (_11098_, _13111_, _05141_);
  and (_13112_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_13113_, _07619_, _06459_);
  or (_13114_, _13113_, _13112_);
  and (_11100_, _13114_, _05141_);
  and (_13115_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_13116_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_13117_, pc_log_change, _13116_);
  or (_13118_, _13117_, _13115_);
  and (_11104_, _13118_, _05141_);
  and (_13119_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_13120_, _07619_, _06376_);
  or (_13121_, _13120_, _13119_);
  and (_11107_, _13121_, _05141_);
  or (_13122_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_13123_, _07619_, _06306_);
  and (_13124_, _13123_, _05141_);
  and (_11161_, _13124_, _13122_);
  or (_13125_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_13126_, _07619_, _06516_);
  and (_13127_, _13126_, _05141_);
  and (_11163_, _13127_, _13125_);
  or (_13128_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_13129_, _07619_, _06484_);
  and (_13130_, _13129_, _05141_);
  and (_11166_, _13130_, _13128_);
  or (_13131_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not (_13132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_13133_, _06728_, _13132_);
  and (_13134_, _13133_, _13131_);
  or (_13135_, _13134_, _06738_);
  nand (_13136_, _06738_, _05604_);
  and (_13137_, _13136_, _13135_);
  or (_13138_, _13137_, _06743_);
  nand (_13139_, _06743_, _08441_);
  and (_13140_, _13139_, _05141_);
  and (_11180_, _13140_, _13138_);
  or (_13141_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_13142_, _07619_, _06311_);
  and (_13143_, _13142_, _05141_);
  and (_11214_, _13143_, _13141_);
  and (_13144_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_13145_, _07619_, _06399_);
  or (_13146_, _13145_, _13144_);
  and (_11217_, _13146_, _05141_);
  and (_13147_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_13148_, _07619_, _06403_);
  or (_13149_, _13148_, _13147_);
  and (_11221_, _13149_, _05141_);
  and (_11229_, _11737_, _05141_);
  or (_13150_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_13151_, _07619_, _06374_);
  and (_13152_, _13151_, _05141_);
  and (_11236_, _13152_, _13150_);
  or (_13153_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not (_13154_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_13155_, pc_log_change, _13154_);
  and (_13156_, _13155_, _05141_);
  and (_11239_, _13156_, _13153_);
  and (_13157_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_13158_, _13157_, _11815_);
  not (_13159_, _08439_);
  nor (_13160_, _11811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_13161_, _13160_, _11812_);
  or (_13162_, _13161_, _13159_);
  or (_13163_, _13162_, _13158_);
  or (_13164_, _08439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_13165_, _13164_, _13163_);
  or (_13166_, _13165_, _08463_);
  nor (_13167_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_13168_, _13167_, _08471_);
  and (_13169_, _13168_, _13166_);
  and (_13170_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_13171_, _13170_, _08478_);
  or (_13172_, _13171_, _13169_);
  or (_13173_, _11789_, _05522_);
  and (_13175_, _13173_, _05141_);
  and (_11254_, _13175_, _13172_);
  or (_13176_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_13177_, _07619_, _06370_);
  and (_13178_, _13177_, _05141_);
  and (_11259_, _13178_, _13176_);
  and (_13179_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_13180_, _07619_, _06427_);
  or (_13181_, _13180_, _13179_);
  and (_11263_, _13181_, _05141_);
  or (_13182_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand (_13183_, _07619_, _06510_);
  and (_13184_, _13183_, _05141_);
  and (_11281_, _13184_, _13182_);
  nand (_13185_, _11418_, _06617_);
  or (_13186_, _11418_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_13187_, _13186_, _05141_);
  and (_11300_, _13187_, _13185_);
  or (_13188_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_13189_, _07619_, _06406_);
  and (_13190_, _13189_, _05141_);
  and (_11310_, _13190_, _13188_);
  and (_13191_, _07611_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_13192_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_13193_, _13192_, _13191_);
  and (_11319_, _13193_, _05141_);
  and (_13194_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _07611_);
  and (_13195_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_13196_, _13195_, _13194_);
  and (_11323_, _13196_, _05141_);
  and (_13197_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07611_);
  and (_13198_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_13199_, _13198_, _13197_);
  and (_11335_, _13199_, _05141_);
  and (_13200_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07611_);
  and (_13201_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_13202_, _13201_, _13200_);
  and (_11346_, _13202_, _05141_);
  or (_13203_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand (_13204_, _07619_, _06429_);
  and (_13206_, _13204_, _05141_);
  and (_11356_, _13206_, _13203_);
  and (_13208_, _06290_, _05617_);
  and (_13209_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or (_13210_, _13209_, _13208_);
  and (_11360_, _13210_, _05141_);
  or (_13211_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_13212_, _07619_, _06395_);
  and (_13213_, _13212_, _05141_);
  and (_11363_, _13213_, _13211_);
  or (_13214_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_13215_, _07619_, _06489_);
  and (_13216_, _13215_, _05141_);
  and (_11376_, _13216_, _13214_);
  or (_13217_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand (_13218_, _07619_, _06438_);
  and (_13219_, _13218_, _05141_);
  and (_11389_, _13219_, _13217_);
  or (_13220_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_13221_, _07619_, _06343_);
  and (_13222_, _13221_, _05141_);
  and (_11409_, _13222_, _13220_);
  or (_13223_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand (_13224_, _07619_, _06464_);
  and (_13225_, _13224_, _05141_);
  and (_11416_, _13225_, _13223_);
  and (_11515_, _11745_, _05141_);
  nor (_11523_, _11742_, rst);
  nand (_13226_, _08305_, _05560_);
  or (_13227_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_13228_, _13227_, _05141_);
  and (_11526_, _13228_, _13226_);
  nor (_13229_, _11619_, _11617_);
  nor (_13230_, _13229_, _11620_);
  or (_13231_, _13230_, _07516_);
  or (_13232_, _06271_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_13233_, _13232_, _12108_);
  and (_11616_, _13233_, _13231_);
  and (_13234_, _11615_, _06271_);
  nand (_13235_, _13234_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_13236_, _13234_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_13237_, _13236_, _12108_);
  and (_11632_, _13237_, _13235_);
  or (_13238_, _11477_, _07011_);
  and (_13239_, _06524_, _06497_);
  and (_13240_, _13239_, _07014_);
  or (_13241_, _13240_, _11501_);
  and (_13242_, _13241_, _13238_);
  not (_13243_, _11546_);
  or (_13244_, _13243_, _07029_);
  or (_13245_, _13244_, _13242_);
  and (_13246_, _11511_, _07012_);
  nor (_13247_, _11596_, _11478_);
  or (_13248_, _13247_, _07013_);
  or (_13249_, _13248_, _13246_);
  and (_13250_, _11477_, _11549_);
  and (_13251_, _11543_, _07009_);
  or (_13252_, _11609_, _13251_);
  or (_13253_, _13252_, _13250_);
  or (_13254_, _11504_, _11585_);
  or (_13255_, _11564_, _11548_);
  or (_13256_, _13255_, _13254_);
  or (_13257_, _13256_, _13253_);
  or (_13258_, _13257_, _13249_);
  or (_13259_, _13258_, _13245_);
  and (_13261_, _13259_, _06272_);
  nor (_13262_, _07005_, _06790_);
  or (_13263_, _13262_, rst);
  or (_11638_, _13263_, _13261_);
  and (_13264_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_13265_, _07619_, _06301_);
  or (_13266_, _13265_, _13264_);
  and (_11641_, _13266_, _05141_);
  and (_13267_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_13268_, _07619_, _06351_);
  or (_13269_, _13268_, _13267_);
  and (_11645_, _13269_, _05141_);
  nand (_13270_, _06832_, _06449_);
  and (_13271_, _13270_, _06830_);
  or (_13272_, _06541_, _06831_);
  or (_11658_, _13272_, _13271_);
  and (_13273_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_13274_, _07619_, _06514_);
  or (_13275_, _13274_, _13273_);
  and (_11664_, _13275_, _05141_);
  and (_13276_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_13277_, _07619_, _06487_);
  or (_13278_, _13277_, _13276_);
  and (_11666_, _13278_, _05141_);
  and (_13279_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_13280_, _07619_, _06324_);
  or (_13281_, _13280_, _13279_);
  and (_11670_, _13281_, _05141_);
  and (_13282_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_13283_, _07619_, _06347_);
  or (_13284_, _13283_, _13282_);
  and (_11675_, _13284_, _05141_);
  nand (_13285_, _06472_, _06270_);
  or (_13286_, _06270_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_13287_, _13286_, _05141_);
  and (_11677_, _13287_, _13285_);
  and (_13288_, _06755_, _06547_);
  or (_13289_, _13288_, _07060_);
  or (_13290_, _13289_, _06785_);
  and (_13291_, _13290_, _06296_);
  and (_13292_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_13293_, _13292_, _06798_);
  and (_13294_, _13293_, _05141_);
  or (_11679_, _13294_, _13291_);
  and (_13295_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_13296_, _07619_, _06482_);
  or (_13297_, _13296_, _13295_);
  and (_11682_, _13297_, _05141_);
  or (_13298_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand (_13299_, _07619_, _06434_);
  and (_13300_, _13299_, _05141_);
  and (_11688_, _13300_, _13298_);
  and (_13301_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_13302_, _07619_, _06457_);
  or (_13303_, _13302_, _13301_);
  and (_11695_, _13303_, _05141_);
  and (_11697_, _11454_, _05141_);
  nand (_13304_, _08305_, _06178_);
  or (_13305_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_13306_, _13305_, _05141_);
  and (_11700_, _13306_, _13304_);
  and (_13307_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_13308_, _07619_, _06508_);
  or (_13309_, _13308_, _13307_);
  and (_11703_, _13309_, _05141_);
  or (_13310_, _08306_, _05522_);
  or (_13311_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_13312_, _13311_, _05141_);
  and (_11717_, _13312_, _13310_);
  and (_11719_, _12158_, _05141_);
  nand (_13313_, _06707_, _06062_);
  or (_13314_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_13315_, _13314_, _05141_);
  and (_11890_, _13315_, _13313_);
  nand (_13316_, _11418_, _07496_);
  or (_13317_, _11418_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_13318_, _13317_, _05141_);
  and (_11921_, _13318_, _13316_);
  nand (_13319_, _11418_, _07350_);
  or (_13320_, _11418_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_13321_, _13320_, _05141_);
  and (_11947_, _13321_, _13319_);
  and (_13322_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_13323_, _13322_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_11968_, _13323_, _05141_);
  and (_13324_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_13325_, _13324_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_11975_, _13325_, _05141_);
  or (_13326_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand (_13327_, _07619_, _06351_);
  and (_13328_, _13327_, _05141_);
  and (_11979_, _13328_, _13326_);
  or (_13329_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand (_13330_, _07619_, _06482_);
  and (_13331_, _13330_, _05141_);
  and (_11987_, _13331_, _13329_);
  and (_13333_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_13334_, _13333_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_11993_, _13334_, _05141_);
  or (_13335_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand (_13336_, _07619_, _06459_);
  and (_13337_, _13336_, _05141_);
  and (_11995_, _13337_, _13335_);
  and (_13338_, _05287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_13339_, _13338_, _10356_);
  and (_13340_, _13339_, _11458_);
  nand (_13341_, _11458_, _08283_);
  and (_13342_, _13341_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_13343_, _13342_, _11462_);
  or (_13344_, _13343_, _13340_);
  nand (_13345_, _11462_, _05560_);
  and (_13346_, _13345_, _05141_);
  and (_12002_, _13346_, _13344_);
  and (_13347_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_13348_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or (_13349_, _13348_, _13347_);
  and (_12008_, _13349_, _05141_);
  and (_13350_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _05141_);
  and (_13351_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _05141_);
  and (_13353_, _13351_, _11643_);
  or (_12013_, _13353_, _13350_);
  and (_13354_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_13355_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or (_13356_, _13355_, _13354_);
  and (_12016_, _13356_, _05141_);
  and (_13357_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_13358_, _13357_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_12018_, _13358_, _05141_);
  or (_13359_, _06745_, _06004_);
  and (_13360_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_13361_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_13362_, _13361_, _13360_);
  or (_13363_, _13362_, _06743_);
  and (_13364_, _13363_, _05141_);
  and (_12058_, _13364_, _13359_);
  and (_13365_, _06742_, _05649_);
  not (_13366_, _13365_);
  or (_13368_, _13366_, _06004_);
  not (_13369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_13370_, _13369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_13371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_13372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _13371_);
  nor (_13373_, _13372_, _13370_);
  not (_13374_, _13373_);
  nand (_13375_, _08476_, _05649_);
  and (_13376_, _13375_, _13374_);
  not (_13377_, _13376_);
  and (_13378_, _13377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  not (_13379_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_13381_, _13379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  not (_13382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_13383_, \oc8051_top_1.oc8051_sfr1.pres_ow , _13382_);
  not (_13384_, t1_i);
  and (_13385_, _13384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_13386_, _13385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or (_13388_, _13386_, _13383_);
  and (_13389_, _13388_, _13381_);
  and (_13391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_13392_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_13393_, _13392_, _13391_);
  and (_13394_, _13393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_13395_, _13394_, _13389_);
  nor (_13396_, _13395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_13397_, _13395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_13398_, _13397_, _13396_);
  and (_13399_, _13374_, _13398_);
  and (_13400_, _13397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_13401_, _13400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_13402_, _13401_, _13370_);
  and (_13403_, _13402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_13404_, _13403_, _13399_);
  and (_13405_, _13404_, _13375_);
  or (_13406_, _13405_, _13378_);
  or (_13407_, _13365_, _13406_);
  and (_13408_, _13407_, _05141_);
  and (_12067_, _13408_, _13368_);
  and (_13409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_13410_, _13409_);
  and (_13412_, _13410_, _13375_);
  and (_13413_, _13393_, _13389_);
  and (_13414_, _13413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_13415_, _13413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_13416_, _13415_, _13414_);
  and (_13417_, _13416_, _13412_);
  not (_13418_, _13412_);
  and (_13419_, _13418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or (_13420_, _13419_, _13417_);
  and (_13421_, _13402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_13422_, _13421_, _13375_);
  or (_13423_, _13422_, _13365_);
  or (_13424_, _13423_, _13420_);
  or (_13425_, _13366_, _05522_);
  and (_13426_, _13425_, _05141_);
  and (_12070_, _13426_, _13424_);
  and (_13427_, _13389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_13428_, _13427_, _13391_);
  nor (_13429_, _13428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_13430_, _13429_, _13413_);
  nand (_13432_, _13430_, _13412_);
  or (_13433_, _13412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_13434_, _13433_, _13432_);
  and (_13435_, _05649_, _05173_);
  and (_13437_, _13435_, _06032_);
  and (_13438_, _13437_, _05925_);
  and (_13439_, _05965_, _05925_);
  and (_13440_, _13414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_13441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_13442_, _13441_, _13440_);
  and (_13443_, _13442_, _13370_);
  nand (_13444_, _13443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_13445_, _13444_, _13439_);
  or (_13446_, _13445_, _13438_);
  or (_13447_, _13446_, _13434_);
  nand (_13448_, _13438_, _06062_);
  and (_13449_, _13448_, _05141_);
  and (_12073_, _13449_, _13447_);
  nor (_12076_, _12287_, rst);
  nand (_13450_, _13365_, _06244_);
  nor (_13451_, _13397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_13452_, _13451_, _13400_);
  and (_13453_, _13452_, _13376_);
  and (_13454_, _13377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_13455_, _13443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_13456_, _13455_, _13439_);
  or (_13457_, _13456_, _13454_);
  or (_13458_, _13457_, _13453_);
  or (_13459_, _13458_, _13365_);
  and (_13460_, _13459_, _05141_);
  and (_12080_, _13460_, _13450_);
  nor (_12082_, _12425_, rst);
  nand (_13461_, _08305_, _06062_);
  or (_13462_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_13463_, _13462_, _05141_);
  and (_12085_, _13463_, _13461_);
  not (_13464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_13465_, _13412_, _13464_);
  or (_13466_, _13389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_13467_, _13427_, _13409_);
  and (_13468_, _13467_, _13466_);
  and (_13469_, _13370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_13470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_13471_, _13470_, _13441_);
  and (_13472_, _13471_, _13393_);
  and (_13473_, _13472_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_13474_, _13473_, _13469_);
  or (_00003_, _13474_, _13468_);
  and (_00004_, _00003_, _13375_);
  or (_00005_, _00004_, _13365_);
  or (_00006_, _00005_, _13465_);
  nand (_00007_, _13365_, _05604_);
  and (_00008_, _00007_, _05141_);
  and (_12090_, _00008_, _00006_);
  and (_00009_, _13427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_00010_, _13427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_00011_, _00010_, _00009_);
  and (_00012_, _00011_, _13412_);
  nand (_00013_, _13443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_00014_, _00013_, _13439_);
  or (_00015_, _00014_, _00012_);
  and (_00016_, _13418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_00017_, _00016_, _13365_);
  or (_00018_, _00017_, _00015_);
  nand (_00019_, _13365_, _06178_);
  and (_00020_, _00019_, _05141_);
  and (_12098_, _00020_, _00018_);
  nor (_00021_, _00009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_00022_, _00021_, _13428_);
  and (_00023_, _00022_, _13412_);
  and (_00024_, _13418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_00025_, _00024_, _00023_);
  and (_00026_, _13402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00027_, _00026_, _13375_);
  or (_00028_, _00027_, _13365_);
  or (_00029_, _00028_, _00025_);
  nand (_00030_, _13365_, _05560_);
  and (_00031_, _00030_, _05141_);
  and (_12102_, _00031_, _00029_);
  nor (_12104_, _12186_, rst);
  nor (_12109_, _12796_, rst);
  nor (_12113_, _12368_, rst);
  nor (_12116_, _12604_, rst);
  or (_00032_, _13375_, _06179_);
  not (_00033_, _13372_);
  and (_00034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00035_, _13441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_00036_, _00035_, _00034_);
  and (_00037_, _00036_, _13393_);
  and (_00038_, _00037_, _13389_);
  nor (_00039_, _00038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00040_, _13473_, _13389_);
  and (_00041_, _00040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_00042_, _00041_, _00039_);
  or (_00043_, _00042_, _00033_);
  and (_00044_, _00034_, _13393_);
  and (_00045_, _00044_, _13389_);
  nor (_00046_, _00045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_00047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_00048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_00050_, _00049_, _13414_);
  nand (_00051_, _00050_, _00048_);
  and (_00052_, _00051_, _00047_);
  or (_00053_, _00052_, _00046_);
  and (_00054_, _00053_, _00043_);
  nand (_00055_, _00054_, _13375_);
  and (_00056_, _00055_, _13366_);
  and (_00057_, _00056_, _00032_);
  and (_00058_, _13438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_00059_, _00058_, _00057_);
  and (_12119_, _00059_, _05141_);
  not (_00060_, _13438_);
  and (_00061_, _13439_, _05560_);
  or (_00062_, _00041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00064_, _00063_, _00040_);
  nor (_00065_, _00064_, _00033_);
  nand (_00066_, _00065_, _00062_);
  nor (_00067_, _00050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_00068_, _00067_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00069_, _00034_, _13413_);
  and (_00070_, _00063_, _13371_);
  and (_00071_, _00070_, _00069_);
  nor (_00072_, _00071_, _13372_);
  nand (_00073_, _00072_, _00068_);
  and (_00074_, _00073_, _00066_);
  and (_00075_, _00074_, _13375_);
  or (_00076_, _00075_, _00061_);
  nand (_00077_, _00076_, _00060_);
  or (_00078_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00079_, _00078_, _05141_);
  and (_12122_, _00079_, _00077_);
  not (_00080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00081_, _00048_, _13414_);
  and (_00082_, _13442_, _13372_);
  nor (_00083_, _00082_, _00081_);
  nand (_00084_, _00083_, _00080_);
  or (_00085_, _00083_, _00080_);
  nand (_00086_, _00085_, _00084_);
  nor (_00087_, _00086_, _13439_);
  and (_00088_, _13439_, _06703_);
  or (_00089_, _00088_, _00087_);
  or (_00090_, _00089_, _13365_);
  nand (_00091_, _13365_, _00080_);
  and (_00092_, _00091_, _05141_);
  and (_12125_, _00092_, _00090_);
  and (_00093_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_00094_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_00095_, _00094_, _00093_);
  or (_00096_, _00095_, _06743_);
  nand (_00097_, _06743_, _05560_);
  and (_00098_, _00097_, _05141_);
  and (_12128_, _00098_, _00096_);
  or (_00099_, _13375_, _05522_);
  nand (_00100_, _00071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00101_, _00100_, _00033_);
  and (_00102_, _00063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00103_, _00102_, _00038_);
  nor (_00104_, _00103_, _00033_);
  nor (_00105_, _00104_, _00101_);
  or (_00106_, _00105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_00107_, _00105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_00108_, _00107_, _00106_);
  and (_00109_, _00108_, _13375_);
  nor (_00110_, _00109_, _13365_);
  and (_00111_, _00110_, _00099_);
  and (_00112_, _06034_, _05925_);
  and (_00113_, _00112_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_00114_, _00113_, _00111_);
  and (_12134_, _00114_, _05141_);
  and (_00115_, _13439_, _06244_);
  not (_00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_00117_, _00107_, _00116_);
  and (_00118_, _00117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00119_, _00117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_00120_, _00119_, _00118_);
  nor (_00121_, _00120_, _13439_);
  or (_00122_, _00121_, _00115_);
  nand (_00123_, _00122_, _00060_);
  or (_00124_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_00125_, _00124_, _05141_);
  and (_12137_, _00125_, _00123_);
  or (_00126_, _13375_, _06004_);
  nand (_00127_, _00107_, _00116_);
  and (_00128_, _00127_, _00117_);
  nor (_00129_, _00128_, _13439_);
  nor (_00130_, _00129_, _13365_);
  and (_00131_, _00130_, _00126_);
  and (_00132_, _00112_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_00133_, _00132_, _00131_);
  and (_12140_, _00133_, _05141_);
  and (_00134_, _13439_, _06062_);
  nor (_00135_, _00072_, _00065_);
  not (_00136_, _00135_);
  nand (_00137_, _00136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_00138_, _00136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00139_, _00138_, _00137_);
  and (_00140_, _00139_, _13375_);
  or (_00141_, _00140_, _00134_);
  nand (_00142_, _00141_, _00060_);
  or (_00143_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00144_, _00143_, _05141_);
  and (_12143_, _00144_, _00142_);
  or (_00145_, _12912_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00146_, _00145_, _12913_);
  or (_00148_, _00146_, _12773_);
  nand (_00149_, _12904_, _05455_);
  and (_00150_, _00149_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_00151_, _00150_, _12969_);
  and (_00152_, _00151_, _12973_);
  and (_00153_, _00152_, _00148_);
  and (_00154_, _12701_, _07319_);
  and (_00155_, _12707_, _12843_);
  nor (_00156_, _12703_, _07350_);
  or (_00157_, _00156_, _00155_);
  or (_00159_, _12985_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00160_, _00159_, _12724_);
  and (_00161_, _00160_, _12713_);
  and (_00162_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_00163_, _00162_, _00161_);
  or (_00164_, _00163_, _00157_);
  nor (_00165_, _00164_, _00154_);
  nand (_00166_, _00165_, _12700_);
  or (_00167_, _00166_, _00153_);
  nor (_00168_, _13002_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00169_, _00168_, _13003_);
  or (_00170_, _00169_, _12700_);
  and (_00171_, _00170_, _05141_);
  and (_12146_, _00171_, _00167_);
  not (_00173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_00174_, t0_i);
  and (_00175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _00174_);
  nor (_00176_, _00175_, _00173_);
  not (_00177_, _00176_);
  not (_00178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_00179_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_00180_, _00179_, _00178_);
  and (_00181_, _00180_, _00177_);
  and (_00182_, _00181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_00183_, _00182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_00184_, _00182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_00185_, _00184_, _00183_);
  not (_00186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _00186_);
  and (_00188_, _00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00189_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_00190_, _00189_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_00191_, _00190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_00192_, _00191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_00193_, _00192_, _00181_);
  and (_00194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00195_, _00194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_00196_, _00195_, _00193_);
  and (_00197_, _00196_, _00188_);
  nor (_00198_, _00197_, _00185_);
  and (_00199_, _08470_, _05649_);
  nor (_00200_, _00199_, _00198_);
  and (_00201_, _00199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_00202_, _00201_, _00200_);
  and (_00203_, _06737_, _05649_);
  not (_00204_, _00203_);
  and (_00205_, _00204_, _00202_);
  nor (_00206_, _00204_, _06178_);
  or (_00207_, _00206_, _00205_);
  and (_12154_, _00207_, _05141_);
  not (_00208_, _12796_);
  and (_00210_, _00208_, _12707_);
  and (_00211_, _13058_, _06669_);
  and (_00212_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_00213_, _12713_, _12776_);
  or (_00214_, _00213_, _00212_);
  or (_00215_, _00214_, _00211_);
  and (_00216_, _12899_, _12896_);
  or (_00217_, _00216_, _12840_);
  or (_00218_, _00217_, _12806_);
  and (_00219_, _00217_, _12806_);
  not (_00220_, _00219_);
  and (_00221_, _00220_, _12940_);
  and (_00222_, _00221_, _00218_);
  or (_00223_, _00222_, _00215_);
  or (_00224_, _00223_, _00210_);
  and (_00225_, _00224_, _12700_);
  and (_00226_, _07622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_00227_, _00226_, _12943_);
  and (_00228_, _00226_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00229_, _00228_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00230_, _00229_, _00227_);
  nor (_00231_, _00230_, _12700_);
  or (_00232_, _00231_, _00225_);
  and (_12157_, _00232_, _05141_);
  not (_00233_, _00181_);
  nor (_00234_, _00199_, _00233_);
  or (_00235_, _00234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_00236_, _00195_, _00192_);
  and (_00237_, _00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_00238_, _00237_, _00236_);
  nand (_00239_, _00238_, _00182_);
  or (_00240_, _00239_, _00199_);
  and (_00241_, _00240_, _00235_);
  or (_00242_, _00241_, _00203_);
  nand (_00243_, _00203_, _05604_);
  and (_00244_, _00243_, _05141_);
  and (_12160_, _00244_, _00242_);
  or (_00245_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_00246_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_00247_, _00246_, _00245_);
  or (_00248_, _00247_, _06743_);
  nand (_00249_, _06743_, _06178_);
  and (_00250_, _00249_, _05141_);
  and (_12163_, _00250_, _00248_);
  and (_00251_, _00190_, _00181_);
  nor (_00252_, _00184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_00253_, _00252_, _00251_);
  and (_00254_, _00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00255_, _00254_, _00196_);
  nor (_00256_, _00255_, _00253_);
  nor (_00257_, _00256_, _00199_);
  and (_00258_, _00199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_00259_, _00258_, _00257_);
  and (_00260_, _00259_, _00204_);
  nor (_00261_, _00204_, _05560_);
  or (_00262_, _00261_, _00260_);
  and (_12180_, _00262_, _05141_);
  or (_00263_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_00264_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_00265_, _08417_, _00264_);
  and (_00266_, _00265_, _00263_);
  or (_00267_, _00266_, _06743_);
  nand (_00268_, _06743_, _05604_);
  and (_00269_, _00268_, _05141_);
  and (_12183_, _00269_, _00267_);
  and (_00270_, _00251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_00271_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_00272_, _00271_, _00193_);
  and (_00273_, _00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00274_, _00273_, _00196_);
  nor (_00275_, _00274_, _00272_);
  nor (_00276_, _00275_, _00199_);
  and (_00277_, _00199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_00278_, _00277_, _00276_);
  and (_00279_, _00278_, _00204_);
  and (_00280_, _00203_, _05522_);
  or (_00281_, _00280_, _00279_);
  and (_12187_, _00281_, _05141_);
  nor (_00282_, _00251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_00283_, _00282_, _00270_);
  and (_00284_, _00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00285_, _00284_, _00196_);
  nor (_00286_, _00285_, _00283_);
  nor (_00287_, _00286_, _00199_);
  and (_00288_, _00199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_00289_, _00288_, _00287_);
  and (_00290_, _00289_, _00204_);
  nor (_00291_, _00204_, _06062_);
  or (_00292_, _00291_, _00290_);
  and (_12190_, _00292_, _05141_);
  or (_00293_, _08345_, _06004_);
  and (_00294_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_00295_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_00296_, _00295_, _00294_);
  or (_00297_, _00296_, _06738_);
  and (_00298_, _00297_, _06745_);
  and (_00299_, _00298_, _00293_);
  and (_00300_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_00301_, _00300_, _00299_);
  and (_12198_, _00301_, _05141_);
  or (_00303_, _08345_, _05522_);
  and (_00304_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_00305_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_00306_, _00305_, _00304_);
  or (_00307_, _00306_, _06738_);
  and (_00308_, _00307_, _06745_);
  and (_00309_, _00308_, _00303_);
  and (_00310_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_00311_, _00310_, _00309_);
  and (_12203_, _00311_, _05141_);
  nand (_00312_, _06738_, _06062_);
  and (_00313_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_00314_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_00315_, _00314_, _00313_);
  or (_00316_, _00315_, _06738_);
  and (_00317_, _00316_, _06745_);
  and (_00318_, _00317_, _00312_);
  and (_00319_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_00320_, _00319_, _00318_);
  and (_12206_, _00320_, _05141_);
  nand (_00321_, _06738_, _05560_);
  and (_00322_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_00323_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_00324_, _00323_, _00322_);
  or (_00325_, _00324_, _06738_);
  and (_00326_, _00325_, _06745_);
  and (_00327_, _00326_, _00321_);
  and (_00328_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_00329_, _00328_, _00327_);
  and (_12210_, _00329_, _05141_);
  nor (_00330_, _12088_, _12060_);
  nor (_00331_, _00330_, _12089_);
  or (_00332_, _00331_, _07135_);
  or (_00333_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_00334_, _00333_, _12108_);
  and (_00335_, _00334_, _00332_);
  and (_00336_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_12212_, _00336_, _00335_);
  nor (_00337_, _12071_, _11615_);
  nor (_00338_, _00337_, _12072_);
  or (_00339_, _00338_, _07135_);
  or (_00340_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_00342_, _00340_, _12108_);
  and (_00344_, _00342_, _00339_);
  and (_00346_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_12218_, _00346_, _00344_);
  nor (_00347_, _12095_, _12034_);
  nor (_00348_, _00347_, _12096_);
  or (_00350_, _00348_, _07135_);
  or (_00351_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00352_, _00351_, _12108_);
  and (_00353_, _00352_, _00350_);
  and (_00354_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_12227_, _00354_, _00353_);
  nor (_00356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not (_00358_, _00356_);
  and (_00359_, _00358_, _00193_);
  and (_00360_, _00359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_00361_, _00360_);
  nor (_00362_, _00361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00363_, _00196_, _00187_);
  and (_00364_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_00365_, _00364_, _00362_);
  nor (_00367_, _00365_, _00199_);
  or (_00368_, _00361_, _00199_);
  and (_00369_, _00368_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_00371_, _00369_, _00367_);
  and (_00372_, _00371_, _00204_);
  nor (_00373_, _00204_, _06244_);
  or (_00375_, _00373_, _00372_);
  and (_12242_, _00375_, _05141_);
  not (_00378_, _00199_);
  or (_00380_, _00378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_00381_, _00380_, _00204_);
  and (_00382_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_00383_, _00359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_00384_, _00383_, _00368_);
  or (_00385_, _00384_, _00382_);
  and (_00386_, _00385_, _00381_);
  and (_00388_, _00203_, _06004_);
  or (_00389_, _00388_, _00386_);
  and (_12246_, _00389_, _05141_);
  nand (_00390_, _00199_, _06244_);
  not (_00391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00392_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00394_, _00393_, _00193_);
  and (_00395_, _00394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00396_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00397_, _00396_, _00392_);
  nor (_00398_, _00397_, _00391_);
  and (_00399_, _00397_, _00391_);
  or (_00400_, _00399_, _00398_);
  and (_00401_, _00400_, _00356_);
  and (_00402_, _00393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00403_, _00402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00404_, _00403_, _00392_);
  and (_00405_, _00236_, _00181_);
  and (_00406_, _00405_, _00404_);
  or (_00407_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_00408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00409_, _00408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00410_, _00404_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_00411_, _00410_, _00405_);
  and (_00412_, _00411_, _00409_);
  and (_00413_, _00412_, _00407_);
  and (_00414_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_00415_, _00414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00416_, _00415_, _00404_);
  nand (_00417_, _00416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_00418_, _00416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00419_, _00418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00420_, _00419_, _00417_);
  or (_00421_, _00420_, _00413_);
  or (_00422_, _00421_, _00401_);
  or (_00423_, _00422_, _00199_);
  and (_00424_, _00423_, _00204_);
  and (_00425_, _00424_, _00390_);
  and (_00426_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_00427_, _00426_, _00425_);
  and (_12284_, _00427_, _05141_);
  nand (_00428_, _00199_, _05560_);
  or (_00429_, _00394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_00430_, _00395_, _00358_);
  and (_00431_, _00430_, _00429_);
  and (_00432_, _00405_, _00393_);
  or (_00433_, _00432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_00434_, _00405_, _00402_);
  and (_00435_, _00434_, _00409_);
  and (_00436_, _00435_, _00433_);
  and (_00437_, _00414_, _00402_);
  nand (_00438_, _00437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00439_, _00414_, _00393_);
  and (_00440_, _00439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_00441_, _00440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00442_, _00441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00443_, _00442_, _00438_);
  or (_00444_, _00443_, _00436_);
  or (_00445_, _00444_, _00431_);
  or (_00446_, _00445_, _00199_);
  and (_00447_, _00446_, _00204_);
  and (_00448_, _00447_, _00428_);
  and (_00449_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_00450_, _00449_, _00448_);
  and (_12295_, _00450_, _05141_);
  nand (_00451_, _00199_, _06062_);
  and (_00452_, _00405_, _00408_);
  and (_00453_, _00452_, _00402_);
  nand (_00454_, _00453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_00455_, _00409_, _00187_);
  or (_00456_, _00453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00458_, _00456_, _00455_);
  and (_00459_, _00458_, _00454_);
  or (_00460_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_00461_, _00396_, _00358_);
  and (_00462_, _00461_, _00460_);
  or (_00463_, _00437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00465_, _00414_, _00403_);
  not (_00466_, _00465_);
  and (_00467_, _00466_, _00464_);
  and (_00468_, _00467_, _00463_);
  or (_00469_, _00468_, _00462_);
  or (_00470_, _00469_, _00459_);
  or (_00471_, _00470_, _00199_);
  and (_00472_, _00471_, _00204_);
  and (_00473_, _00472_, _00451_);
  and (_00474_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_00475_, _00474_, _00473_);
  and (_12298_, _00475_, _05141_);
  or (_00476_, _00378_, _05522_);
  and (_00477_, _00403_, _00193_);
  or (_00478_, _00477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00479_, _00477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_00480_, _00479_, _00358_);
  and (_00481_, _00480_, _00478_);
  and (_00482_, _00192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_00483_, _00482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00484_, _00483_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_00485_, _00403_, _00181_);
  and (_00487_, _00485_, _00484_);
  and (_00488_, _00487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00489_, _00487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_00490_, _00489_, _00409_);
  nor (_00491_, _00490_, _00488_);
  and (_00492_, _00415_, _00403_);
  nand (_00493_, _00492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00494_, _00492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00495_, _00494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00496_, _00495_, _00493_);
  or (_00497_, _00496_, _00491_);
  or (_00498_, _00497_, _00481_);
  or (_00499_, _00498_, _00199_);
  and (_00500_, _00499_, _00204_);
  and (_00501_, _00500_, _00476_);
  and (_00502_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00503_, _00502_, _00501_);
  and (_12307_, _00503_, _05141_);
  or (_00504_, _00378_, _06004_);
  and (_00505_, _00488_, _00408_);
  nor (_00506_, _00505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00507_, _00505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_00508_, _00507_, _00506_);
  and (_00509_, _00508_, _00455_);
  and (_00510_, _00465_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_00511_, _00510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_00512_, _00510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00513_, _00512_, _00511_);
  and (_00514_, _00513_, _00464_);
  or (_00515_, _00479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_00516_, _00397_, _00358_);
  and (_00517_, _00516_, _00515_);
  or (_00518_, _00517_, _00514_);
  or (_00519_, _00518_, _00509_);
  or (_00520_, _00519_, _00199_);
  and (_00521_, _00520_, _00204_);
  and (_00522_, _00521_, _00504_);
  and (_00523_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_00524_, _00523_, _00522_);
  and (_12311_, _00524_, _05141_);
  nand (_00525_, _00199_, _06178_);
  and (_00526_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00527_, _00526_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_00528_, _00432_);
  and (_00529_, _00528_, _00409_);
  or (_00530_, _00529_, _00187_);
  and (_00531_, _00530_, _00527_);
  and (_00532_, _00414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00533_, _00532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_00534_, _00533_, _00464_);
  nor (_00535_, _00534_, _00439_);
  and (_00536_, _00193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00537_, _00536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_00538_, _00394_, _00358_);
  and (_00539_, _00538_, _00537_);
  or (_00540_, _00539_, _00535_);
  or (_00541_, _00540_, _00531_);
  or (_00542_, _00541_, _00199_);
  and (_00543_, _00542_, _00525_);
  or (_00544_, _00543_, _00203_);
  or (_00545_, _00204_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00546_, _00545_, _05141_);
  and (_12324_, _00546_, _00544_);
  or (_00547_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not (_00548_, _00526_);
  and (_00549_, _00548_, _00455_);
  and (_00550_, _00549_, _00547_);
  nor (_00551_, _00414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_00552_, _00551_, _00532_);
  and (_00553_, _00552_, _00464_);
  or (_00554_, _00193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_00555_, _00536_, _00358_);
  and (_00556_, _00555_, _00554_);
  or (_00557_, _00556_, _00553_);
  or (_00558_, _00557_, _00550_);
  or (_00559_, _00558_, _00199_);
  nand (_00560_, _00199_, _05604_);
  and (_00561_, _00560_, _00559_);
  or (_00562_, _00561_, _00203_);
  not (_00563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_00564_, _00203_, _00563_);
  and (_00565_, _00564_, _05141_);
  and (_12328_, _00565_, _00562_);
  and (_00566_, _08242_, _05649_);
  nand (_00567_, _00566_, _05604_);
  or (_00568_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00569_, _00568_, _05141_);
  and (_12334_, _00569_, _00567_);
  nand (_00570_, _00566_, _06178_);
  or (_00571_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00572_, _00571_, _05141_);
  and (_12337_, _00572_, _00570_);
  or (_00573_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_00574_, _00573_, _05141_);
  and (_00575_, _06184_, _05925_);
  nand (_00576_, _00575_, _06062_);
  and (_12342_, _00576_, _00574_);
  or (_00577_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_00578_, _00577_, _05141_);
  not (_00579_, _00575_);
  or (_00580_, _00579_, _05522_);
  and (_12345_, _00580_, _00578_);
  nand (_00581_, _00566_, _05560_);
  or (_00582_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_00583_, _00582_, _05141_);
  and (_12348_, _00583_, _00581_);
  or (_00584_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00585_, _00584_, _05141_);
  nand (_00586_, _00575_, _06244_);
  and (_12353_, _00586_, _00585_);
  or (_00587_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00588_, _00587_, _05141_);
  or (_00589_, _00579_, _06004_);
  and (_12360_, _00589_, _00588_);
  nand (_00590_, _08305_, _06244_);
  or (_00591_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_00592_, _00591_, _05141_);
  and (_12406_, _00592_, _00590_);
  and (_00593_, _05614_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_00594_, _06179_, _05617_);
  nand (_00595_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_00596_, _00595_, _05609_);
  or (_00597_, _00596_, _00594_);
  or (_00598_, _00597_, _00593_);
  and (_12536_, _00598_, _05141_);
  not (_00599_, _05576_);
  nor (_00600_, _05960_, _00599_);
  and (_00601_, _00599_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_00602_, _00601_, _05572_);
  or (_00603_, _00602_, _00600_);
  or (_00604_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_00605_, _00604_, _05141_);
  and (_12620_, _00605_, _00603_);
  or (_00606_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand (_00607_, _07619_, _06427_);
  and (_00608_, _00607_, _05141_);
  and (_12623_, _00608_, _00606_);
  nor (_00609_, _12628_, _06791_);
  not (_00610_, _12115_);
  or (_00611_, _12118_, _12130_);
  or (_00612_, _00611_, _00610_);
  and (_00613_, _07051_, _12627_);
  nand (_00614_, _00613_, _07034_);
  or (_00615_, _00614_, _12129_);
  or (_00616_, _00615_, _00612_);
  and (_00617_, _00616_, _06821_);
  or (_00618_, _00617_, _00609_);
  and (_12630_, _00618_, _05141_);
  and (_00619_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _07611_);
  and (_00620_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00621_, _00620_, _00619_);
  and (_12648_, _00621_, _05141_);
  nor (_12656_, _12827_, rst);
  and (_00622_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07611_);
  and (_00623_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00624_, _00623_, _00622_);
  and (_12661_, _00624_, _05141_);
  not (_00625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_00626_, _06683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_00627_, _00626_, _00625_);
  and (_00628_, _00627_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_00629_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_00630_, _00627_, _00629_);
  or (_00631_, _00630_, _00628_);
  or (_00632_, _00631_, _08280_);
  or (_00633_, _06620_, _00629_);
  nand (_00634_, _00633_, _08280_);
  or (_00635_, _00634_, _10356_);
  and (_00636_, _00635_, _00632_);
  or (_00637_, _00636_, _08289_);
  nand (_00638_, _08289_, _05560_);
  and (_00639_, _00638_, _05141_);
  and (_12722_, _00639_, _00637_);
  and (_00640_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _05141_);
  and (_00641_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _05141_);
  and (_00642_, _00641_, _11644_);
  or (_12734_, _00642_, _00640_);
  and (_00643_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_00644_, _00643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_12738_, _00644_, _05141_);
  and (_00645_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _07611_);
  and (_00646_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00647_, _00646_, _00645_);
  and (_12767_, _00647_, _05141_);
  and (_12788_, _12409_, _05141_);
  nor (_12791_, _12876_, rst);
  or (_00648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_00649_, _00648_, _08280_);
  not (_00650_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_00651_, _05288_, _00650_);
  nand (_00652_, _00651_, _08280_);
  or (_00653_, _00652_, _08178_);
  and (_00654_, _00653_, _00649_);
  or (_00655_, _00654_, _08289_);
  nand (_00656_, _08289_, _06178_);
  and (_00658_, _00656_, _05141_);
  and (_12815_, _00658_, _00655_);
  and (_12854_, _12257_, _05141_);
  and (_12856_, _12325_, _05141_);
  nand (_12858_, _12569_, _05141_);
  nand (_12861_, _12515_, _05141_);
  and (_00659_, _08280_, _10407_);
  and (_00661_, _00659_, _05963_);
  nor (_00662_, _00659_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_00663_, _00662_, _00661_);
  nand (_00664_, _00663_, _08360_);
  or (_00665_, _08360_, _06004_);
  and (_00667_, _00665_, _05141_);
  and (_12925_, _00667_, _00664_);
  or (_00668_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  not (_00669_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_00671_, pc_log_change, _00669_);
  and (_00672_, _00671_, _05141_);
  and (_13021_, _00672_, _00668_);
  and (_00673_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_00674_, pc_log_change, _00669_);
  or (_00675_, _00674_, _00673_);
  and (_13030_, _00675_, _05141_);
  and (_00676_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_00677_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_00678_, pc_log_change, _00677_);
  or (_00679_, _00678_, _00676_);
  and (_13067_, _00679_, _05141_);
  nand (_00680_, _06707_, _05560_);
  or (_00681_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_00682_, _00681_, _05141_);
  and (_13174_, _00682_, _00680_);
  and (_13205_, _12390_, _05141_);
  and (_13207_, _10319_, _12164_);
  and (_00683_, _05299_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_00685_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_00686_, _00685_, _05303_);
  and (_00687_, _05605_, _05284_);
  or (_00688_, _00687_, _00686_);
  or (_00689_, _00688_, _00683_);
  and (_13260_, _00689_, _05141_);
  and (_00690_, _10342_, _06879_);
  and (_00691_, _00690_, _06207_);
  nand (_00692_, _00691_, _05963_);
  or (_00693_, _00691_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_00694_, _00693_, _05647_);
  and (_00695_, _00694_, _00692_);
  not (_00696_, _05646_);
  and (_00697_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_00698_, _00690_, _05210_);
  not (_00699_, _00698_);
  or (_00700_, _00699_, _06669_);
  or (_00701_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_00702_, _00701_, _05925_);
  and (_00703_, _00702_, _00700_);
  or (_00704_, _00703_, _00697_);
  or (_00705_, _00704_, _00695_);
  and (_13332_, _00705_, _05141_);
  and (_00707_, _00690_, _05288_);
  nand (_00708_, _00707_, _05963_);
  or (_00709_, _00707_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_00710_, _00709_, _05647_);
  and (_00711_, _00710_, _00708_);
  and (_00712_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_00713_, _00699_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_00714_, _00699_, _07434_);
  or (_00715_, _00714_, _00713_);
  and (_00716_, _00715_, _05925_);
  or (_00717_, _00716_, _00712_);
  or (_00718_, _00717_, _00711_);
  and (_13352_, _00718_, _05141_);
  or (_00719_, _00699_, _05922_);
  or (_00720_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_00721_, _00720_, _05647_);
  and (_00722_, _00721_, _00719_);
  and (_00723_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_00724_, _00698_, _07496_);
  and (_00725_, _00720_, _05925_);
  and (_00726_, _00725_, _00724_);
  or (_00727_, _00726_, _00723_);
  or (_00728_, _00727_, _00722_);
  and (_13367_, _00728_, _05141_);
  not (_00729_, _00690_);
  or (_00730_, _00729_, _10375_);
  and (_00731_, _00730_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_00732_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_00733_, _00732_, _10380_);
  and (_00734_, _00733_, _00690_);
  or (_00735_, _00734_, _00731_);
  and (_00736_, _00735_, _05647_);
  not (_00737_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_00738_, _05646_, _00737_);
  nand (_00739_, _00698_, _07259_);
  or (_00740_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_00741_, _00740_, _05925_);
  and (_00742_, _00741_, _00739_);
  or (_00743_, _00742_, _00738_);
  or (_00744_, _00743_, _00736_);
  and (_13380_, _00744_, _05141_);
  nand (_00745_, _00690_, _05186_);
  and (_00746_, _00745_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not (_00747_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_00748_, _08282_, _00747_);
  or (_00749_, _00748_, _08281_);
  and (_00750_, _00749_, _00690_);
  or (_00751_, _00750_, _00746_);
  and (_00752_, _00751_, _05647_);
  nor (_00753_, _05646_, _00747_);
  nand (_00754_, _00698_, _07350_);
  or (_00755_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_00756_, _00755_, _05925_);
  and (_00757_, _00756_, _00754_);
  or (_00758_, _00757_, _00753_);
  or (_00759_, _00758_, _00752_);
  and (_13387_, _00759_, _05141_);
  and (_00760_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_00761_, _00760_, _10380_);
  and (_00762_, _00761_, _08280_);
  not (_00763_, _08280_);
  or (_00764_, _00763_, _10375_);
  and (_00765_, _00764_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_00766_, _00765_, _08289_);
  or (_00767_, _00766_, _00762_);
  or (_00768_, _08360_, _05522_);
  and (_00769_, _00768_, _05141_);
  and (_13390_, _00769_, _00767_);
  or (_00770_, _12096_, _12030_);
  and (_00771_, _00770_, _12097_);
  or (_00772_, _00771_, _07135_);
  or (_00773_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00774_, _00773_, _12108_);
  and (_00775_, _00774_, _00772_);
  and (_00776_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_13411_, _00776_, _00775_);
  nand (_00777_, _12099_, _12025_);
  and (_00779_, _00777_, _12100_);
  or (_00780_, _00779_, _07135_);
  or (_00781_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00782_, _00781_, _12108_);
  and (_00783_, _00782_, _00780_);
  and (_00784_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_13431_, _00784_, _00783_);
  nand (_00785_, _12097_, _12027_);
  and (_00786_, _00785_, _12099_);
  or (_00787_, _00786_, _07135_);
  or (_00789_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00790_, _00789_, _12108_);
  and (_00791_, _00790_, _00787_);
  and (_00792_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_13436_, _00792_, _00791_);
  nor (_00793_, _12075_, _12072_);
  nor (_00794_, _00793_, _12077_);
  or (_00795_, _00794_, _07135_);
  or (_00796_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_00797_, _00796_, _12108_);
  and (_00798_, _00797_, _00795_);
  and (_00799_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00147_, _00799_, _00798_);
  nor (_00800_, _12087_, _12084_);
  nor (_00801_, _00800_, _12088_);
  or (_00802_, _00801_, _07135_);
  or (_00803_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00804_, _00803_, _12108_);
  and (_00805_, _00804_, _00802_);
  and (_00806_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00158_, _00806_, _00805_);
  nor (_00808_, _12083_, _12063_);
  nor (_00809_, _00808_, _12084_);
  or (_00810_, _00809_, _07135_);
  or (_00811_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00812_, _00811_, _12108_);
  and (_00813_, _00812_, _00810_);
  and (_00814_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_00172_, _00814_, _00813_);
  and (_00815_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00816_, _12081_, _12078_);
  nor (_00817_, _00816_, _12083_);
  or (_00818_, _00817_, _07135_);
  or (_00819_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00820_, _00819_, _12108_);
  and (_00821_, _00820_, _00818_);
  or (_00209_, _00821_, _00815_);
  nand (_00822_, _00203_, _05960_);
  and (_00823_, _00358_, _00194_);
  nand (_00824_, _00823_, _00193_);
  nor (_00825_, _00824_, _00199_);
  or (_00827_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_00828_, _00408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_00829_, _00828_, _00186_);
  nand (_00830_, _00829_, _00196_);
  or (_00831_, _00830_, _00199_);
  and (_00832_, _00831_, _00827_);
  or (_00833_, _00832_, _00203_);
  and (_00834_, _00833_, _05141_);
  and (_00341_, _00834_, _00822_);
  or (_00835_, _00414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_00836_, _00464_, _05141_);
  and (_00837_, _00836_, _00835_);
  not (_00838_, _00414_);
  and (_00839_, _00410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_00840_, _00839_, _00838_);
  nand (_00841_, _00840_, _00837_);
  nor (_00842_, _00841_, _00203_);
  and (_00343_, _00842_, _00378_);
  nand (_00843_, _00199_, _05960_);
  and (_00844_, _00507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_00845_, _00844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_00846_, _00844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_00847_, _00846_, _00845_);
  and (_00848_, _00847_, _00455_);
  not (_00849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_00850_, _00414_, _00410_);
  and (_00851_, _00850_, _00849_);
  nor (_00852_, _00850_, _00849_);
  or (_00854_, _00852_, _00851_);
  and (_00856_, _00854_, _00464_);
  and (_00857_, _00410_, _00193_);
  or (_00858_, _00857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_00859_, _00858_, _00356_);
  and (_00860_, _00839_, _00193_);
  nor (_00861_, _00860_, _00859_);
  or (_00862_, _00861_, _00856_);
  or (_00864_, _00862_, _00199_);
  or (_00865_, _00864_, _00848_);
  and (_00866_, _00865_, _00204_);
  and (_00867_, _00866_, _00843_);
  and (_00868_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_00869_, _00868_, _00867_);
  and (_00345_, _00869_, _05141_);
  nand (_00870_, _06707_, _06244_);
  or (_00871_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_00872_, _00871_, _05141_);
  and (_00349_, _00872_, _00870_);
  or (_00873_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_00874_, _00873_, _05141_);
  nand (_00875_, _00575_, _05960_);
  and (_00355_, _00875_, _00874_);
  or (_00876_, _12914_, _12773_);
  or (_00877_, _00876_, _05739_);
  nor (_00878_, _12772_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_00879_, _00878_, _12906_);
  and (_00880_, _00879_, _00877_);
  nor (_00881_, _00880_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00882_, _00880_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_00883_, _00882_, _00881_);
  and (_00884_, _00883_, _12973_);
  and (_00885_, _12701_, _07288_);
  and (_00886_, _11451_, _06669_);
  and (_00887_, _12707_, _12776_);
  nand (_00888_, _12726_, _05699_);
  and (_00889_, _00888_, _12727_);
  and (_00891_, _00889_, _12713_);
  or (_00892_, _00891_, _00887_);
  and (_00893_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_00894_, _00893_, _00892_);
  or (_00895_, _00894_, _00886_);
  or (_00896_, _00895_, _00885_);
  or (_00897_, _00896_, _00884_);
  or (_00898_, _00897_, _13052_);
  nor (_00900_, _12955_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_00901_, _00900_, _12956_);
  or (_00902_, _00901_, _12700_);
  and (_00903_, _00902_, _05141_);
  and (_00357_, _00903_, _00898_);
  and (_00366_, t0_i, _05141_);
  and (_00370_, t1_i, _05141_);
  and (_00904_, _13439_, _05960_);
  and (_00905_, _00102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00906_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_00907_, _00906_, _00905_);
  and (_00908_, _00907_, _00038_);
  or (_00909_, _00908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_00910_, _00908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_00912_, _00910_, _00033_);
  and (_00913_, _00912_, _00909_);
  and (_00914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_00915_, _00907_, _00069_);
  or (_00916_, _00915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  not (_00917_, _00048_);
  and (_00918_, _00915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_00919_, _00918_, _00917_);
  and (_00920_, _00919_, _00916_);
  or (_00921_, _00920_, _00914_);
  nor (_00922_, _00921_, _00913_);
  and (_00923_, _00922_, _13375_);
  or (_00924_, _00923_, _00904_);
  nand (_00925_, _00924_, _00060_);
  or (_00926_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_00927_, _00926_, _05141_);
  and (_00374_, _00927_, _00925_);
  and (_00928_, _00233_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  or (_00929_, _00928_, _00860_);
  and (_00930_, _00929_, _00356_);
  or (_00931_, _00928_, _00196_);
  or (_00932_, _00928_, _00839_);
  and (_00933_, _00932_, _00409_);
  and (_00934_, _00933_, _00931_);
  and (_00935_, _00931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_00936_, _00935_, _00934_);
  or (_00937_, _00936_, _00930_);
  nand (_00938_, _00937_, _05141_);
  nor (_00939_, _00938_, _00203_);
  and (_00376_, _00939_, _00378_);
  not (_00940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_00941_, _13389_, _00940_);
  or (_00942_, _00941_, _00918_);
  and (_00943_, _00942_, _00048_);
  or (_00944_, _00941_, _00910_);
  and (_00945_, _00944_, _13372_);
  nand (_00946_, _13389_, _13369_);
  and (_00947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00948_, _00947_, _00946_);
  or (_00949_, _00948_, _13443_);
  or (_00950_, _00949_, _00945_);
  or (_00951_, _00950_, _00943_);
  and (_00952_, _13366_, _13375_);
  and (_00953_, _00952_, _05141_);
  and (_00377_, _00953_, _00951_);
  nor (_00954_, _13400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_00955_, _00954_, _13401_);
  and (_00956_, _00955_, _13374_);
  and (_00957_, _13402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_00958_, _00957_, _00956_);
  and (_00959_, _00958_, _00953_);
  and (_00960_, _13377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_00961_, _00960_, _13366_);
  nor (_00962_, _00060_, _05960_);
  or (_00963_, _00962_, _00961_);
  and (_00964_, _00963_, _05141_);
  or (_00379_, _00964_, _00959_);
  nand (_00965_, _12906_, _12773_);
  and (_00966_, _00965_, _00876_);
  nand (_00967_, _00966_, _05739_);
  or (_00968_, _00966_, _05739_);
  and (_00969_, _00968_, _12973_);
  and (_00970_, _00969_, _00967_);
  and (_00971_, _12701_, _07166_);
  nand (_00972_, _12725_, _05739_);
  and (_00973_, _00972_, _12726_);
  and (_00974_, _00973_, _12713_);
  nor (_00975_, _12703_, _07200_);
  or (_00976_, _00975_, _00974_);
  and (_00977_, _12707_, _12808_);
  and (_00979_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_00981_, _00979_, _00977_);
  or (_00982_, _00981_, _00976_);
  nor (_00983_, _00982_, _00971_);
  nand (_00984_, _00983_, _12700_);
  or (_00985_, _00984_, _00970_);
  nor (_00986_, _12954_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_00988_, _00986_, _12955_);
  or (_00989_, _00988_, _12700_);
  and (_00990_, _00989_, _05141_);
  and (_00387_, _00990_, _00985_);
  and (_00991_, _05568_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_00992_, _05522_, _05291_);
  or (_00993_, _00992_, _05572_);
  or (_00994_, _00993_, _00991_);
  or (_00995_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_00996_, _00995_, _05141_);
  and (_00457_, _00996_, _00994_);
  and (_00997_, _06154_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_00998_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_00999_, _00998_, _06156_);
  and (_01000_, _06180_, _05561_);
  or (_01001_, _01000_, _00999_);
  or (_01002_, _01001_, _00997_);
  and (_00486_, _01002_, _05141_);
  not (_01003_, _12827_);
  and (_01004_, _01003_, _12707_);
  not (_01006_, _07200_);
  and (_01007_, _13058_, _01006_);
  and (_01008_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_01009_, _12713_, _12808_);
  or (_01010_, _01009_, _01008_);
  or (_01011_, _01010_, _01007_);
  nand (_01012_, _12898_, _12896_);
  nand (_01013_, _01012_, _12835_);
  nand (_01014_, _12837_, _01013_);
  or (_01015_, _12837_, _01013_);
  and (_01016_, _01015_, _12940_);
  and (_01017_, _01016_, _01014_);
  or (_01018_, _01017_, _01011_);
  or (_01019_, _01018_, _01004_);
  and (_01020_, _01019_, _12700_);
  nor (_01021_, _00226_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_01022_, _01021_, _00228_);
  nor (_01023_, _01022_, _12700_);
  or (_01024_, _01023_, _01020_);
  and (_00657_, _01024_, _05141_);
  not (_01026_, _07593_);
  and (_01028_, _12707_, _01026_);
  not (_01029_, _07259_);
  and (_01031_, _13058_, _01029_);
  and (_01033_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_01034_, _12713_, _12831_);
  or (_01035_, _01034_, _01033_);
  or (_01036_, _01035_, _01031_);
  or (_01037_, _01036_, _01028_);
  or (_01038_, _12898_, _12896_);
  and (_01039_, _01038_, _01012_);
  and (_01040_, _01039_, _12940_);
  or (_01041_, _01040_, _01037_);
  and (_01042_, _01041_, _12700_);
  nor (_01043_, _07622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_01044_, _01043_, _00226_);
  nor (_01045_, _01044_, _12700_);
  or (_01046_, _01045_, _01042_);
  and (_00660_, _01046_, _05141_);
  not (_01047_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_01048_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_01049_, _01048_, _01047_);
  nor (_01050_, _01049_, rst);
  nand (_01051_, _01048_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_01052_, _01048_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_01053_, _01052_, _01051_);
  and (_00666_, _01053_, _01050_);
  or (_01054_, _12847_, _12848_);
  not (_01055_, _01054_);
  nand (_01056_, _01055_, _12894_);
  or (_01057_, _01055_, _12894_);
  and (_01058_, _01057_, _12973_);
  and (_01059_, _01058_, _01056_);
  not (_01060_, _07350_);
  and (_01061_, _13058_, _01060_);
  not (_01062_, _07572_);
  and (_01063_, _12707_, _01062_);
  and (_01064_, _12713_, _12843_);
  and (_01065_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_01066_, _01065_, _01064_);
  or (_01067_, _01066_, _01063_);
  or (_01068_, _01067_, _01061_);
  or (_01069_, _01068_, _01059_);
  and (_01070_, _01069_, _12700_);
  and (_01071_, _13052_, _07623_);
  or (_01072_, _01071_, _01070_);
  and (_00670_, _01072_, _05141_);
  not (_01073_, _07550_);
  and (_01074_, _12707_, _01073_);
  not (_01075_, _06617_);
  and (_01076_, _13058_, _01075_);
  and (_01077_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_01078_, _12713_, _12849_);
  or (_01079_, _01078_, _01077_);
  or (_01080_, _01079_, _01076_);
  or (_01081_, _12892_, _12889_);
  not (_01082_, _12893_);
  and (_01083_, _12940_, _01082_);
  and (_01084_, _01083_, _01081_);
  or (_01085_, _01084_, _01080_);
  or (_01086_, _01085_, _01074_);
  and (_01087_, _01086_, _12700_);
  and (_01088_, _13052_, _07636_);
  or (_01089_, _01088_, _01087_);
  and (_00684_, _01089_, _05141_);
  not (_01090_, _07434_);
  and (_01091_, _13058_, _01090_);
  not (_01092_, _12876_);
  and (_01093_, _01092_, _12707_);
  and (_01094_, _12713_, _12855_);
  and (_01095_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_01096_, _01095_, _01094_);
  or (_01097_, _01096_, _01093_);
  or (_01098_, _01097_, _01091_);
  nor (_01099_, _12887_, _12884_);
  nor (_01100_, _01099_, _12888_);
  and (_01101_, _01100_, _12940_);
  or (_01102_, _01101_, _01098_);
  or (_01103_, _01102_, _13052_);
  or (_01104_, _12700_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_01105_, _01104_, _05141_);
  and (_00706_, _01105_, _01103_);
  and (_01106_, _12701_, _07378_);
  and (_01107_, _12707_, _12849_);
  nor (_01108_, _12703_, _06617_);
  or (_01109_, _01108_, _01107_);
  and (_01110_, _12713_, _07014_);
  and (_01111_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_01112_, _01111_, _01110_);
  or (_01113_, _01112_, _01109_);
  or (_01114_, _01113_, _01106_);
  nor (_01115_, _12904_, _12772_);
  and (_01116_, _12902_, _12910_);
  nor (_01117_, _01116_, _12773_);
  or (_01118_, _01117_, _01115_);
  nand (_01119_, _01118_, _05455_);
  or (_01120_, _01118_, _05455_);
  and (_01121_, _01120_, _01119_);
  and (_01122_, _01121_, _12940_);
  or (_01123_, _01122_, _01114_);
  or (_01124_, _01123_, _13052_);
  nor (_01125_, _13001_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01126_, _01125_, _13002_);
  or (_01127_, _01126_, _12700_);
  and (_01128_, _01127_, _05141_);
  and (_00778_, _01128_, _01124_);
  and (_01129_, _12701_, _07406_);
  and (_01130_, _12707_, _12855_);
  and (_01131_, _12713_, _06524_);
  or (_01132_, _01131_, _01130_);
  and (_01133_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01134_, _11451_, _01090_);
  or (_01135_, _01134_, _01133_);
  or (_01136_, _01135_, _01132_);
  or (_01137_, _01136_, _01129_);
  and (_01138_, _12902_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_01139_, _01138_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_01140_, _01139_, _01117_);
  and (_01141_, _12903_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_01142_, _01141_, _12904_);
  and (_01143_, _01142_, _12773_);
  or (_01144_, _01143_, _01140_);
  and (_01145_, _01144_, _12940_);
  or (_01146_, _01145_, _01137_);
  or (_01147_, _01146_, _13052_);
  nor (_01148_, _13000_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_01150_, _01148_, _13001_);
  or (_01151_, _01150_, _12700_);
  and (_01152_, _01151_, _05141_);
  and (_00788_, _01152_, _01147_);
  and (_01153_, _12701_, _07466_);
  and (_01154_, _12707_, _12880_);
  and (_01155_, _11451_, _13057_);
  or (_01156_, _01155_, _01154_);
  and (_01157_, _12713_, _06497_);
  and (_01158_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_01159_, _01158_, _01157_);
  or (_01160_, _01159_, _01156_);
  or (_01161_, _01160_, _01153_);
  and (_01162_, _12902_, _05411_);
  nor (_01163_, _12902_, _05411_);
  nor (_01164_, _01163_, _01162_);
  nand (_01165_, _01164_, _12772_);
  or (_01166_, _01164_, _12772_);
  and (_01167_, _01166_, _01165_);
  and (_01168_, _01167_, _12940_);
  nor (_01169_, _01168_, _01161_);
  nand (_01170_, _01169_, _12700_);
  nor (_01171_, _12999_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_01172_, _01171_, _13000_);
  or (_01173_, _01172_, _12700_);
  and (_01174_, _01173_, _05141_);
  and (_00807_, _01174_, _01170_);
  not (_01175_, _06875_);
  and (_01176_, _13058_, _01175_);
  not (_01177_, _12770_);
  and (_01178_, _01177_, _12707_);
  and (_01179_, _12713_, _12732_);
  and (_01180_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_01181_, _01180_, _01179_);
  or (_01182_, _01181_, _01178_);
  or (_01184_, _01182_, _01176_);
  nor (_01185_, _00219_, _12800_);
  nor (_01186_, _01185_, _12802_);
  and (_01187_, _01185_, _12802_);
  or (_01189_, _01187_, _01186_);
  and (_01190_, _01189_, _12940_);
  or (_01191_, _01190_, _01184_);
  and (_01192_, _01191_, _12700_);
  nor (_01193_, _00227_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_01194_, _01193_, _12999_);
  nor (_01195_, _01194_, _12700_);
  or (_01196_, _01195_, _01192_);
  and (_00826_, _01196_, _05141_);
  and (_01197_, _11667_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_01198_, _01197_, _11665_);
  and (_01199_, _01198_, _06013_);
  not (_01200_, _06013_);
  or (_01201_, _06209_, _01200_);
  and (_01202_, _01201_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_01203_, _01202_, _06020_);
  or (_01204_, _01203_, _01199_);
  or (_01205_, _06021_, _06004_);
  and (_01206_, _01205_, _05141_);
  and (_00853_, _01206_, _01204_);
  and (_01208_, _05287_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01209_, _01208_, _10356_);
  and (_01210_, _01209_, _06013_);
  nand (_01211_, _06013_, _08283_);
  and (_01212_, _01211_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01213_, _01212_, _06020_);
  or (_01214_, _01213_, _01210_);
  nand (_01215_, _06020_, _05560_);
  and (_01216_, _01215_, _05141_);
  and (_00863_, _01216_, _01214_);
  and (_01217_, _11667_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_01218_, _01217_, _11665_);
  and (_01219_, _01218_, _06255_);
  not (_01220_, _06255_);
  or (_01221_, _01220_, _06209_);
  and (_01222_, _01221_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_01223_, _01222_, _06262_);
  or (_01224_, _01223_, _01219_);
  or (_01225_, _06263_, _06004_);
  and (_01226_, _01225_, _05141_);
  and (_00890_, _01226_, _01224_);
  and (_01227_, _05287_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_01228_, _01227_, _10356_);
  and (_01229_, _01228_, _06255_);
  nand (_01230_, _06255_, _08283_);
  and (_01231_, _01230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_01232_, _01231_, _06262_);
  or (_01233_, _01232_, _01229_);
  nand (_01234_, _06262_, _05560_);
  and (_01235_, _01234_, _05141_);
  and (_00899_, _01235_, _01233_);
  or (_01236_, \oc8051_top_1.oc8051_sfr1.prescaler [2], rst);
  nor (_00911_, _01236_, _01051_);
  and (_00978_, _00640_, _06065_);
  not (_01237_, _06114_);
  nor (_01238_, _06102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_01239_, _01238_, _06100_);
  or (_01240_, _01239_, _06105_);
  and (_01241_, _01240_, _01237_);
  or (_01242_, _01241_, _06112_);
  and (_01243_, _06133_, _06110_);
  and (_01244_, _01243_, _01242_);
  not (_01245_, _06078_);
  or (_01246_, _06089_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01247_, _01246_, _06085_);
  or (_01248_, _01247_, _06093_);
  and (_01249_, _01248_, _01245_);
  or (_01250_, _01249_, _06076_);
  and (_01251_, _06097_, _06074_);
  and (_01252_, _01251_, _01250_);
  or (_01253_, _01252_, _06065_);
  or (_01254_, _01253_, _01244_);
  or (_01255_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01256_, _01255_, _05141_);
  and (_00980_, _01256_, _01254_);
  and (_01257_, _06878_, _06009_);
  and (_01258_, _01257_, _06008_);
  nand (_01259_, _01258_, _05963_);
  or (_01260_, _01258_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_01261_, _01260_, _05647_);
  and (_01262_, _01261_, _01259_);
  and (_01263_, _06261_, _05272_);
  not (_01264_, _01263_);
  nor (_01265_, _01264_, _05960_);
  and (_01266_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_01267_, _01266_, _01265_);
  and (_01268_, _01267_, _05925_);
  and (_01269_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_01270_, _01269_, rst);
  or (_01271_, _01270_, _01268_);
  or (_00987_, _01271_, _01262_);
  and (_01272_, _06205_, _05210_);
  nand (_01273_, _01272_, _05963_);
  or (_01274_, _01272_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_01275_, _01274_, _05928_);
  and (_01276_, _01275_, _01273_);
  and (_01277_, _05927_, _06703_);
  or (_01278_, _01277_, _01276_);
  and (_01005_, _01278_, _05141_);
  and (_01279_, _12559_, _12502_);
  nand (_01280_, _12397_, _12391_);
  and (_01281_, _01280_, _12450_);
  and (_01282_, _12261_, _12310_);
  and (_01283_, _01282_, _01281_);
  and (_01284_, _12608_, _12372_);
  and (_01285_, _01284_, _01283_);
  and (_01286_, _01285_, _01279_);
  and (_01287_, _01286_, _06619_);
  and (_01288_, _12557_, _12502_);
  and (_01289_, _12610_, _12374_);
  and (_01290_, _01289_, _01288_);
  and (_01291_, _01280_, _12448_);
  and (_01292_, _01291_, _01282_);
  and (_01293_, _01292_, _01290_);
  and (_01294_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_01295_, _12608_, _12374_);
  and (_01296_, _01288_, _01295_);
  and (_01297_, _01296_, _01292_);
  and (_01298_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_01299_, _01298_, _01294_);
  and (_01300_, _01279_, _01295_);
  and (_01301_, _01300_, _01292_);
  and (_01302_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_01303_, _12557_, _12504_);
  and (_01304_, _01303_, _01289_);
  and (_01305_, _01304_, _01292_);
  and (_01306_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_01307_, _01306_, _01302_);
  or (_01308_, _01307_, _01299_);
  and (_01309_, _12559_, _12504_);
  and (_01310_, _01295_, _01309_);
  and (_01311_, _01292_, _01310_);
  and (_01312_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_01313_, _01296_, _01283_);
  and (_01314_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_01315_, _01314_, _01312_);
  not (_01316_, _01296_);
  nand (_01317_, _01281_, _12313_);
  or (_01318_, _01317_, _12263_);
  nor (_01319_, _01318_, _01316_);
  and (_01320_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_01321_, _12263_, _12313_);
  and (_01322_, _01321_, _01281_);
  and (_01323_, _01309_, _12610_);
  and (_01324_, _01323_, _12372_);
  and (_01325_, _01324_, _01322_);
  and (_01326_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_01327_, _01326_, _01320_);
  or (_01328_, _01327_, _01315_);
  or (_01329_, _01328_, _01308_);
  and (_01330_, _01310_, _01283_);
  and (_01331_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_01332_, _01303_, _01295_);
  and (_01333_, _01332_, _01283_);
  and (_01334_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_01335_, _01334_, _01331_);
  and (_01336_, _01300_, _01283_);
  and (_01337_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_01338_, _01304_, _01283_);
  and (_01339_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_01340_, _01339_, _01337_);
  or (_01341_, _01340_, _01335_);
  nand (_01342_, _01281_, _12310_);
  nor (_01343_, _01342_, _12261_);
  and (_01344_, _01343_, _01296_);
  and (_01345_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_01346_, _01343_, _01332_);
  and (_01347_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_01348_, _01347_, _01345_);
  and (_01349_, _01290_, _01283_);
  and (_01350_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_01351_, _01324_, _01283_);
  and (_01352_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_01353_, _01352_, _01350_);
  or (_01354_, _01353_, _01348_);
  or (_01355_, _01354_, _01341_);
  or (_01356_, _01355_, _01329_);
  and (_01357_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_01358_, _01284_, _01309_);
  and (_01359_, _01358_, _01283_);
  and (_01360_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01361_, _01360_, _01357_);
  and (_01362_, _01291_, _12313_);
  and (_01363_, _01284_, _01288_);
  and (_01364_, _01363_, _12263_);
  and (_01365_, _01364_, _01362_);
  and (_01366_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_01367_, _01303_, _01284_);
  and (_01368_, _01367_, _01283_);
  and (_01369_, _01368_, _12390_);
  or (_01370_, _01369_, _01366_);
  or (_01371_, _01370_, _01361_);
  not (_01372_, _01363_);
  nor (_01373_, _01318_, _01372_);
  and (_01374_, _07053_, _06417_);
  or (_01375_, _01374_, _06563_);
  or (_01376_, _01375_, _06777_);
  and (_01377_, _01376_, _06773_);
  not (_01378_, _01377_);
  and (_01379_, _06755_, _06564_);
  or (_01380_, _01379_, _07073_);
  or (_01381_, _01380_, _12130_);
  or (_01382_, _06779_, _06772_);
  and (_01383_, _07074_, _06574_);
  or (_01384_, _12136_, _01383_);
  or (_01385_, _01384_, _01382_);
  or (_01386_, _01385_, _07056_);
  nor (_01387_, _01386_, _01381_);
  and (_01388_, _01387_, _01378_);
  and (_01390_, _01388_, _12123_);
  nor (_01391_, _01390_, _08330_);
  or (_01393_, _01391_, p2_in[7]);
  not (_01394_, _01391_);
  or (_01396_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_01397_, _01396_, _01393_);
  and (_01398_, _01397_, _01373_);
  and (_01399_, _01322_, _01363_);
  or (_01400_, _01391_, p3_in[7]);
  or (_01401_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_01402_, _01401_, _01400_);
  and (_01403_, _01402_, _01399_);
  or (_01404_, _01403_, _01398_);
  and (_01405_, _01363_, _01283_);
  or (_01406_, _01391_, p0_in[7]);
  or (_01407_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_01408_, _01407_, _01406_);
  and (_01409_, _01408_, _01405_);
  or (_01410_, _01391_, p1_in[7]);
  or (_01411_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_01412_, _01411_, _01410_);
  and (_01413_, _01343_, _01363_);
  and (_01414_, _01413_, _01412_);
  or (_01415_, _01414_, _01409_);
  or (_01416_, _01415_, _01404_);
  or (_01417_, _01416_, _01371_);
  and (_01418_, _01363_, _01280_);
  or (_01419_, _12450_, _12313_);
  or (_01420_, _01419_, _12261_);
  not (_01421_, _01420_);
  and (_01422_, _01421_, _01418_);
  and (_01423_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_01424_, _01363_, _12261_);
  and (_01425_, _01424_, _01362_);
  and (_01426_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_01427_, _01426_, _01423_);
  or (_01428_, _01427_, _01417_);
  or (_01429_, _01428_, _01356_);
  nand (_01430_, _01422_, _12690_);
  nand (_01431_, _01285_, _01309_);
  or (_01432_, _01431_, _07138_);
  and (_01433_, _01432_, _01430_);
  or (_01434_, _01433_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_01435_, _06010_);
  nor (_01436_, _01323_, _01435_);
  nand (_01437_, _01436_, _12455_);
  nand (_01438_, _01425_, _08161_);
  and (_01439_, _01438_, _01437_);
  and (_01440_, _01439_, _12617_);
  and (_01441_, _01440_, _01434_);
  and (_01442_, _01441_, _01429_);
  not (_01443_, _01441_);
  nor (_01444_, _01297_, _01293_);
  nor (_01445_, _01305_, _01301_);
  and (_01446_, _01445_, _01444_);
  nor (_01447_, _01313_, _01311_);
  nor (_01448_, _01325_, _01319_);
  and (_01449_, _01448_, _01447_);
  and (_01450_, _01449_, _01446_);
  nor (_01452_, _01346_, _01344_);
  nor (_01453_, _01351_, _01349_);
  and (_01454_, _01453_, _01452_);
  nor (_01455_, _01333_, _01330_);
  nor (_01456_, _01338_, _01336_);
  and (_01457_, _01456_, _01455_);
  and (_01458_, _01457_, _01454_);
  and (_01460_, _01458_, _01450_);
  nor (_01461_, _01425_, _01422_);
  nor (_01462_, _01359_, _01286_);
  nor (_01463_, _01368_, _01365_);
  and (_01464_, _01463_, _01462_);
  nor (_01466_, _01399_, _01373_);
  nor (_01468_, _01413_, _01405_);
  and (_01469_, _01468_, _01466_);
  and (_01470_, _01469_, _01464_);
  and (_01471_, _01470_, _01461_);
  and (_01472_, _01471_, _01460_);
  or (_01474_, _01472_, _01443_);
  and (_01475_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_01476_, _01475_, _01442_);
  or (_01477_, _01476_, _01287_);
  nand (_01478_, _01287_, _06875_);
  and (_01480_, _01478_, _05141_);
  and (_01025_, _01480_, _01477_);
  and (_01481_, _06004_, _05277_);
  and (_01482_, _08484_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_01483_, _01482_, _05572_);
  or (_01485_, _01483_, _01481_);
  or (_01486_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_01487_, _01486_, _05141_);
  and (_01027_, _01487_, _01485_);
  and (_01488_, _06013_, _06207_);
  nand (_01489_, _01488_, _05963_);
  or (_01490_, _01488_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_01491_, _01490_, _01489_);
  or (_01492_, _01491_, _06020_);
  nand (_01493_, _06244_, _06020_);
  and (_01494_, _01493_, _05141_);
  and (_01030_, _01494_, _01492_);
  and (_01495_, _06255_, _06207_);
  nand (_01496_, _01495_, _05963_);
  or (_01497_, _01495_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_01498_, _01497_, _06263_);
  and (_01499_, _01498_, _01496_);
  nor (_01501_, _06263_, _06244_);
  or (_01502_, _01501_, _01499_);
  and (_01032_, _01502_, _05141_);
  and (_01504_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_01505_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_01506_, _01505_, _01504_);
  and (_01507_, _01506_, _08355_);
  and (_01508_, _08348_, _05522_);
  or (_01509_, _01508_, _01507_);
  and (_01149_, _01509_, _05141_);
  and (_01510_, _06281_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_01512_, _06275_, _06179_);
  or (_01513_, _01512_, _01510_);
  and (_01183_, _01513_, _05141_);
  nor (_01514_, _06121_, _06065_);
  and (_01515_, _06065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_01517_, _01515_, _01514_);
  and (_01389_, _01517_, _05141_);
  not (_01518_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_01519_, _06089_, _05630_);
  or (_01520_, _01519_, _01518_);
  nor (_01521_, _06085_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_01522_, _01521_, _06093_);
  nand (_01524_, _01522_, _01520_);
  or (_01525_, _06094_, _05629_);
  and (_01526_, _01525_, _01524_);
  or (_01527_, _01526_, _06078_);
  not (_01528_, _06076_);
  or (_01529_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _05630_);
  or (_01530_, _01529_, _01245_);
  and (_01531_, _01530_, _01528_);
  and (_01532_, _01531_, _01527_);
  and (_01533_, _06076_, _05629_);
  or (_01534_, _01533_, _06073_);
  or (_01535_, _01534_, _01532_);
  or (_01536_, _01529_, _06074_);
  and (_01537_, _01536_, _01535_);
  or (_01538_, _01537_, _06123_);
  and (_01539_, _06102_, _05630_);
  or (_01541_, _01539_, _01518_);
  and (_01542_, _06100_, _05630_);
  nor (_01544_, _01542_, _06105_);
  nand (_01546_, _01544_, _01541_);
  or (_01547_, _06106_, _05629_);
  and (_01549_, _01547_, _01546_);
  or (_01550_, _01549_, _06114_);
  not (_01551_, _06112_);
  or (_01552_, _01529_, _01237_);
  and (_01554_, _01552_, _01551_);
  and (_01555_, _01554_, _01550_);
  and (_01556_, _06112_, _05629_);
  or (_01557_, _01556_, _06109_);
  or (_01558_, _01557_, _01555_);
  or (_01559_, _01529_, _06110_);
  and (_01560_, _01559_, _01558_);
  or (_01561_, _01560_, _06134_);
  and (_01562_, _01561_, _01538_);
  or (_01563_, _01562_, _06065_);
  or (_01565_, _01514_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_01566_, _01565_, _05141_);
  and (_01392_, _01566_, _01563_);
  and (_01567_, _06205_, _06620_);
  nand (_01568_, _01567_, _05963_);
  or (_01569_, _01567_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_01570_, _01569_, _05928_);
  and (_01571_, _01570_, _01568_);
  nor (_01572_, _05928_, _05560_);
  or (_01573_, _01572_, _01571_);
  and (_01395_, _01573_, _05141_);
  and (_01451_, _11861_, _05141_);
  or (_01574_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _05630_);
  and (_01575_, _01574_, _06110_);
  or (_01576_, _01575_, _06116_);
  and (_01577_, _06105_, _05639_);
  not (_01579_, _06115_);
  or (_01580_, _01539_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01581_, _01580_, _01544_);
  or (_01583_, _01581_, _01579_);
  or (_01584_, _01583_, _01577_);
  and (_01586_, _01584_, _01576_);
  and (_01587_, _06109_, _05639_);
  or (_01588_, _01587_, _06119_);
  or (_01589_, _01588_, _01586_);
  or (_01590_, _06120_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01591_, _01590_, _01589_);
  and (_01592_, _01591_, _06123_);
  and (_01593_, _01574_, _06074_);
  or (_01594_, _01593_, _06081_);
  and (_01595_, _06093_, _05639_);
  or (_01596_, _01519_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nand (_01597_, _01596_, _01522_);
  nand (_01598_, _01597_, _06080_);
  or (_01599_, _01598_, _01595_);
  and (_01600_, _01599_, _01594_);
  and (_01601_, _06073_, _05639_);
  or (_01602_, _01601_, _01600_);
  and (_01603_, _01602_, _06097_);
  or (_01604_, _01603_, _06065_);
  or (_01605_, _01604_, _01592_);
  or (_01606_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01607_, _01606_, _05141_);
  and (_01459_, _01607_, _01605_);
  and (_01608_, _06205_, _08469_);
  or (_01609_, _01608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_01610_, _01609_, _05928_);
  nand (_01611_, _01608_, _05963_);
  and (_01612_, _01611_, _01610_);
  and (_01613_, _05927_, _05522_);
  or (_01614_, _01613_, _01612_);
  and (_01465_, _01614_, _05141_);
  and (_01467_, _06391_, _05141_);
  and (_01473_, _13350_, _06065_);
  and (_01615_, _06065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_01616_, _01615_, _01514_);
  and (_01479_, _01616_, _05141_);
  nand (_01617_, _06117_, _06141_);
  nor (_01618_, _01617_, _06097_);
  and (_01619_, _06065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor (_01620_, _06093_, _06071_);
  not (_01621_, _06081_);
  nor (_01622_, _06091_, _01621_);
  and (_01623_, _01622_, _01620_);
  and (_01624_, _01623_, _06066_);
  or (_01625_, _01624_, _01619_);
  or (_01627_, _01625_, _01618_);
  and (_01484_, _01627_, _05141_);
  or (_01628_, _06093_, _06078_);
  and (_01629_, _06091_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_01630_, _01629_, _01628_);
  and (_01631_, _01630_, _01528_);
  and (_01632_, _01631_, _01251_);
  nor (_01633_, _06112_, _06109_);
  or (_01634_, _06114_, _06105_);
  and (_01635_, _06103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_01636_, _01635_, _01634_);
  and (_01637_, _01636_, _01633_);
  and (_01638_, _01637_, _06133_);
  or (_01639_, _01638_, _06065_);
  or (_01640_, _01639_, _01632_);
  or (_01641_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_01642_, _01641_, _05141_);
  and (_01500_, _01642_, _01640_);
  nor (_01643_, _06097_, _06065_);
  or (_01644_, _01643_, _05630_);
  nand (_01645_, _06247_, _06121_);
  and (_01646_, _01645_, _05141_);
  and (_01503_, _01646_, _01644_);
  or (_01647_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01648_, _01647_, _05141_);
  or (_01649_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01650_, _01649_, _06074_);
  or (_01652_, _01650_, _06081_);
  and (_01653_, _06089_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_01654_, _01653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor (_01655_, _06085_, _05630_);
  nor (_01656_, _01655_, _06093_);
  and (_01657_, _01656_, _01654_);
  nand (_01658_, _06093_, _05640_);
  nand (_01659_, _01658_, _06080_);
  or (_01660_, _01659_, _01657_);
  and (_01661_, _01660_, _01652_);
  and (_01662_, _06073_, _05640_);
  or (_01663_, _01662_, _01661_);
  and (_01664_, _01663_, _06097_);
  and (_01665_, _01649_, _06110_);
  or (_01666_, _01665_, _06116_);
  and (_01667_, _06105_, _05640_);
  and (_01668_, _06100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_01669_, _01668_, _06105_);
  and (_01670_, _06102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_01671_, _01670_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01672_, _01671_, _01669_);
  or (_01673_, _01672_, _01579_);
  or (_01674_, _01673_, _01667_);
  and (_01675_, _01674_, _01666_);
  and (_01676_, _06109_, _05640_);
  or (_01677_, _01676_, _06119_);
  or (_01678_, _01677_, _01675_);
  or (_01679_, _06120_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01680_, _01679_, _01678_);
  and (_01682_, _01680_, _06123_);
  or (_01683_, _01682_, _01664_);
  or (_01684_, _01683_, _06065_);
  and (_01511_, _01684_, _01648_);
  not (_01685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor (_01686_, _01514_, _01685_);
  or (_01687_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_01688_, _01687_, _06074_);
  and (_01689_, _01688_, _06097_);
  or (_01690_, _01653_, _01685_);
  nand (_01691_, _01690_, _01656_);
  or (_01692_, _06094_, _05631_);
  and (_01693_, _01692_, _01691_);
  or (_01694_, _01693_, _06078_);
  or (_01695_, _01687_, _01245_);
  and (_01696_, _01695_, _01528_);
  and (_01697_, _01696_, _01694_);
  and (_01698_, _06076_, _05631_);
  or (_01699_, _01698_, _06073_);
  or (_01700_, _01699_, _01697_);
  and (_01701_, _01700_, _01689_);
  or (_01702_, _01670_, _01685_);
  nand (_01703_, _01702_, _01669_);
  or (_01704_, _06106_, _05631_);
  and (_01705_, _01704_, _01703_);
  or (_01706_, _01705_, _06114_);
  or (_01707_, _01687_, _01237_);
  and (_01708_, _01707_, _01551_);
  and (_01709_, _01708_, _01706_);
  and (_01710_, _06112_, _05631_);
  or (_01711_, _01710_, _06109_);
  or (_01712_, _01711_, _01709_);
  or (_01713_, _01687_, _06110_);
  and (_01714_, _01713_, _06133_);
  and (_01715_, _01714_, _01712_);
  or (_01716_, _01715_, _01701_);
  and (_01717_, _01716_, _06066_);
  or (_01718_, _01717_, _01686_);
  and (_01516_, _01718_, _05141_);
  nand (_01719_, _06247_, _06133_);
  and (_01720_, _06247_, _06097_);
  or (_01721_, _01720_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and (_01722_, _01721_, _05141_);
  and (_01523_, _01722_, _01719_);
  nand (_01723_, _06137_, _06133_);
  and (_01724_, _06137_, _06097_);
  or (_01725_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and (_01726_, _01725_, _05141_);
  and (_01540_, _01726_, _01723_);
  and (_01727_, _06255_, _05288_);
  nand (_01728_, _01727_, _05963_);
  or (_01729_, _01727_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_01730_, _01729_, _06263_);
  and (_01731_, _01730_, _01728_);
  nor (_01732_, _06263_, _06178_);
  or (_01734_, _01732_, _01731_);
  and (_01543_, _01734_, _05141_);
  and (_01735_, _06255_, _05210_);
  and (_01736_, _01735_, _05963_);
  nor (_01737_, _01735_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_01738_, _01737_, _01736_);
  nand (_01739_, _01738_, _06263_);
  nand (_01740_, _06262_, _05604_);
  and (_01741_, _01740_, _05141_);
  and (_01545_, _01741_, _01739_);
  and (_01742_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01743_, _01742_, _10380_);
  and (_01744_, _01743_, _06255_);
  or (_01745_, _01220_, _10375_);
  and (_01746_, _01745_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01747_, _01746_, _06262_);
  or (_01748_, _01747_, _01744_);
  or (_01749_, _06263_, _05522_);
  and (_01750_, _01749_, _05141_);
  and (_01548_, _01750_, _01748_);
  and (_01751_, _08283_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_01752_, _01751_, _08281_);
  and (_01753_, _01752_, _06255_);
  nand (_01754_, _06255_, _05186_);
  and (_01755_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_01757_, _01755_, _06262_);
  or (_01759_, _01757_, _01753_);
  nand (_01760_, _06262_, _06062_);
  and (_01761_, _01760_, _05141_);
  and (_01553_, _01761_, _01759_);
  and (_01564_, _06532_, _05141_);
  and (_01763_, _06283_, _06180_);
  and (_01765_, _06154_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_01766_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_01767_, _01766_, _06156_);
  or (_01768_, _01767_, _01765_);
  or (_01769_, _01768_, _01763_);
  and (_01578_, _01769_, _05141_);
  or (_01770_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_01771_, pc_log_change, _05411_);
  and (_01772_, _01771_, _05141_);
  and (_01582_, _01772_, _01770_);
  and (_01773_, _06013_, _05288_);
  nand (_01774_, _01773_, _05963_);
  or (_01775_, _01773_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_01776_, _01775_, _06021_);
  and (_01777_, _01776_, _01774_);
  nor (_01778_, _06178_, _06021_);
  or (_01780_, _01778_, _01777_);
  and (_01585_, _01780_, _05141_);
  or (_01781_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand (_01782_, _07619_, _06379_);
  and (_01784_, _01782_, _05141_);
  and (_01626_, _01784_, _01781_);
  nand (_01785_, _06875_, _06624_);
  or (_01786_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_01787_, _01786_, _05141_);
  and (_01651_, _01787_, _01785_);
  and (_01788_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_01789_, _01788_, _06683_);
  not (_01790_, _01789_);
  and (_01791_, _00626_, _08295_);
  nor (_01792_, _01791_, _06685_);
  nor (_01793_, _09785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  not (_01794_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_01795_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01794_);
  and (_01796_, _01795_, _01793_);
  nor (_01797_, _01796_, _06686_);
  and (_01798_, _01797_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_01799_, _01798_, _01792_);
  and (_01800_, _01799_, _01790_);
  and (_01801_, _01796_, _06685_);
  nor (_01802_, _01801_, _01789_);
  not (_01803_, _01802_);
  nand (_01804_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_01805_, _01804_, _06715_);
  or (_01681_, _01805_, _01800_);
  or (_01806_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand (_01807_, _07619_, _06403_);
  and (_01808_, _01807_, _05141_);
  and (_01733_, _01808_, _01806_);
  and (_01809_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_01810_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_01811_, pc_log_change, _01810_);
  or (_01812_, _01811_, _01809_);
  and (_01756_, _01812_, _05141_);
  and (_01813_, _06013_, _05210_);
  nand (_01814_, _01813_, _05963_);
  or (_01815_, _01813_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_01816_, _01815_, _01814_);
  or (_01817_, _01816_, _06020_);
  nand (_01818_, _06020_, _05604_);
  and (_01819_, _01818_, _05141_);
  and (_01758_, _01819_, _01817_);
  and (_01820_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01821_, _01820_, _10380_);
  and (_01822_, _01821_, _06013_);
  or (_01823_, _10375_, _01200_);
  and (_01825_, _01823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01826_, _01825_, _06020_);
  or (_01827_, _01826_, _01822_);
  or (_01828_, _06021_, _05522_);
  and (_01829_, _01828_, _05141_);
  and (_01762_, _01829_, _01827_);
  nor (_01830_, _08282_, _06104_);
  or (_01831_, _01830_, _08281_);
  and (_01832_, _01831_, _06013_);
  nand (_01833_, _06013_, _05186_);
  and (_01834_, _01833_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_01835_, _01834_, _06020_);
  or (_01836_, _01835_, _01832_);
  nand (_01837_, _06062_, _06020_);
  and (_01838_, _01837_, _05141_);
  and (_01764_, _01838_, _01836_);
  and (_01839_, _10346_, _06032_);
  nand (_01840_, _01839_, _05963_);
  or (_01841_, _01839_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_01843_, _01841_, _10355_);
  nand (_01844_, _01843_, _01840_);
  nand (_01845_, _01844_, _11860_);
  and (_01779_, _01845_, _05141_);
  and (_01846_, _06293_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_01847_, _06766_, _06550_);
  or (_01848_, _13288_, _12117_);
  or (_01849_, _01848_, _01847_);
  or (_01850_, _01374_, _06996_);
  not (_01851_, _07054_);
  or (_01852_, _01851_, _06772_);
  or (_01854_, _01852_, _01850_);
  or (_01855_, _01854_, _01849_);
  or (_01856_, _01855_, _06780_);
  and (_01857_, _07069_, _06546_);
  or (_01858_, _01383_, _01857_);
  or (_01859_, _11431_, _06980_);
  or (_01861_, _01859_, _01858_);
  or (_01862_, _01861_, _06764_);
  and (_01864_, _06565_, _06420_);
  or (_01865_, _12114_, _07037_);
  or (_01866_, _01865_, _01864_);
  and (_01867_, _06556_, _06536_);
  and (_01869_, _06552_, _06536_);
  or (_01870_, _01869_, _01867_);
  and (_01872_, _06755_, _07053_);
  or (_01873_, _01872_, _01870_);
  or (_01875_, _01873_, _01866_);
  or (_01876_, _01875_, _01862_);
  or (_01877_, _01876_, _01856_);
  and (_01878_, _01877_, _06296_);
  or (_01783_, _01878_, _01846_);
  or (_01879_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand (_01880_, _07619_, _06514_);
  and (_01881_, _01880_, _05141_);
  and (_01824_, _01881_, _01879_);
  and (_01882_, _05563_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_01884_, _06290_, _05523_);
  or (_01885_, _01884_, _01882_);
  and (_01842_, _01885_, _05141_);
  nand (_01887_, _06743_, _05960_);
  and (_01889_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_01891_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_01892_, _01891_, _01889_);
  or (_01893_, _01892_, _06743_);
  and (_01894_, _01893_, _05141_);
  and (_01853_, _01894_, _01887_);
  or (_01895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_01896_, _01895_, _11458_);
  and (_01897_, _05922_, _06008_);
  not (_01898_, _06008_);
  nand (_01899_, _01898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_01900_, _01899_, _11458_);
  or (_01901_, _01900_, _01897_);
  and (_01902_, _01901_, _01896_);
  or (_01903_, _01902_, _11462_);
  nand (_01904_, _11462_, _05960_);
  and (_01905_, _01904_, _05141_);
  and (_01860_, _01905_, _01903_);
  nor (_01906_, _11727_, _11651_);
  and (_01907_, _11727_, _08439_);
  and (_01908_, _08462_, _06726_);
  and (_01909_, _01908_, _08457_);
  and (_01910_, _01909_, _01907_);
  or (_01911_, _01910_, _01906_);
  and (_01863_, _01911_, _05141_);
  nand (_01912_, _11726_, _05960_);
  or (_01913_, _11830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_01914_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_01915_, _01914_, _08439_);
  nand (_01916_, _01915_, _08457_);
  and (_01918_, _01916_, _01913_);
  or (_01919_, _01918_, _08463_);
  nor (_01920_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor (_01922_, _01920_, _08471_);
  and (_01923_, _01922_, _01919_);
  nor (_01924_, _11726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor (_01925_, _01924_, _11727_);
  or (_01926_, _01925_, _01923_);
  and (_01928_, _01926_, _05141_);
  and (_01868_, _01928_, _01912_);
  nor (_01929_, _11902_, _05960_);
  and (_01930_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_01931_, _01930_, _08457_);
  nor (_01932_, _08452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor (_01933_, _01932_, _08453_);
  or (_01934_, _01933_, _13159_);
  or (_01935_, _01934_, _01931_);
  or (_01936_, _08439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_01937_, _01936_, _01935_);
  or (_01938_, _01937_, _08463_);
  nor (_01939_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor (_01940_, _01939_, _08471_);
  and (_01941_, _01940_, _01938_);
  or (_01942_, _01941_, _08478_);
  or (_01943_, _01942_, _01929_);
  or (_01944_, _08479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_01945_, _01944_, _05141_);
  and (_01871_, _01945_, _01943_);
  not (_01946_, _08457_);
  and (_01947_, _01907_, _08460_);
  nand (_01948_, _01947_, _01946_);
  or (_01949_, _01947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_01950_, _01949_, _05141_);
  and (_01874_, _01950_, _01948_);
  and (_01883_, t2_i, _05141_);
  nand (_01951_, _06738_, _05960_);
  and (_01952_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_01953_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_01954_, _01953_, _01952_);
  or (_01955_, _01954_, _06738_);
  and (_01956_, _01955_, _06745_);
  and (_01957_, _01956_, _01951_);
  and (_01958_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_01959_, _01958_, _01957_);
  and (_01886_, _01959_, _05141_);
  and (_01888_, t2ex_i, _05141_);
  and (_01890_, _06531_, _05141_);
  nor (_01960_, t2ex_i, rst);
  and (_01917_, _01960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  nor (_01961_, t2_i, rst);
  and (_01921_, _01961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  and (_01962_, _06283_, _05523_);
  and (_01963_, _05303_, _05297_);
  or (_01964_, _01963_, _05299_);
  and (_01965_, _01964_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_01966_, _01965_, _01962_);
  and (_01927_, _01966_, _05141_);
  and (_01967_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_01968_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_01969_, pc_log_change, _01968_);
  or (_01970_, _01969_, _01967_);
  and (_02067_, _01970_, _05141_);
  or (_01971_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_01972_, pc_log_change, _05436_);
  and (_01973_, _01972_, _05141_);
  and (_02103_, _01973_, _01971_);
  nor (_01974_, _05560_, _08484_);
  and (_01975_, _08484_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_01976_, _01975_, _01974_);
  or (_01977_, _01976_, _05572_);
  or (_01978_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_01979_, _01978_, _05141_);
  and (_02137_, _01979_, _01977_);
  nand (_01980_, _06678_, _06244_);
  or (_01981_, _06678_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_01982_, _01981_, _05141_);
  and (_02194_, _01982_, _01980_);
  or (_01983_, _06975_, _07138_);
  nor (_01984_, _07169_, _06875_);
  and (_01985_, _07169_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01986_, _01985_, _06619_);
  or (_01987_, _01986_, _01984_);
  and (_01988_, _01987_, _05141_);
  and (_02221_, _01988_, _01983_);
  and (_01989_, _00690_, _10407_);
  nand (_01990_, _01989_, _05963_);
  or (_01991_, _01989_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01992_, _01991_, _05647_);
  and (_01993_, _01992_, _01990_);
  not (_01994_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_01995_, _05646_, _01994_);
  nand (_01996_, _00698_, _07200_);
  or (_01997_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01998_, _01997_, _05925_);
  and (_01999_, _01998_, _01996_);
  or (_02000_, _01999_, _01995_);
  or (_02001_, _02000_, _01993_);
  and (_02394_, _02001_, _05141_);
  nand (_02002_, _00690_, _08283_);
  and (_02003_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_02004_, _05287_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_02005_, _02004_, _10356_);
  and (_02006_, _02005_, _00690_);
  or (_02007_, _02006_, _02003_);
  and (_02008_, _02007_, _05647_);
  and (_02009_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_02010_, _00698_, _06617_);
  or (_02011_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_02012_, _02011_, _05925_);
  and (_02013_, _02012_, _02010_);
  or (_02014_, _02013_, _02009_);
  or (_02015_, _02014_, _02008_);
  and (_02397_, _02015_, _05141_);
  nor (_02429_, _12304_, rst);
  nand (_02431_, _12463_, _05141_);
  and (_02016_, _10342_, _06009_);
  and (_02017_, _02016_, _05210_);
  nand (_02018_, _02017_, _05963_);
  or (_02019_, _02017_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_02020_, _02019_, _05647_);
  and (_02021_, _02020_, _02018_);
  and (_02022_, _06017_, _05272_);
  and (_02023_, _02022_, _06703_);
  not (_02024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_02025_, _02022_, _02024_);
  or (_02026_, _02025_, _02023_);
  and (_02027_, _02026_, _05925_);
  nor (_02028_, _05646_, _02024_);
  or (_02029_, _02028_, rst);
  or (_02030_, _02029_, _02027_);
  or (_02493_, _02030_, _02021_);
  and (_02031_, _01257_, _06207_);
  nand (_02032_, _02031_, _05963_);
  or (_02033_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_02034_, _02033_, _05647_);
  and (_02035_, _02034_, _02032_);
  nor (_02036_, _01264_, _06244_);
  and (_02037_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02038_, _02037_, _02036_);
  and (_02039_, _02038_, _05925_);
  and (_02040_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02041_, _02040_, rst);
  or (_02042_, _02041_, _02039_);
  or (_02495_, _02042_, _02035_);
  and (_02043_, _10342_, _06202_);
  and (_02044_, _02043_, _06620_);
  nand (_02045_, _02044_, _05963_);
  or (_02046_, _02044_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_02047_, _02046_, _05647_);
  and (_02048_, _02047_, _02045_);
  and (_02049_, _08241_, _05272_);
  nand (_02050_, _02049_, _05560_);
  or (_02051_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_02052_, _02051_, _05925_);
  and (_02053_, _02052_, _02050_);
  and (_02054_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_02055_, _02054_, rst);
  or (_02056_, _02055_, _02053_);
  or (_02499_, _02056_, _02048_);
  or (_02057_, _01264_, _05922_);
  or (_02058_, _01263_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_02059_, _02058_, _05647_);
  and (_02060_, _02059_, _02057_);
  and (_02061_, _01263_, _06703_);
  not (_02062_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_02063_, _01263_, _02062_);
  or (_02064_, _02063_, _02061_);
  and (_02065_, _02064_, _05925_);
  nor (_02066_, _05646_, _02062_);
  or (_02068_, _02066_, rst);
  or (_02069_, _02068_, _02065_);
  or (_02501_, _02069_, _02060_);
  and (_02070_, _06878_, _06202_);
  nand (_02071_, _02070_, _05186_);
  and (_02072_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_02073_, _08283_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_02074_, _02073_, _08281_);
  and (_02075_, _02074_, _02070_);
  or (_02076_, _02075_, _02072_);
  and (_02077_, _02076_, _05647_);
  and (_02078_, _05649_, _05272_);
  nand (_02079_, _02078_, _06062_);
  or (_02080_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_02081_, _02080_, _05925_);
  and (_02082_, _02081_, _02079_);
  and (_02083_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_02084_, _02083_, rst);
  or (_02085_, _02084_, _02082_);
  or (_02502_, _02085_, _02077_);
  not (_02086_, _02078_);
  or (_02087_, _02086_, _05922_);
  or (_02088_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_02089_, _02088_, _05647_);
  and (_02090_, _02089_, _02087_);
  nand (_02091_, _02078_, _05604_);
  and (_02092_, _02088_, _05925_);
  and (_02093_, _02092_, _02091_);
  not (_02094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_02095_, _05646_, _02094_);
  or (_02096_, _02095_, rst);
  or (_02097_, _02096_, _02093_);
  or (_02504_, _02097_, _02090_);
  and (_02098_, _02016_, _10407_);
  nand (_02099_, _02098_, _05963_);
  or (_02100_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_02101_, _02100_, _05647_);
  and (_02102_, _02101_, _02099_);
  and (_02104_, _02022_, _06004_);
  not (_02105_, _02022_);
  and (_02106_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_02107_, _02106_, _02104_);
  and (_02108_, _02107_, _05925_);
  and (_02109_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_02110_, _02109_, rst);
  or (_02111_, _02110_, _02108_);
  or (_02517_, _02111_, _02102_);
  and (_02112_, _01257_, _10407_);
  nand (_02113_, _02112_, _05963_);
  or (_02114_, _02112_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_02115_, _02114_, _05647_);
  and (_02116_, _02115_, _02113_);
  and (_02117_, _01263_, _06004_);
  and (_02118_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_02119_, _02118_, _02117_);
  and (_02120_, _02119_, _05925_);
  and (_02121_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_02122_, _02121_, rst);
  or (_02123_, _02122_, _02120_);
  or (_02519_, _02123_, _02116_);
  and (_02124_, _02043_, _06207_);
  nand (_02125_, _02124_, _05963_);
  or (_02126_, _02124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_02127_, _02126_, _05647_);
  and (_02128_, _02127_, _02125_);
  nand (_02129_, _02049_, _06244_);
  or (_02130_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_02131_, _02130_, _05925_);
  and (_02132_, _02131_, _02129_);
  and (_02133_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_02134_, _02133_, rst);
  or (_02135_, _02134_, _02132_);
  or (_02522_, _02135_, _02128_);
  and (_02136_, _02043_, _05288_);
  nand (_02138_, _02136_, _05963_);
  or (_02139_, _02136_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_02140_, _02139_, _05647_);
  and (_02141_, _02140_, _02138_);
  nand (_02142_, _02049_, _06178_);
  or (_02143_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_02144_, _02143_, _05925_);
  and (_02145_, _02144_, _02142_);
  and (_02146_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_02147_, _02146_, rst);
  or (_02148_, _02147_, _02145_);
  or (_02523_, _02148_, _02141_);
  and (_02149_, _02043_, _08469_);
  nand (_02150_, _02149_, _05963_);
  or (_02151_, _02149_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_02152_, _02151_, _05647_);
  and (_02153_, _02152_, _02150_);
  not (_02154_, _02049_);
  or (_02155_, _02154_, _05522_);
  or (_02156_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_02157_, _02156_, _05925_);
  and (_02158_, _02157_, _02155_);
  and (_02159_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_02160_, _02159_, rst);
  or (_02161_, _02160_, _02158_);
  or (_02525_, _02161_, _02153_);
  nand (_02162_, _02070_, _08283_);
  and (_02163_, _02162_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02164_, _05287_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02165_, _02164_, _10356_);
  and (_02166_, _02165_, _02070_);
  or (_02167_, _02166_, _02163_);
  and (_02168_, _02167_, _05647_);
  nand (_02169_, _02078_, _05560_);
  or (_02170_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02171_, _02170_, _05925_);
  and (_02172_, _02171_, _02169_);
  and (_02173_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02174_, _02173_, rst);
  or (_02175_, _02174_, _02172_);
  or (_02526_, _02175_, _02168_);
  and (_02176_, _02070_, _10407_);
  nand (_02177_, _02176_, _05963_);
  or (_02178_, _02176_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_02179_, _02178_, _05647_);
  and (_02180_, _02179_, _02177_);
  or (_02181_, _02086_, _06004_);
  or (_02182_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_02183_, _02182_, _05925_);
  and (_02184_, _02183_, _02181_);
  and (_02185_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_02186_, _02185_, rst);
  or (_02187_, _02186_, _02184_);
  or (_02529_, _02187_, _02180_);
  and (_02188_, _01257_, _08469_);
  nand (_02189_, _02188_, _05963_);
  or (_02190_, _02188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_02191_, _02190_, _05647_);
  and (_02192_, _02191_, _02189_);
  and (_02193_, _01263_, _05522_);
  and (_02195_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_02196_, _02195_, _02193_);
  and (_02197_, _02196_, _05925_);
  and (_02198_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_02199_, _02198_, rst);
  or (_02200_, _02199_, _02197_);
  or (_02613_, _02200_, _02192_);
  and (_02201_, _01257_, _06032_);
  nand (_02202_, _02201_, _05963_);
  or (_02203_, _02201_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_02204_, _02203_, _05647_);
  and (_02205_, _02204_, _02202_);
  nor (_02206_, _01264_, _06062_);
  and (_02207_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_02208_, _02207_, _02206_);
  and (_02209_, _02208_, _05925_);
  and (_02210_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_02211_, _02210_, rst);
  or (_02212_, _02211_, _02209_);
  or (_02615_, _02212_, _02205_);
  and (_02213_, _01257_, _06620_);
  nand (_02214_, _02213_, _05963_);
  or (_02215_, _02213_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_02216_, _02215_, _05647_);
  and (_02217_, _02216_, _02214_);
  nor (_02218_, _01264_, _05560_);
  and (_02219_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02220_, _02219_, _02218_);
  and (_02222_, _02220_, _05925_);
  and (_02223_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02224_, _02223_, rst);
  or (_02225_, _02224_, _02222_);
  or (_02634_, _02225_, _02217_);
  or (_02226_, _02154_, _05922_);
  or (_02227_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_02228_, _02227_, _05647_);
  and (_02229_, _02228_, _02226_);
  nand (_02230_, _02049_, _05604_);
  and (_02231_, _02227_, _05925_);
  and (_02232_, _02231_, _02230_);
  not (_02233_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_02234_, _05646_, _02233_);
  or (_02235_, _02234_, rst);
  or (_02236_, _02235_, _02232_);
  or (_02635_, _02236_, _02229_);
  and (_02237_, _02016_, _06032_);
  nand (_02238_, _02237_, _05963_);
  or (_02239_, _02237_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_02240_, _02239_, _05647_);
  and (_02241_, _02240_, _02238_);
  nor (_02242_, _02105_, _06062_);
  and (_02243_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_02244_, _02243_, _02242_);
  and (_02245_, _02244_, _05925_);
  and (_02246_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_02247_, _02246_, rst);
  or (_02248_, _02247_, _02245_);
  or (_02638_, _02248_, _02241_);
  and (_02249_, _02016_, _06620_);
  nand (_02250_, _02249_, _05963_);
  or (_02251_, _02249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_02252_, _02251_, _05647_);
  and (_02253_, _02252_, _02250_);
  nor (_02254_, _02105_, _05560_);
  and (_02255_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_02256_, _02255_, _02254_);
  and (_02257_, _02256_, _05925_);
  and (_02258_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_02259_, _02258_, rst);
  or (_02260_, _02259_, _02257_);
  or (_02640_, _02260_, _02253_);
  and (_02261_, _05649_, _05276_);
  nand (_02262_, _02261_, _05963_);
  or (_02263_, _02261_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_02264_, _02263_, _05647_);
  and (_02265_, _02264_, _02262_);
  nand (_02266_, _02078_, _06178_);
  or (_02267_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_02268_, _02267_, _05925_);
  and (_02269_, _02268_, _02266_);
  and (_02270_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_02271_, _02270_, rst);
  or (_02272_, _02271_, _02269_);
  or (_02658_, _02272_, _02265_);
  and (_02273_, _02070_, _06207_);
  nand (_02274_, _02273_, _05963_);
  or (_02275_, _02273_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02276_, _02275_, _05647_);
  and (_02277_, _02276_, _02274_);
  nand (_02278_, _02078_, _06244_);
  or (_02279_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02280_, _02279_, _05925_);
  and (_02281_, _02280_, _02278_);
  and (_02282_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_02283_, _02282_, rst);
  or (_02284_, _02283_, _02281_);
  or (_02661_, _02284_, _02277_);
  and (_02285_, _02070_, _08469_);
  nand (_02286_, _02285_, _05963_);
  or (_02287_, _02285_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02288_, _02287_, _05647_);
  and (_02289_, _02288_, _02286_);
  or (_02290_, _02086_, _05522_);
  or (_02291_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02292_, _02291_, _05925_);
  and (_02293_, _02292_, _02290_);
  and (_02294_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_02295_, _02294_, rst);
  or (_02296_, _02295_, _02293_);
  or (_02664_, _02296_, _02289_);
  and (_02297_, _01257_, _05288_);
  nand (_02298_, _02297_, _05963_);
  or (_02299_, _02297_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_02300_, _02299_, _05647_);
  and (_02301_, _02300_, _02298_);
  nor (_02302_, _01264_, _06178_);
  and (_02303_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_02304_, _02303_, _02302_);
  and (_02305_, _02304_, _05925_);
  and (_02306_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_02307_, _02306_, rst);
  or (_02308_, _02307_, _02305_);
  or (_02666_, _02308_, _02301_);
  and (_02309_, _02043_, _10407_);
  nand (_02310_, _02309_, _05963_);
  or (_02311_, _02309_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_02312_, _02311_, _05647_);
  and (_02313_, _02312_, _02310_);
  or (_02314_, _02154_, _06004_);
  or (_02315_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_02316_, _02315_, _05925_);
  and (_02317_, _02316_, _02314_);
  and (_02318_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_02319_, _02318_, rst);
  or (_02320_, _02319_, _02317_);
  or (_02668_, _02320_, _02313_);
  and (_02321_, _02043_, _06032_);
  nand (_02322_, _02321_, _05963_);
  or (_02323_, _02321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02324_, _02323_, _05647_);
  and (_02325_, _02324_, _02322_);
  nand (_02326_, _02049_, _06062_);
  or (_02327_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02328_, _02327_, _05925_);
  and (_02329_, _02328_, _02326_);
  and (_02330_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_02331_, _02330_, rst);
  or (_02332_, _02331_, _02329_);
  or (_02670_, _02332_, _02325_);
  and (_02333_, _02016_, _05288_);
  nand (_02334_, _02333_, _05963_);
  or (_02335_, _02333_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_02336_, _02335_, _05647_);
  and (_02337_, _02336_, _02334_);
  nor (_02338_, _02105_, _06178_);
  and (_02339_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_02340_, _02339_, _02338_);
  and (_02341_, _02340_, _05925_);
  and (_02342_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_02343_, _02342_, rst);
  or (_02344_, _02343_, _02341_);
  or (_02672_, _02344_, _02337_);
  and (_02345_, _02016_, _06207_);
  nand (_02346_, _02345_, _05963_);
  or (_02347_, _02345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_02348_, _02347_, _05647_);
  and (_02349_, _02348_, _02346_);
  nor (_02350_, _02105_, _06244_);
  and (_02351_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_02352_, _02351_, _02350_);
  and (_02353_, _02352_, _05925_);
  and (_02354_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_02355_, _02354_, rst);
  or (_02356_, _02355_, _02353_);
  or (_02677_, _02356_, _02349_);
  and (_02357_, _02016_, _08469_);
  nand (_02358_, _02357_, _05963_);
  or (_02359_, _02357_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_02360_, _02359_, _05647_);
  and (_02361_, _02360_, _02358_);
  and (_02362_, _02022_, _05522_);
  and (_02363_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_02364_, _02363_, _02362_);
  and (_02365_, _02364_, _05925_);
  and (_02366_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_02367_, _02366_, rst);
  or (_02368_, _02367_, _02365_);
  or (_02679_, _02368_, _02361_);
  or (_02369_, _05277_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nand (_02370_, _06178_, _05277_);
  and (_02371_, _02370_, _02369_);
  or (_02372_, _02371_, _05572_);
  or (_02373_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_02374_, _02373_, _05141_);
  and (_02698_, _02374_, _02372_);
  and (_02375_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_02376_, pc_log_change, _13154_);
  or (_02377_, _02376_, _02375_);
  and (_02701_, _02377_, _05141_);
  or (_02378_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not (_02379_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_02380_, pc_log_change, _02379_);
  and (_02381_, _02380_, _05141_);
  and (_02705_, _02381_, _02378_);
  and (_02382_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  not (_02383_, pc_log_change);
  and (_02384_, _02383_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or (_02385_, _02384_, _02382_);
  and (_02710_, _02385_, _05141_);
  or (_02386_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nand (_02387_, pc_log_change, _01968_);
  and (_02388_, _02387_, _05141_);
  and (_02713_, _02388_, _02386_);
  and (_02389_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_02390_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_02391_, pc_log_change, _02390_);
  or (_02392_, _02391_, _02389_);
  and (_02715_, _02392_, _05141_);
  and (_02393_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_02395_, pc_log_change, _02379_);
  or (_02396_, _02395_, _02393_);
  and (_02723_, _02396_, _05141_);
  and (_02398_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_02399_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_02400_, pc_log_change, _02399_);
  or (_02401_, _02400_, _02398_);
  and (_02726_, _02401_, _05141_);
  and (_02402_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_02403_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_02404_, pc_log_change, _02403_);
  or (_02405_, _02404_, _02402_);
  and (_02730_, _02405_, _05141_);
  and (_02406_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_02407_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_02408_, pc_log_change, _02407_);
  or (_02409_, _02408_, _02406_);
  and (_02734_, _02409_, _05141_);
  and (_02410_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_02411_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_02412_, pc_log_change, _02411_);
  or (_02413_, _02412_, _02410_);
  and (_02738_, _02413_, _05141_);
  and (_02414_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_02415_, _02383_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or (_02416_, _02415_, _02414_);
  and (_02759_, _02416_, _05141_);
  and (_02417_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_02418_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_02419_, pc_log_change, _02418_);
  or (_02420_, _02419_, _02417_);
  and (_02760_, _02420_, _05141_);
  or (_02421_, _06363_, _07117_);
  or (_02422_, _06270_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_02423_, _02422_, _05141_);
  and (_02768_, _02423_, _02421_);
  and (_02424_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_02425_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_02426_, pc_log_change, _02425_);
  or (_02427_, _02426_, _02424_);
  and (_02771_, _02427_, _05141_);
  or (_02428_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nand (_02430_, pc_log_change, _02399_);
  and (_02432_, _02430_, _05141_);
  and (_02797_, _02432_, _02428_);
  or (_02433_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  not (_02434_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_02435_, pc_log_change, _02434_);
  and (_02436_, _02435_, _05141_);
  and (_02804_, _02436_, _02433_);
  and (_02437_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_02438_, pc_log_change, _02434_);
  or (_02439_, _02438_, _02437_);
  and (_02806_, _02439_, _05141_);
  and (_02440_, _02070_, _06008_);
  nand (_02441_, _02440_, _05963_);
  or (_02442_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_02443_, _02442_, _05647_);
  and (_02444_, _02443_, _02441_);
  nand (_02445_, _02078_, _05960_);
  or (_02446_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_02447_, _02446_, _05925_);
  and (_02448_, _02447_, _02445_);
  and (_02449_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_02450_, _02449_, rst);
  or (_02451_, _02450_, _02448_);
  or (_02824_, _02451_, _02444_);
  or (_02452_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand (_02453_, _07619_, _06462_);
  and (_02454_, _02453_, _05141_);
  and (_02828_, _02454_, _02452_);
  nor (_02455_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_02830_, _02455_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_02832_, _01280_, _05141_);
  and (_02456_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_02457_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  or (_02458_, _02457_, _02456_);
  and (_02840_, _02458_, _05141_);
  not (_02459_, _06678_);
  nor (_02460_, _02459_, _05960_);
  and (_02461_, _02459_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or (_02462_, _02461_, _02460_);
  and (_02863_, _02462_, _05141_);
  nor (_02463_, _05960_, _08484_);
  and (_02464_, _08484_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_02465_, _02464_, _05572_);
  or (_02466_, _02465_, _02463_);
  or (_02467_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_02468_, _02467_, _05141_);
  and (_02871_, _02468_, _02466_);
  nand (_02469_, _06707_, _05960_);
  or (_02470_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_02471_, _02470_, _05141_);
  and (_02876_, _02471_, _02469_);
  or (_02472_, _02459_, _05522_);
  or (_02473_, _06678_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_02474_, _02473_, _05141_);
  and (_02888_, _02474_, _02472_);
  and (_02475_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_02476_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or (_02897_, _02476_, _02475_);
  and (_02477_, _06154_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_02478_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_02479_, _02478_, _06156_);
  and (_02480_, _06180_, _06290_);
  or (_02481_, _02480_, _02479_);
  or (_02482_, _02481_, _02477_);
  and (_02915_, _02482_, _05141_);
  and (_02483_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_02484_, _13031_, _05617_);
  or (_02485_, _02484_, _02483_);
  and (_02925_, _02485_, _05141_);
  nor (_02486_, _06180_, _11869_);
  and (_02487_, _06180_, _13031_);
  or (_02488_, _02487_, _02486_);
  and (_02935_, _02488_, _05141_);
  nor (_02489_, _08294_, rxd_i);
  and (_02490_, _02489_, _06693_);
  nor (_02491_, _06693_, _06682_);
  not (_02492_, _06684_);
  and (_02494_, _08374_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand (_02496_, _02494_, _06683_);
  nand (_02497_, _02496_, _02492_);
  or (_02498_, _02497_, _02491_);
  or (_02500_, _02498_, _02490_);
  and (_02973_, _02500_, _06715_);
  and (_02503_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_02505_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_02987_, _02505_, _02503_);
  and (_02999_, _12483_, _05141_);
  and (_03006_, _12220_, _05141_);
  and (_03011_, _12351_, _05141_);
  or (_02506_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_02507_, _08447_, _08439_);
  or (_02508_, _02507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_02509_, _02508_, _11907_);
  or (_02510_, _02509_, _08463_);
  and (_02511_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_02512_, _02511_, _08457_);
  or (_02513_, _02512_, _02510_);
  nand (_02514_, _02513_, _02506_);
  nand (_02515_, _02514_, _11727_);
  nand (_02516_, _08471_, _05560_);
  or (_02518_, _11789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_02520_, _02518_, _05141_);
  and (_02521_, _02520_, _02516_);
  and (_03017_, _02521_, _02515_);
  and (_03021_, _12588_, _05141_);
  nor (_02524_, _11451_, rst);
  and (_03031_, _02524_, _12700_);
  and (_02527_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_02528_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_02530_, _02528_, _02527_);
  and (_03033_, _02530_, _05141_);
  nor (_03035_, _12770_, rst);
  or (_02531_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05143_);
  and (_02532_, _02531_, _06814_);
  or (_02533_, _11443_, _07105_);
  and (_02534_, _06995_, _06528_);
  and (_02535_, _06995_, _08339_);
  or (_02536_, _02535_, _02534_);
  or (_02537_, _02536_, _06530_);
  or (_02538_, _02537_, _02533_);
  and (_02539_, _06778_, _06540_);
  and (_02540_, _06771_, _06556_);
  nor (_02541_, _02540_, _02539_);
  nand (_02542_, _11434_, _02541_);
  or (_02543_, _02542_, _02538_);
  or (_02544_, _07110_, _06784_);
  or (_02545_, _12144_, _11430_);
  and (_02546_, _07041_, _06420_);
  or (_02547_, _02546_, _01379_);
  or (_02548_, _02547_, _02545_);
  or (_02549_, _02548_, _02544_);
  or (_02550_, _02549_, _02543_);
  and (_02551_, _06755_, _06565_);
  or (_02552_, _02551_, _06781_);
  and (_02553_, _11428_, _06417_);
  or (_02554_, _06570_, _06552_);
  and (_02555_, _02554_, _06420_);
  or (_02556_, _02555_, _02553_);
  or (_02557_, _02556_, _02552_);
  or (_02558_, _02557_, _01873_);
  or (_02559_, _02558_, _02550_);
  and (_02560_, _02559_, _06271_);
  or (_02561_, _02560_, _02532_);
  and (_03039_, _02561_, _05141_);
  and (_03045_, _12534_, _05141_);
  nor (_02562_, _06244_, _08484_);
  and (_02563_, _08484_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_02564_, _02563_, _05572_);
  or (_02565_, _02564_, _02562_);
  or (_02566_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_02567_, _02566_, _05141_);
  and (_03049_, _02567_, _02565_);
  and (_02568_, _08280_, _06008_);
  nand (_02569_, _02568_, _05963_);
  or (_02570_, _02568_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_02571_, _02570_, _08360_);
  and (_02572_, _02571_, _02569_);
  nor (_02573_, _08360_, _05960_);
  or (_02574_, _02573_, _02572_);
  and (_03067_, _02574_, _05141_);
  and (_02575_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02576_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_03074_, _02576_, _02575_);
  and (_02577_, _06293_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_02578_, _07053_, _06565_);
  and (_02579_, _02578_, _06544_);
  or (_02580_, _02579_, _02552_);
  and (_02581_, _11428_, _06420_);
  and (_02582_, _06574_, _06420_);
  and (_02583_, _02582_, _06450_);
  or (_02584_, _02583_, _02581_);
  or (_02585_, _02584_, _02580_);
  or (_02586_, _06774_, _06769_);
  or (_02587_, _01850_, _12138_);
  or (_02588_, _02587_, _02586_);
  or (_02589_, _02588_, _02585_);
  or (_02590_, _01861_, _06543_);
  or (_02591_, _02590_, _02589_);
  and (_02592_, _02591_, _06296_);
  or (_03080_, _02592_, _02577_);
  and (_03087_, _11633_, _06065_);
  and (_02593_, _06688_, _01794_);
  and (_02594_, _02593_, _06697_);
  or (_02595_, _02594_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not (_02596_, rxd_i);
  nand (_02597_, _02594_, _02596_);
  and (_02598_, _02597_, _05141_);
  and (_03090_, _02598_, _02595_);
  and (_02599_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_02600_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_03098_, _02600_, _02599_);
  and (_02601_, _02016_, _06008_);
  nand (_02602_, _02601_, _05963_);
  or (_02603_, _02601_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_02604_, _02603_, _05647_);
  and (_02605_, _02604_, _02602_);
  nor (_02606_, _02105_, _05960_);
  and (_02607_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_02608_, _02607_, _02606_);
  and (_02609_, _02608_, _05925_);
  and (_02610_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_02611_, _02610_, rst);
  or (_02612_, _02611_, _02609_);
  or (_03119_, _02612_, _02605_);
  and (_02614_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor (_02616_, _01802_, _08366_);
  not (_02617_, _06693_);
  or (_02618_, _02496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_02619_, _02618_, _06686_);
  and (_02620_, _02619_, _02617_);
  nor (_02621_, _02620_, _01797_);
  nand (_02622_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor (_02623_, _02622_, _02621_);
  or (_02624_, _02623_, _02616_);
  and (_02625_, _02624_, _06715_);
  or (_03123_, _02625_, _02614_);
  nand (_02626_, _08305_, _05960_);
  or (_02627_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_02628_, _02627_, _05141_);
  and (_03126_, _02628_, _02626_);
  and (_02629_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand (_02630_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor (_02631_, _02630_, _02621_);
  or (_02632_, _02631_, _02629_);
  and (_02633_, _02632_, _06715_);
  or (_03132_, _02633_, _02475_);
  and (_02636_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_02637_, _01797_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_02639_, _02637_, _02619_);
  or (_02641_, _06693_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_02642_, _02641_, _01790_);
  and (_02643_, _02642_, _02639_);
  or (_02644_, _02643_, _02636_);
  and (_02645_, _02644_, _06715_);
  or (_03134_, _02645_, _02503_);
  or (_02646_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_02647_, _02646_, _02621_);
  or (_02648_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_02649_, _02648_, _06715_);
  and (_02650_, _02649_, _02647_);
  or (_03136_, _02650_, _02575_);
  and (_02651_, _01898_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_02652_, _02651_, _01897_);
  and (_02653_, _02652_, _10346_);
  or (_02654_, _12689_, _05922_);
  nor (_02655_, _12690_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_02656_, _02655_, _10346_);
  and (_02657_, _02656_, _02654_);
  or (_02659_, _02657_, _10354_);
  or (_02662_, _02659_, _02653_);
  nand (_02663_, _10354_, _05960_);
  and (_02665_, _02663_, _05141_);
  and (_03139_, _02665_, _02662_);
  or (_02667_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_02669_, _02667_, _02621_);
  or (_02671_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02673_, _02671_, _06715_);
  and (_02674_, _02673_, _02669_);
  or (_03141_, _02674_, _02599_);
  and (_02675_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_02676_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_02678_, _02676_, _02621_);
  or (_02680_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_02681_, _02680_, _06715_);
  and (_02682_, _02681_, _02678_);
  or (_03143_, _02682_, _02675_);
  or (_02683_, _07080_, _07059_);
  and (_02684_, _02683_, _06271_);
  and (_02685_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02686_, _02685_, _07092_);
  or (_02687_, _02686_, _02684_);
  and (_03150_, _02687_, _05141_);
  and (_02688_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_02689_, _07044_, _06450_);
  or (_02690_, _02689_, _06979_);
  or (_02691_, _02690_, _07072_);
  or (_02692_, _02691_, _06820_);
  and (_02693_, _02692_, _06271_);
  or (_02694_, _02693_, _02688_);
  or (_02695_, _02694_, _07090_);
  and (_03152_, _02695_, _05141_);
  nand (_02696_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_02697_, _02696_, _08243_);
  and (_02699_, _08243_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_02700_, _02699_, _02697_);
  and (_03160_, _02700_, _05141_);
  or (_02702_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_02703_, _02702_, _02621_);
  or (_02704_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02706_, _02704_, _06715_);
  and (_02707_, _02706_, _02703_);
  or (_03168_, _02707_, _06714_);
  or (_02708_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_02709_, _02708_, _02621_);
  or (_02711_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_02712_, _02711_, _06715_);
  and (_02714_, _02712_, _02709_);
  or (_03170_, _02714_, _10324_);
  or (_02716_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_02717_, _02716_, _02621_);
  and (_02718_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_02719_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_02720_, _02719_, _06715_);
  or (_02721_, _02720_, _02718_);
  and (_03172_, _02721_, _02717_);
  or (_02722_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_02724_, _02722_, _02621_);
  and (_02725_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_02727_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  and (_02728_, _02727_, _06715_);
  or (_02729_, _02728_, _02725_);
  and (_03175_, _02729_, _02724_);
  or (_02731_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_02732_, _02731_, _02621_);
  and (_02733_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_02735_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  and (_02736_, _02735_, _06715_);
  or (_02737_, _02736_, _02733_);
  and (_03178_, _02737_, _02732_);
  nor (_02739_, _10407_, _05751_);
  or (_02740_, _02739_, _11665_);
  nand (_02741_, _02740_, _08163_);
  nor (_02742_, _07200_, _06842_);
  and (_02743_, _08171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_02744_, _02743_, _02742_);
  nand (_02745_, _02744_, _02741_);
  nand (_02746_, _02745_, _08158_);
  nand (_02747_, _07166_, _06836_);
  nand (_02748_, _02747_, _02746_);
  and (_03180_, _02748_, _05141_);
  and (_03183_, _12444_, _05141_);
  nor (_02749_, _06620_, _05464_);
  or (_02750_, _02749_, _10356_);
  nand (_02751_, _02750_, _08163_);
  nor (_02752_, _06842_, _06617_);
  and (_02753_, _08171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_02754_, _02753_, _02752_);
  and (_02755_, _02754_, _08158_);
  nand (_02756_, _02755_, _02751_);
  or (_02757_, _07378_, _08158_);
  and (_02758_, _02757_, _02756_);
  and (_03193_, _02758_, _05141_);
  or (_02761_, _11443_, _07070_);
  and (_02762_, _06755_, _06557_);
  or (_02763_, _02762_, _02582_);
  or (_02764_, _02763_, _02761_);
  or (_02765_, _07062_, _06818_);
  or (_02766_, _08334_, _02765_);
  or (_02767_, _02766_, _02764_);
  or (_02769_, _11429_, _02539_);
  or (_02770_, _02769_, _06819_);
  or (_02772_, _02770_, _02767_);
  or (_02773_, _12671_, _06530_);
  and (_02774_, _06828_, _06420_);
  or (_02775_, _02774_, _06795_);
  or (_02776_, _02775_, _02555_);
  or (_02777_, _02776_, _02773_);
  and (_02778_, _06755_, _06765_);
  and (_02779_, _06547_, _06420_);
  or (_02781_, _02779_, _02778_);
  or (_02782_, _02781_, _01864_);
  and (_02783_, _06828_, _06760_);
  and (_02784_, _06564_, _06544_);
  or (_02785_, _02784_, _02783_);
  or (_02786_, _02785_, _02782_);
  or (_02787_, _02786_, _02777_);
  or (_02788_, _02553_, _01870_);
  and (_02789_, _06755_, _06566_);
  or (_02790_, _01379_, _06793_);
  or (_02791_, _02790_, _02789_);
  or (_02792_, _02791_, _06541_);
  or (_02793_, _02792_, _02788_);
  or (_02794_, _02793_, _02787_);
  or (_02795_, _02794_, _02772_);
  and (_02796_, _02795_, _06271_);
  and (_02798_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_02799_, _06796_, _06821_);
  or (_02800_, _02799_, _06813_);
  or (_02801_, _02800_, _02798_);
  or (_02802_, _02801_, _02796_);
  and (_03195_, _02802_, _05141_);
  or (_02803_, _01851_, _07037_);
  and (_02805_, _02803_, _06531_);
  or (_02807_, _02769_, _08332_);
  or (_02808_, _02807_, _02805_);
  or (_02809_, _12139_, _08334_);
  or (_02810_, _02809_, _02781_);
  and (_02811_, _07069_, _06528_);
  or (_02812_, _11443_, _07042_);
  or (_02813_, _02812_, _02811_);
  and (_02814_, _06778_, _06528_);
  or (_02815_, _02814_, _06781_);
  or (_02816_, _07073_, _06793_);
  or (_02817_, _02816_, _02815_);
  or (_02818_, _02817_, _02813_);
  or (_02819_, _02818_, _02810_);
  or (_02820_, _02788_, _02777_);
  or (_02821_, _02820_, _02819_);
  or (_02822_, _02821_, _02808_);
  and (_02823_, _02822_, _06271_);
  and (_02825_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02826_, _02825_, _02800_);
  or (_02827_, _02826_, _02823_);
  and (_03198_, _02827_, _05141_);
  and (_02829_, _06154_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_02831_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_02833_, _02831_, _06156_);
  and (_02834_, _05605_, _05291_);
  or (_02835_, _02834_, _02833_);
  or (_02836_, _02835_, _02829_);
  and (_03300_, _02836_, _05141_);
  nor (_02837_, _07259_, _06842_);
  and (_02838_, _08171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_02839_, _02838_, _02837_);
  nor (_02841_, _02839_, _06836_);
  not (_02842_, _02841_);
  not (_02843_, _08163_);
  nor (_02844_, _08469_, _05339_);
  nor (_02845_, _02844_, _10380_);
  or (_02846_, _02845_, _02843_);
  nand (_02847_, _07229_, _06836_);
  and (_02848_, _02847_, _02846_);
  and (_02849_, _02848_, _02842_);
  nor (_03305_, _02849_, rst);
  and (_02850_, _06293_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_02851_, _06570_, _06566_);
  or (_02852_, _06767_, _06553_);
  or (_02853_, _02852_, _02851_);
  and (_02854_, _02853_, _06536_);
  or (_02855_, _02854_, _00612_);
  or (_02856_, _02789_, _11443_);
  or (_02857_, _02856_, _06989_);
  or (_02858_, _02857_, _07048_);
  or (_02859_, _02858_, _02544_);
  nand (_02860_, _06773_, _06566_);
  nand (_02861_, _02860_, _07051_);
  and (_02862_, _06570_, _06420_);
  or (_02864_, _02862_, _06756_);
  or (_02865_, _02539_, _06997_);
  or (_02866_, _02865_, _02864_);
  or (_02867_, _02866_, _02861_);
  or (_02868_, _02867_, _06985_);
  or (_02869_, _02868_, _02859_);
  or (_02870_, _02869_, _02855_);
  and (_02872_, _02870_, _06296_);
  or (_03316_, _02872_, _02850_);
  and (_02873_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_02874_, pc_log_change, _08551_);
  or (_02875_, _02874_, _02873_);
  and (_03319_, _02875_, _05141_);
  and (_02877_, _06283_, _05617_);
  and (_02878_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or (_02879_, _02878_, _02877_);
  and (_03372_, _02879_, _05141_);
  nand (_02880_, _08265_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or (_02881_, _08265_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_02882_, _02881_, _05141_);
  nand (_02883_, _02882_, _02880_);
  nor (_03519_, _02883_, _08243_);
  and (_02884_, _09451_, _08385_);
  and (_02885_, _08388_, _09438_);
  and (_02886_, _02885_, _09451_);
  nor (_02887_, _08388_, _00625_);
  or (_02889_, _02887_, _02886_);
  and (_02890_, _02889_, _08246_);
  nand (_02891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_02892_, _02891_, _08245_);
  or (_02893_, _02892_, _02890_);
  and (_02894_, _02893_, _09437_);
  or (_02895_, _02894_, _02884_);
  nand (_02896_, _02895_, _05141_);
  nor (_03523_, _02896_, _08243_);
  or (_02898_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nand (_02899_, pc_log_change, _02425_);
  and (_02900_, _02899_, _05141_);
  and (_03601_, _02900_, _02898_);
  and (_02901_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_02902_, _05617_, _05561_);
  or (_02903_, _02902_, _02901_);
  and (_03623_, _02903_, _05141_);
  or (_02904_, _12117_, _06996_);
  or (_02905_, _02904_, _11429_);
  or (_02906_, _02905_, _02553_);
  or (_02907_, _02906_, _01866_);
  or (_02908_, _02907_, _02792_);
  or (_02909_, _01870_, _06979_);
  and (_02910_, _02909_, _06449_);
  or (_02911_, _02762_, _13288_);
  or (_02912_, _02911_, _02862_);
  or (_02913_, _02912_, _08336_);
  or (_02914_, _01859_, _12131_);
  or (_02916_, _02914_, _02913_);
  or (_02917_, _02916_, _02910_);
  or (_02918_, _02917_, _02908_);
  and (_02919_, _02918_, _06296_);
  nor (_02920_, _06821_, rst);
  and (_02921_, _02920_, _06793_);
  and (_02922_, _06293_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_02923_, _02922_, _02921_);
  or (_03634_, _02923_, _02919_);
  nor (_02924_, _02773_, _01867_);
  nand (_02926_, _02924_, _11445_);
  or (_02927_, _06994_, _12927_);
  or (_02928_, _02927_, _12112_);
  or (_02929_, _02928_, _01381_);
  or (_02930_, _02929_, _02926_);
  and (_02931_, _06767_, _06535_);
  or (_02932_, _02931_, _02774_);
  or (_02933_, _02932_, _06780_);
  and (_02934_, _06773_, _06564_);
  or (_02936_, _02865_, _02781_);
  or (_02937_, _02936_, _02934_);
  or (_02938_, _02937_, _06764_);
  or (_02939_, _02938_, _02933_);
  or (_02940_, _02939_, _02930_);
  and (_02941_, _02940_, _06271_);
  and (_02942_, _06793_, _05143_);
  and (_02943_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02944_, _02943_, _02942_);
  or (_02945_, _02944_, _02941_);
  and (_03637_, _02945_, _05141_);
  and (_02946_, _12261_, _12372_);
  and (_02947_, _02946_, _01362_);
  and (_02948_, _02947_, _06838_);
  nor (_02949_, _02948_, _12697_);
  and (_02950_, _01288_, _06703_);
  or (_02951_, _02950_, _12610_);
  and (_02952_, _01303_, _06179_);
  and (_02953_, _01279_, _05561_);
  and (_02954_, _01309_, _06290_);
  or (_02955_, _02954_, _02953_);
  or (_02956_, _02955_, _02952_);
  or (_02957_, _02956_, _02951_);
  and (_02958_, _01288_, _05522_);
  or (_02959_, _02958_, _12608_);
  and (_02960_, _01309_, _13031_);
  and (_02961_, _01279_, _06283_);
  and (_02962_, _01303_, _06004_);
  or (_02963_, _02962_, _02961_);
  or (_02964_, _02963_, _02960_);
  or (_02965_, _02964_, _02959_);
  nand (_02966_, _02965_, _02957_);
  nor (_02967_, _02966_, _02949_);
  and (_02968_, _12372_, _01280_);
  nand (_02969_, _02968_, _12263_);
  or (_02970_, _02969_, _01419_);
  nand (_02971_, _02757_, _02756_);
  nand (_02972_, _02971_, _08415_);
  or (_02974_, _02971_, _08415_);
  nand (_02975_, _02974_, _02972_);
  nand (_02976_, _08187_, _08186_);
  nand (_02977_, _08509_, _02976_);
  or (_02978_, _08509_, _02976_);
  and (_02979_, _02978_, _02977_);
  nand (_02980_, _02979_, _02975_);
  or (_02981_, _02979_, _02975_);
  nand (_02982_, _02981_, _02980_);
  nand (_02983_, _02748_, _08177_);
  or (_02984_, _02748_, _08177_);
  and (_02985_, _02984_, _02983_);
  nand (_02986_, _02985_, _02982_);
  or (_02988_, _02985_, _02982_);
  and (_02989_, _02988_, _02986_);
  nand (_02990_, _02849_, _06977_);
  or (_02991_, _02849_, _06977_);
  and (_02992_, _02991_, _02990_);
  nand (_02993_, _02992_, _02989_);
  or (_02994_, _02992_, _02989_);
  and (_02995_, _02994_, _02993_);
  nand (_02996_, _02995_, _12608_);
  or (_02997_, _12608_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_02998_, _02997_, _01288_);
  and (_03000_, _02998_, _02996_);
  and (_03001_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_03002_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03003_, _03002_, _03001_);
  and (_03004_, _03003_, _12610_);
  and (_03005_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_03007_, _12608_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03008_, _03007_, _03005_);
  and (_03009_, _03008_, _01279_);
  and (_03010_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03012_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_03013_, _03012_, _03010_);
  and (_03014_, _03013_, _12608_);
  or (_03015_, _03014_, _03009_);
  or (_03016_, _03015_, _03004_);
  nor (_03018_, _03016_, _03000_);
  nor (_03019_, _03018_, _02970_);
  and (_03020_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_03022_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_03023_, _03022_, _03020_);
  and (_03024_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_03025_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_03026_, _03025_, _03024_);
  or (_03027_, _03026_, _03023_);
  and (_03028_, _03027_, _12608_);
  and (_03029_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_03030_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_03032_, _03030_, _03029_);
  and (_03034_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03036_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_03038_, _03036_, _03034_);
  or (_03040_, _03038_, _03032_);
  and (_03041_, _03040_, _12610_);
  nor (_03042_, _03041_, _03028_);
  nor (_03043_, _03042_, _01318_);
  and (_03044_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_03046_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_03047_, _03046_, _03044_);
  and (_03048_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_03050_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_03051_, _03050_, _03048_);
  or (_03052_, _03051_, _03047_);
  and (_03053_, _03052_, _12608_);
  and (_03054_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03055_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03056_, _03055_, _03054_);
  and (_03057_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_03058_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_03059_, _03058_, _03057_);
  or (_03060_, _03059_, _03056_);
  and (_03061_, _03060_, _12610_);
  or (_03062_, _03061_, _03053_);
  and (_03063_, _03062_, _01283_);
  and (_03064_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_03065_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_03066_, _03065_, _03064_);
  and (_03068_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_03069_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03070_, _03069_, _03068_);
  or (_03071_, _03070_, _03066_);
  and (_03072_, _03071_, _12608_);
  and (_03073_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_03075_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_03076_, _03075_, _03073_);
  and (_03077_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_03078_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_03079_, _03078_, _03077_);
  or (_03081_, _03079_, _03076_);
  and (_03082_, _03081_, _12610_);
  or (_03083_, _03082_, _03072_);
  and (_03084_, _03083_, _01343_);
  or (_03085_, _03084_, _03063_);
  or (_03086_, _03085_, _03043_);
  and (_03088_, _03086_, _12374_);
  or (_03089_, _01391_, p3_in[6]);
  or (_03091_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03092_, _03091_, _03089_);
  and (_03093_, _03092_, _01279_);
  or (_03094_, _03093_, _12608_);
  and (_03095_, _01402_, _01309_);
  or (_03096_, _01391_, p3_in[4]);
  or (_03097_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_03099_, _03097_, _03096_);
  and (_03100_, _03099_, _01288_);
  or (_03101_, _01391_, p3_in[5]);
  or (_03102_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03103_, _03102_, _03101_);
  and (_03104_, _03103_, _01303_);
  or (_03105_, _03104_, _03100_);
  or (_03106_, _03105_, _03095_);
  or (_03107_, _03106_, _03094_);
  nor (_03108_, _01391_, p3_in[0]);
  and (_03109_, _01391_, _02024_);
  nor (_03110_, _03109_, _03108_);
  and (_03111_, _03110_, _01288_);
  or (_03112_, _03111_, _12610_);
  or (_03113_, _01391_, p3_in[3]);
  or (_03114_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03115_, _03114_, _03113_);
  and (_03116_, _03115_, _01309_);
  or (_03117_, _01391_, p3_in[2]);
  or (_03118_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03120_, _03118_, _03117_);
  and (_03121_, _03120_, _01279_);
  or (_03122_, _01391_, p3_in[1]);
  or (_03124_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03125_, _03124_, _03122_);
  and (_03127_, _03125_, _01303_);
  or (_03128_, _03127_, _03121_);
  or (_03129_, _03128_, _03116_);
  or (_03130_, _03129_, _03112_);
  and (_03131_, _03130_, _03107_);
  or (_03133_, _03131_, _12261_);
  or (_03135_, _01317_, _12374_);
  or (_03137_, _01391_, p2_in[4]);
  or (_03138_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_03140_, _03138_, _03137_);
  and (_03142_, _03140_, _01288_);
  or (_03144_, _03142_, _12608_);
  or (_03145_, _01391_, p2_in[6]);
  or (_03146_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03147_, _03146_, _03145_);
  and (_03148_, _03147_, _01279_);
  or (_03149_, _01391_, p2_in[5]);
  or (_03151_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03153_, _03151_, _03149_);
  and (_03154_, _03153_, _01303_);
  and (_03155_, _01397_, _01309_);
  or (_03156_, _03155_, _03154_);
  or (_03157_, _03156_, _03148_);
  or (_03158_, _03157_, _03144_);
  or (_03159_, _01391_, p2_in[1]);
  or (_03161_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_03162_, _03161_, _03159_);
  and (_03163_, _03162_, _01303_);
  or (_03164_, _03163_, _12610_);
  or (_03165_, _01391_, p2_in[2]);
  or (_03166_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03167_, _03166_, _03165_);
  and (_03169_, _03167_, _01279_);
  nor (_03171_, _01391_, p2_in[0]);
  and (_03173_, _01391_, _02062_);
  nor (_03174_, _03173_, _03171_);
  and (_03176_, _03174_, _01288_);
  or (_03177_, _01391_, p2_in[3]);
  or (_03179_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03181_, _03179_, _03177_);
  and (_03182_, _03181_, _01309_);
  or (_03184_, _03182_, _03176_);
  or (_03185_, _03184_, _03169_);
  or (_03186_, _03185_, _03164_);
  and (_03187_, _03186_, _03158_);
  nor (_03188_, _03187_, _12263_);
  nor (_03189_, _03188_, _03135_);
  and (_03190_, _03189_, _03133_);
  or (_03191_, _01391_, p1_in[3]);
  or (_03192_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03194_, _03192_, _03191_);
  and (_03196_, _03194_, _01309_);
  or (_03197_, _03196_, _12610_);
  or (_03199_, _01391_, p1_in[1]);
  or (_03200_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03201_, _03200_, _03199_);
  and (_03202_, _03201_, _01303_);
  or (_03203_, _01391_, p1_in[2]);
  or (_03204_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03205_, _03204_, _03203_);
  and (_03206_, _03205_, _01279_);
  nor (_03207_, _01391_, p1_in[0]);
  and (_03208_, _01391_, _02233_);
  nor (_03209_, _03208_, _03207_);
  and (_03210_, _03209_, _01288_);
  or (_03211_, _03210_, _03206_);
  or (_03212_, _03211_, _03202_);
  or (_03213_, _03212_, _03197_);
  and (_03214_, _01343_, _12372_);
  and (_03215_, _01412_, _01309_);
  or (_03216_, _03215_, _12608_);
  or (_03217_, _01391_, p1_in[5]);
  or (_03218_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03219_, _03218_, _03217_);
  and (_03220_, _03219_, _01303_);
  or (_03221_, _01391_, p1_in[6]);
  or (_03222_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03223_, _03222_, _03221_);
  and (_03224_, _03223_, _01279_);
  or (_03225_, _01391_, p1_in[4]);
  or (_03226_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03227_, _03226_, _03225_);
  and (_03228_, _03227_, _01288_);
  or (_03229_, _03228_, _03224_);
  or (_03230_, _03229_, _03220_);
  or (_03231_, _03230_, _03216_);
  and (_03232_, _03231_, _03214_);
  and (_03233_, _03232_, _03213_);
  and (_03234_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_03235_, _03234_, _12608_);
  and (_03236_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03237_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_03238_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03239_, _03238_, _03237_);
  or (_03240_, _03239_, _03236_);
  or (_03241_, _03240_, _03235_);
  and (_03242_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03243_, _03242_, _12610_);
  and (_03244_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_03245_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_03246_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_03247_, _03246_, _03245_);
  or (_03248_, _03247_, _03244_);
  or (_03249_, _03248_, _03243_);
  and (_03250_, _03249_, _02947_);
  and (_03251_, _03250_, _03241_);
  or (_03252_, _03251_, _03233_);
  and (_03253_, _12261_, _12374_);
  nand (_03254_, _03253_, _01280_);
  or (_03255_, _03254_, _01419_);
  and (_03256_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_03257_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03258_, _03257_, _03256_);
  and (_03259_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_03260_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03261_, _03260_, _03259_);
  or (_03262_, _03261_, _03258_);
  and (_03263_, _03262_, _12608_);
  and (_03264_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03265_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_03266_, _03265_, _03264_);
  and (_03267_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03268_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_03269_, _03268_, _03267_);
  or (_03270_, _03269_, _03266_);
  and (_03271_, _03270_, _12610_);
  nor (_03272_, _03271_, _03263_);
  nor (_03273_, _03272_, _03255_);
  and (_03274_, _01322_, _12374_);
  and (_03275_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_03276_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03277_, _03276_, _03275_);
  and (_03278_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_03279_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_03280_, _03279_, _03278_);
  or (_03281_, _03280_, _03277_);
  and (_03282_, _03281_, _12608_);
  and (_03283_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_03284_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_03285_, _03284_, _03283_);
  and (_03286_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_03287_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_03288_, _03287_, _03286_);
  or (_03289_, _03288_, _03285_);
  and (_03290_, _03289_, _12610_);
  or (_03291_, _03290_, _03282_);
  and (_03292_, _03291_, _03274_);
  or (_03293_, _03292_, _03273_);
  or (_03294_, _03293_, _03252_);
  and (_03295_, _12615_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  nand (_03296_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_03297_, _03296_, _12610_);
  not (_03298_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_03299_, _12557_, _12502_);
  or (_03301_, _03299_, _03298_);
  nand (_03302_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_03303_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_03304_, _03303_, _03302_);
  and (_03306_, _03304_, _03301_);
  and (_03307_, _03306_, _03297_);
  and (_03308_, _12448_, _12313_);
  not (_03309_, _03308_);
  or (_03310_, _02969_, _03309_);
  nand (_03311_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_03312_, _03311_, _12608_);
  nand (_03313_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_03314_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_03315_, _03299_, _00747_);
  and (_03317_, _03315_, _03314_);
  and (_03318_, _03317_, _03313_);
  and (_03320_, _03318_, _03312_);
  or (_03321_, _03320_, _03310_);
  nor (_03322_, _03321_, _03307_);
  or (_03323_, _03322_, _03295_);
  or (_03324_, _01342_, _12374_);
  and (_03325_, _03310_, _03135_);
  and (_03326_, _03325_, _03324_);
  not (_03327_, _02970_);
  nor (_03328_, _03327_, _02947_);
  nand (_03329_, _01281_, _12374_);
  and (_03330_, _03329_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_03331_, _03330_, _03255_);
  and (_03332_, _03331_, _03328_);
  and (_03333_, _03332_, _03326_);
  or (_03334_, _01391_, p0_in[4]);
  or (_03335_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_03336_, _03335_, _03334_);
  and (_03337_, _03336_, _01288_);
  or (_03338_, _03337_, _12608_);
  or (_03339_, _01391_, p0_in[5]);
  or (_03340_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03341_, _03340_, _03339_);
  and (_03342_, _03341_, _01303_);
  and (_03343_, _01408_, _01309_);
  or (_03344_, _01391_, p0_in[6]);
  or (_03345_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03346_, _03345_, _03344_);
  and (_03347_, _03346_, _01279_);
  or (_03348_, _03347_, _03343_);
  or (_03349_, _03348_, _03342_);
  or (_03350_, _03349_, _03338_);
  and (_03351_, _01283_, _12372_);
  nor (_03352_, _01391_, p0_in[0]);
  and (_03353_, _01391_, _02094_);
  nor (_03354_, _03353_, _03352_);
  and (_03355_, _03354_, _01288_);
  or (_03356_, _03355_, _12610_);
  or (_03357_, _01391_, p0_in[2]);
  or (_03358_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_03359_, _03358_, _03357_);
  and (_03360_, _03359_, _01279_);
  or (_03361_, _01391_, p0_in[3]);
  or (_03362_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03363_, _03362_, _03361_);
  and (_03364_, _03363_, _01309_);
  or (_03365_, _01391_, p0_in[1]);
  or (_03366_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03367_, _03366_, _03365_);
  and (_03368_, _03367_, _01303_);
  or (_03369_, _03368_, _03364_);
  or (_03370_, _03369_, _03360_);
  or (_03371_, _03370_, _03356_);
  and (_03373_, _03371_, _03351_);
  and (_03374_, _03373_, _03350_);
  or (_03375_, _03374_, _03333_);
  or (_03376_, _03375_, _03323_);
  or (_03377_, _03376_, _03294_);
  or (_03378_, _03377_, _03190_);
  or (_03379_, _03378_, _03088_);
  or (_03380_, _03379_, _03019_);
  nand (_03381_, _03295_, _05963_);
  and (_03382_, _03381_, _02949_);
  and (_03383_, _03382_, _03380_);
  or (_03384_, _03383_, _02967_);
  and (_03643_, _03384_, _05141_);
  nand (_03385_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_03386_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_03387_, _03386_, _03385_);
  nand (_03388_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_03389_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_03390_, _03389_, _03388_);
  and (_03391_, _03390_, _03387_);
  nand (_03392_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_03393_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_03394_, _03393_, _03392_);
  nand (_03395_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_03396_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_03397_, _03396_, _03395_);
  and (_03398_, _03397_, _03394_);
  and (_03399_, _03398_, _03391_);
  nand (_03400_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_03401_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_03402_, _03401_, _03400_);
  nand (_03403_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand (_03404_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_03405_, _03404_, _03403_);
  and (_03406_, _03405_, _03402_);
  nand (_03407_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_03408_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_03409_, _03408_, _03407_);
  nand (_03410_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_03411_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_03412_, _03411_, _03410_);
  and (_03413_, _03412_, _03409_);
  and (_03414_, _03413_, _03406_);
  and (_03415_, _03414_, _03399_);
  nand (_03416_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_03417_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_03418_, _03417_, _03416_);
  nand (_03419_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not (_03420_, _12463_);
  nand (_03421_, _01368_, _03420_);
  and (_03422_, _03421_, _03419_);
  and (_03423_, _03422_, _03418_);
  nand (_03424_, _03110_, _01399_);
  nand (_03425_, _03174_, _01373_);
  and (_03426_, _03425_, _03424_);
  nand (_03427_, _03354_, _01405_);
  nand (_03428_, _03209_, _01413_);
  and (_03429_, _03428_, _03427_);
  and (_03430_, _03429_, _03426_);
  and (_03431_, _03430_, _03423_);
  not (_03432_, _01422_);
  or (_03433_, _02995_, _03432_);
  nand (_03434_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_03435_, _03434_, _03433_);
  and (_03436_, _03435_, _03431_);
  and (_03437_, _03436_, _03415_);
  nor (_03438_, _03437_, _01443_);
  not (_03439_, _01287_);
  nand (_03440_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_03441_, _03440_, _03439_);
  or (_03442_, _03441_, _03438_);
  nand (_03443_, _01287_, _07496_);
  and (_03444_, _03443_, _05141_);
  and (_03688_, _03444_, _03442_);
  or (_03445_, _06979_, _06772_);
  or (_03446_, _03445_, _06998_);
  or (_03447_, _03446_, _06763_);
  or (_03448_, _03447_, _00611_);
  or (_03449_, _01869_, _01380_);
  or (_03450_, _02934_, _02864_);
  or (_03451_, _03450_, _03449_);
  or (_03452_, _03451_, _02933_);
  or (_03453_, _03452_, _03448_);
  and (_03454_, _03453_, _06271_);
  and (_03455_, _06795_, _05143_);
  and (_03456_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_03457_, _03456_, _03455_);
  or (_03458_, _03457_, _03454_);
  and (_03698_, _03458_, _05141_);
  or (_03459_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_03460_, _01048_, rst);
  and (_03700_, _03460_, _03459_);
  or (_03461_, _01287_, rst);
  nor (_03709_, _03461_, _01441_);
  nand (_03462_, _02886_, _08245_);
  nand (_03463_, _03462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_03464_, _03463_, _02884_);
  or (_03465_, _03464_, _08243_);
  and (_03713_, _03465_, _05141_);
  and (_03466_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_03467_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_03468_, _03467_, _03466_);
  and (_03469_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_03470_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_03471_, _03470_, _03469_);
  or (_03472_, _03471_, _03468_);
  and (_03473_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_03474_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_03475_, _03474_, _03473_);
  and (_03476_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_03477_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_03478_, _03477_, _03476_);
  or (_03479_, _03478_, _03475_);
  or (_03480_, _03479_, _03472_);
  and (_03481_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_03482_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_03483_, _03482_, _03481_);
  and (_03484_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_03485_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_03486_, _03485_, _03484_);
  or (_03487_, _03486_, _03483_);
  and (_03488_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_03489_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03490_, _03489_, _03488_);
  and (_03491_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_03492_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_03493_, _03492_, _03491_);
  or (_03494_, _03493_, _03490_);
  or (_03495_, _03494_, _03487_);
  or (_03496_, _03495_, _03480_);
  and (_03497_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_03498_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_03499_, _03498_, _03497_);
  and (_03500_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not (_03501_, _12515_);
  and (_03502_, _01368_, _03501_);
  or (_03503_, _03502_, _03500_);
  or (_03504_, _03503_, _03499_);
  and (_03505_, _03162_, _01373_);
  and (_03506_, _03125_, _01399_);
  or (_03507_, _03506_, _03505_);
  and (_03508_, _03367_, _01405_);
  and (_03509_, _03201_, _01413_);
  or (_03510_, _03509_, _03508_);
  or (_03511_, _03510_, _03507_);
  or (_03512_, _03511_, _03504_);
  and (_03513_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03514_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03515_, _03514_, _03513_);
  or (_03516_, _03515_, _03512_);
  or (_03517_, _03516_, _03496_);
  and (_03518_, _03517_, _01441_);
  and (_03520_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or (_03521_, _03520_, _03518_);
  or (_03522_, _03521_, _01287_);
  nand (_03524_, _01287_, _07434_);
  and (_03525_, _03524_, _05141_);
  and (_03716_, _03525_, _03522_);
  and (_03526_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_03527_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_03528_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_03529_, _03528_, _03527_);
  and (_03530_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_03531_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_03532_, _03531_, _03530_);
  or (_03533_, _03532_, _03529_);
  and (_03534_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_03535_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_03536_, _03535_, _03534_);
  and (_03537_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_03538_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_03539_, _03538_, _03537_);
  or (_03540_, _03539_, _03536_);
  or (_03541_, _03540_, _03533_);
  and (_03542_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_03543_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_03544_, _03543_, _03542_);
  and (_03545_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_03546_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_03547_, _03546_, _03545_);
  or (_03548_, _03547_, _03544_);
  and (_03549_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_03550_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_03551_, _03550_, _03549_);
  and (_03552_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_03553_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03554_, _03553_, _03552_);
  or (_03555_, _03554_, _03551_);
  or (_03556_, _03555_, _03548_);
  or (_03557_, _03556_, _03541_);
  and (_03558_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_03559_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_03560_, _03559_, _03558_);
  and (_03561_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_03562_, _12569_);
  and (_03563_, _01368_, _03562_);
  or (_03564_, _03563_, _03561_);
  or (_03565_, _03564_, _03560_);
  and (_03566_, _03120_, _01399_);
  and (_03567_, _03167_, _01373_);
  or (_03568_, _03567_, _03566_);
  and (_03569_, _03359_, _01405_);
  and (_03570_, _03205_, _01413_);
  or (_03571_, _03570_, _03569_);
  or (_03572_, _03571_, _03568_);
  or (_03573_, _03572_, _03565_);
  and (_03574_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_03575_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03576_, _03575_, _03574_);
  or (_03577_, _03576_, _03573_);
  or (_03578_, _03577_, _03557_);
  and (_03579_, _03578_, _01441_);
  or (_03580_, _03579_, _01287_);
  or (_03581_, _03580_, _03526_);
  nand (_03582_, _01287_, _06617_);
  and (_03583_, _03582_, _05141_);
  and (_03728_, _03583_, _03581_);
  nor (_03584_, _01048_, _01047_);
  or (_03585_, _03584_, _01049_);
  and (_03586_, _01051_, _05141_);
  and (_03731_, _03586_, _03585_);
  or (_03587_, _02459_, _06004_);
  or (_03588_, _06678_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_03589_, _03588_, _05141_);
  and (_03745_, _03589_, _03587_);
  not (_03590_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_03591_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_03592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03593_, _05626_, _03592_);
  or (_03594_, _03593_, _08654_);
  nor (_03595_, _03594_, _03591_);
  nand (_03596_, _03595_, _03590_);
  nor (_03597_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor (_03598_, _03597_, _03595_);
  nand (_03599_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_03600_, _03599_, _03598_);
  and (_03602_, _03600_, _05141_);
  and (_03777_, _03602_, _03596_);
  and (_03604_, _06674_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nand (_03605_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_03606_, _03605_, _05278_);
  nor (_03607_, _02459_, _06062_);
  or (_03608_, _03607_, _03606_);
  or (_03609_, _03608_, _03604_);
  and (_03779_, _03609_, _05141_);
  and (_03610_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_03611_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  or (_03612_, _03611_, _03610_);
  and (_03795_, _03612_, _05141_);
  and (_03613_, _06293_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_03614_, _06774_, _06560_);
  or (_03615_, _03614_, _06990_);
  or (_03616_, _12671_, _02778_);
  or (_03617_, _03616_, _02862_);
  or (_03618_, _03617_, _07107_);
  or (_03619_, _03618_, _03615_);
  or (_03620_, _03619_, _02855_);
  and (_03621_, _03620_, _06296_);
  or (_03806_, _03621_, _03613_);
  and (_03816_, _03598_, _05141_);
  nor (_03624_, _02621_, _08366_);
  and (_03625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or (_03626_, _03625_, rxd_i);
  or (_03627_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_03628_, _03627_, _01801_);
  or (_03629_, _03628_, _01789_);
  and (_03630_, _03629_, _03626_);
  or (_03631_, _03630_, _03624_);
  nand (_03632_, _01789_, _02596_);
  and (_03633_, _03632_, _06715_);
  and (_03635_, _03633_, _03631_);
  and (_03636_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_03818_, _03636_, _03635_);
  nor (_03835_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  nand (_03638_, _06707_, _05604_);
  or (_03639_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_03640_, _03639_, _05141_);
  and (_03849_, _03640_, _03638_);
  or (_03641_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nand (_03642_, pc_log_change, _02403_);
  and (_03644_, _03642_, _05141_);
  and (_03854_, _03644_, _03641_);
  and (_03645_, _02043_, _06008_);
  nand (_03646_, _03645_, _05963_);
  or (_03647_, _03645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_03648_, _03647_, _05647_);
  and (_03649_, _03648_, _03646_);
  nand (_03650_, _02049_, _05960_);
  or (_03651_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_03652_, _03651_, _05925_);
  and (_03653_, _03652_, _03650_);
  and (_03654_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_03655_, _03654_, rst);
  or (_03656_, _03655_, _03653_);
  or (_03856_, _03656_, _03649_);
  or (_03657_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand (_03658_, _07619_, _06457_);
  and (_03659_, _03658_, _05141_);
  and (_03871_, _03659_, _03657_);
  and (_03660_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_03661_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  or (_03662_, _03661_, _03660_);
  and (_03876_, _03662_, _05141_);
  and (_03663_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_03664_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  or (_03665_, _03664_, _03663_);
  and (_03882_, _03665_, _05141_);
  or (_03666_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand (_03667_, _07619_, _06487_);
  and (_03668_, _03667_, _05141_);
  and (_03884_, _03668_, _03666_);
  and (_03669_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_03670_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or (_03671_, _03670_, _03669_);
  and (_03886_, _03671_, _05141_);
  and (_03672_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_03673_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or (_03674_, _03673_, _03672_);
  and (_03888_, _03674_, _05141_);
  and (_03675_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_03890_, _03675_, _02614_);
  and (_03676_, _06696_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_03677_, _03676_, _02594_);
  and (_03894_, _03677_, _05141_);
  and (_03678_, _01795_, _09587_);
  and (_03679_, _03678_, _06697_);
  nand (_03680_, _03679_, _02596_);
  or (_03681_, _03679_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_03682_, _03681_, _05141_);
  and (_03899_, _03682_, _03680_);
  and (_03683_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_03904_, _03683_, _02675_);
  nor (_03684_, _08440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor (_03685_, _03684_, _02507_);
  and (_03686_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_03687_, _03686_, _08457_);
  or (_03689_, _03687_, _03685_);
  and (_03690_, _03689_, _08464_);
  nand (_03691_, _08463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nand (_03692_, _03691_, _11727_);
  or (_03693_, _03692_, _03690_);
  nand (_03694_, _08471_, _06178_);
  or (_03695_, _11789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_03696_, _03695_, _05141_);
  and (_03697_, _03696_, _03694_);
  and (_03908_, _03697_, _03693_);
  nand (_03699_, _06707_, _06178_);
  or (_03701_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_03702_, _03701_, _05141_);
  and (_03910_, _03702_, _03699_);
  and (_03703_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_03704_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or (_03705_, _03704_, _03703_);
  and (_03912_, _03705_, _05141_);
  and (_03706_, _08078_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_03707_, _06244_, _08078_);
  or (_03708_, _03707_, _03706_);
  and (_03920_, _03708_, _05141_);
  nand (_03710_, _00698_, _06875_);
  or (_03711_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03712_, _03711_, _05925_);
  and (_03714_, _03712_, _03710_);
  nor (_03715_, _05646_, _03298_);
  and (_03717_, _00690_, _06008_);
  nand (_03718_, _03717_, _05963_);
  or (_03719_, _03717_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03720_, _03719_, _05647_);
  and (_03721_, _03720_, _03718_);
  or (_03722_, _03721_, _03715_);
  or (_03723_, _03722_, _03714_);
  and (_03923_, _03723_, _05141_);
  and (_03724_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_03725_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or (_03726_, _03725_, _03724_);
  and (_03933_, _03726_, _05141_);
  and (_03727_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_03729_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03730_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_03732_, _03730_, _03729_);
  and (_03733_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_03734_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_03735_, _03734_, _03733_);
  or (_03736_, _03735_, _03732_);
  and (_03737_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_03738_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_03739_, _03738_, _03737_);
  and (_03740_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_03741_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_03742_, _03741_, _03740_);
  or (_03743_, _03742_, _03739_);
  or (_03744_, _03743_, _03736_);
  and (_03746_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_03747_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_03748_, _03747_, _03746_);
  and (_03749_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_03750_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or (_03751_, _03750_, _03749_);
  or (_03752_, _03751_, _03748_);
  and (_03753_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_03754_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_03755_, _03754_, _03753_);
  and (_03756_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_03757_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_03758_, _03757_, _03756_);
  or (_03759_, _03758_, _03755_);
  or (_03760_, _03759_, _03752_);
  or (_03761_, _03760_, _03744_);
  and (_03762_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_03763_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_03764_, _03763_, _03762_);
  and (_03765_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_03766_, _01368_, _12257_);
  or (_03767_, _03766_, _03765_);
  or (_03768_, _03767_, _03764_);
  and (_03769_, _03099_, _01399_);
  and (_03770_, _03140_, _01373_);
  or (_03771_, _03770_, _03769_);
  and (_03772_, _03336_, _01405_);
  and (_03773_, _03227_, _01413_);
  or (_03774_, _03773_, _03772_);
  or (_03775_, _03774_, _03771_);
  or (_03776_, _03775_, _03768_);
  and (_03778_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_03780_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_03781_, _03780_, _03778_);
  or (_03782_, _03781_, _03776_);
  or (_03783_, _03782_, _03761_);
  and (_03784_, _03783_, _01441_);
  or (_03785_, _03784_, _01287_);
  or (_03786_, _03785_, _03727_);
  nand (_03787_, _01287_, _07259_);
  and (_03788_, _03787_, _05141_);
  and (_03979_, _03788_, _03786_);
  and (_03789_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_03790_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_03791_, _03790_, _03789_);
  and (_03792_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03793_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03794_, _03793_, _03792_);
  or (_03796_, _03794_, _03791_);
  and (_03797_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_03798_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_03799_, _03798_, _03797_);
  and (_03800_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_03801_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_03802_, _03801_, _03800_);
  or (_03803_, _03802_, _03799_);
  or (_03804_, _03803_, _03796_);
  and (_03805_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_03807_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_03808_, _03807_, _03805_);
  and (_03809_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_03810_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_03811_, _03810_, _03809_);
  or (_03812_, _03811_, _03808_);
  and (_03813_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_03814_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_03815_, _03814_, _03813_);
  and (_03817_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_03819_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or (_03820_, _03819_, _03817_);
  or (_03821_, _03820_, _03815_);
  or (_03822_, _03821_, _03812_);
  or (_03823_, _03822_, _03804_);
  and (_03824_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_03825_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_03826_, _03825_, _03824_);
  and (_03827_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_03828_, _01368_, _12325_);
  or (_03829_, _03828_, _03827_);
  or (_03830_, _03829_, _03826_);
  and (_03831_, _03181_, _01373_);
  and (_03832_, _03115_, _01399_);
  or (_03833_, _03832_, _03831_);
  and (_03834_, _03363_, _01405_);
  and (_03836_, _03194_, _01413_);
  or (_03837_, _03836_, _03834_);
  or (_03838_, _03837_, _03833_);
  or (_03839_, _03838_, _03830_);
  and (_03840_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_03841_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_03842_, _03841_, _03840_);
  or (_03843_, _03842_, _03839_);
  or (_03844_, _03843_, _03823_);
  and (_03845_, _03844_, _01441_);
  and (_03846_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or (_03847_, _03846_, _03845_);
  or (_03848_, _03847_, _01287_);
  nand (_03850_, _01287_, _07350_);
  and (_03851_, _03850_, _05141_);
  and (_03983_, _03851_, _03848_);
  and (_03852_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_03853_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_03855_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_03857_, _03855_, _03853_);
  and (_03858_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03859_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_03860_, _03859_, _03858_);
  or (_03861_, _03860_, _03857_);
  and (_03862_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_03863_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_03864_, _03863_, _03862_);
  and (_03865_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_03866_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_03867_, _03866_, _03865_);
  or (_03868_, _03867_, _03864_);
  or (_03869_, _03868_, _03861_);
  and (_03870_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_03872_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_03873_, _03872_, _03870_);
  and (_03874_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_03875_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_03877_, _03875_, _03874_);
  or (_03878_, _03877_, _03873_);
  and (_03879_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_03880_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_03881_, _03880_, _03879_);
  and (_03883_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_03885_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_03887_, _03885_, _03883_);
  or (_03889_, _03887_, _03881_);
  or (_03891_, _03889_, _03878_);
  or (_03892_, _03891_, _03869_);
  and (_03893_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_03895_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_03896_, _03895_, _03893_);
  and (_03897_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_03898_, _01368_, _12409_);
  or (_03900_, _03898_, _03897_);
  or (_03901_, _03900_, _03896_);
  and (_03902_, _03092_, _01399_);
  and (_03903_, _03147_, _01373_);
  or (_03905_, _03903_, _03902_);
  and (_03906_, _03346_, _01405_);
  and (_03907_, _03223_, _01413_);
  or (_03909_, _03907_, _03906_);
  or (_03911_, _03909_, _03905_);
  or (_03913_, _03911_, _03901_);
  and (_03914_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_03915_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_03916_, _03915_, _03914_);
  or (_03917_, _03916_, _03913_);
  or (_03918_, _03917_, _03892_);
  and (_03919_, _03918_, _01441_);
  or (_03921_, _03919_, _01287_);
  or (_03922_, _03921_, _03852_);
  or (_03924_, _03439_, _06669_);
  and (_03925_, _03924_, _05141_);
  and (_03989_, _03925_, _03922_);
  and (_03926_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_03927_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_03928_, _03927_, _03926_);
  and (_03929_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_03930_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_03931_, _03930_, _03929_);
  or (_03932_, _03931_, _03928_);
  and (_03934_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_03935_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03937_, _03935_, _03934_);
  and (_03938_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_03939_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_03940_, _03939_, _03938_);
  or (_03941_, _03940_, _03937_);
  or (_03942_, _03941_, _03932_);
  and (_03943_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_03944_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_03945_, _03944_, _03943_);
  and (_03946_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_03947_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_03948_, _03947_, _03946_);
  or (_03949_, _03948_, _03945_);
  and (_03950_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_03951_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_03952_, _03951_, _03950_);
  and (_03953_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_03954_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_03955_, _03954_, _03953_);
  or (_03956_, _03955_, _03952_);
  or (_03957_, _03956_, _03949_);
  or (_03958_, _03957_, _03942_);
  and (_03959_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_03960_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_03961_, _03960_, _03959_);
  and (_03962_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_03963_, _12304_);
  and (_03964_, _01368_, _03963_);
  or (_03965_, _03964_, _03962_);
  or (_03966_, _03965_, _03961_);
  and (_03967_, _03103_, _01399_);
  and (_03968_, _03153_, _01373_);
  or (_03969_, _03968_, _03967_);
  and (_03970_, _03341_, _01405_);
  and (_03971_, _03219_, _01413_);
  or (_03972_, _03971_, _03970_);
  or (_03973_, _03972_, _03969_);
  or (_03974_, _03973_, _03966_);
  and (_03975_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_03976_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_03977_, _03976_, _03975_);
  or (_03978_, _03977_, _03974_);
  or (_03980_, _03978_, _03958_);
  and (_03981_, _03980_, _01441_);
  and (_03982_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or (_03984_, _03982_, _03981_);
  or (_03985_, _03984_, _01287_);
  nand (_03986_, _01287_, _07200_);
  and (_03987_, _03986_, _05141_);
  and (_03993_, _03987_, _03985_);
  nor (_03988_, _05960_, _08078_);
  and (_03990_, _08078_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_03991_, _03990_, _03988_);
  and (_03995_, _03991_, _05141_);
  and (_03992_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_03994_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or (_03996_, _03994_, _03992_);
  and (_03997_, _03996_, _05141_);
  and (_03999_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_04000_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or (_04001_, _04000_, _03999_);
  and (_03998_, _04001_, _05141_);
  and (_04002_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_04003_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or (_04004_, _04003_, _04002_);
  and (_04059_, _04004_, _05141_);
  and (_04005_, _13031_, _05523_);
  and (_04006_, _01964_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or (_04007_, _04006_, _04005_);
  and (_04083_, _04007_, _05141_);
  and (_04008_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_04009_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04010_, pc_log_change, _04009_);
  or (_04011_, _04010_, _04008_);
  and (_04103_, _04011_, _05141_);
  and (_04012_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_04013_, _04012_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04014_, _04013_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_04015_, _04014_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_04016_, _04015_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_04017_, _04016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_04018_, _04017_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_04019_, _04018_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_04020_, _04019_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_04021_, _04020_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_04022_, _04021_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_04023_, _04022_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_04024_, _04022_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_04025_, _04024_, _04023_);
  nor (_04026_, _04025_, cy_reg);
  and (_04027_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_04028_, _04027_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  not (_04029_, _04028_);
  or (_04030_, _04027_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04031_, _04030_, _04029_);
  not (_04032_, _04031_);
  or (_04033_, _04028_, _07607_);
  nand (_04034_, _04028_, _07607_);
  and (_04035_, _04034_, _04033_);
  nand (_04036_, _04035_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_04038_, _04035_, _08192_);
  nand (_04039_, _04038_, _04036_);
  nand (_04040_, _04039_, _04032_);
  not (_04041_, _04035_);
  or (_04042_, _04041_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_04043_, _04035_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_04044_, _04043_, _04031_);
  nand (_04045_, _04044_, _04042_);
  nand (_04046_, _04045_, _04040_);
  nand (_04047_, _04046_, _04027_);
  nor (_04048_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nand (_04049_, _04035_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_04050_, _04035_, _07661_);
  nand (_04051_, _04050_, _04049_);
  nand (_04052_, _04051_, _04032_);
  or (_04053_, _04041_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_04054_, _04035_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_04055_, _04054_, _04031_);
  nand (_04056_, _04055_, _04053_);
  nand (_04057_, _04056_, _04052_);
  nand (_04058_, _04057_, _04048_);
  and (_04060_, _04058_, _04047_);
  and (_04061_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _02390_);
  nand (_04062_, _04035_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_04063_, _04035_, _07691_);
  and (_04064_, _04063_, _04062_);
  or (_04065_, _04064_, _04032_);
  or (_04066_, _04035_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_04067_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_04068_, _04035_, _04067_);
  and (_04069_, _04068_, _04066_);
  nand (_04070_, _04069_, _04032_);
  nand (_04071_, _04070_, _04065_);
  nand (_04072_, _04071_, _04061_);
  and (_04073_, _04009_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nand (_04074_, _04035_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_04075_, _04035_, _08257_);
  nand (_04076_, _04075_, _04074_);
  nand (_04077_, _04076_, _04032_);
  or (_04078_, _04035_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand (_04079_, _04035_, _07652_);
  and (_04080_, _04079_, _04031_);
  nand (_04081_, _04080_, _04078_);
  nand (_04082_, _04081_, _04077_);
  nand (_04084_, _04082_, _04073_);
  and (_04085_, _04084_, _04072_);
  and (_04086_, _04085_, _04060_);
  and (_04087_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_04088_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor (_04089_, _04088_, _04087_);
  and (_04090_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_04091_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_04092_, _04091_, _04090_);
  and (_04093_, _04092_, _04089_);
  and (_04094_, _04093_, _04032_);
  and (_04095_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_04096_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nor (_04097_, _04096_, _04095_);
  and (_04098_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_04099_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_04100_, _04099_, _04098_);
  and (_04101_, _04100_, _04097_);
  and (_04102_, _04101_, _04031_);
  or (_04104_, _04102_, _04041_);
  nor (_04105_, _04104_, _04094_);
  and (_04106_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_04107_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor (_04108_, _04107_, _04106_);
  and (_04109_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_04110_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_04111_, _04110_, _04109_);
  and (_04112_, _04111_, _04108_);
  and (_04113_, _04112_, _04032_);
  and (_04114_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_04115_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nor (_04116_, _04115_, _04114_);
  and (_04117_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_04118_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_04119_, _04118_, _04117_);
  and (_04120_, _04119_, _04116_);
  and (_04121_, _04120_, _04031_);
  or (_04122_, _04121_, _04035_);
  nor (_04123_, _04122_, _04113_);
  nor (_04124_, _04123_, _04105_);
  nor (_04125_, _04124_, _04086_);
  and (_04126_, _04125_, _04025_);
  nor (_04127_, _04125_, _04025_);
  nor (_04128_, _04127_, _04126_);
  not (_04129_, _04128_);
  nor (_04130_, _04021_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_04131_, _04130_, _04022_);
  and (_04132_, _04131_, _04125_);
  not (_04133_, _04132_);
  nor (_04134_, _04020_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_04135_, _04134_, _04021_);
  and (_04136_, _04135_, _04125_);
  nor (_04137_, _04019_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_04138_, _04137_, _04020_);
  and (_04139_, _04138_, _04125_);
  nor (_04140_, _04139_, _04136_);
  nor (_04142_, _04135_, _04125_);
  nor (_04143_, _04142_, _04136_);
  not (_04144_, _04143_);
  nor (_04145_, _04138_, _04125_);
  nor (_04146_, _04145_, _04139_);
  nor (_04147_, _04018_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_04148_, _04147_, _04019_);
  and (_04149_, _04148_, _04125_);
  nor (_04150_, _04017_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_04151_, _04150_, _04018_);
  and (_04152_, _04151_, _04125_);
  nor (_04153_, _04152_, _04149_);
  nor (_04154_, _04148_, _04125_);
  nor (_04155_, _04154_, _04149_);
  not (_04156_, _04155_);
  nor (_04157_, _04016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_04158_, _04157_, _04017_);
  and (_04159_, _04158_, _04125_);
  nor (_04160_, _04158_, _04125_);
  nor (_04161_, _04015_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_04162_, _04161_, _04016_);
  and (_04163_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_04164_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_04165_, _04164_, _04163_);
  and (_04166_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_04167_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_04168_, _04167_, _04166_);
  and (_04169_, _04168_, _04165_);
  nor (_04170_, _04169_, _04031_);
  and (_04171_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_04172_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_04173_, _04172_, _04171_);
  and (_04174_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_04175_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_04176_, _04175_, _04174_);
  and (_04177_, _04176_, _04173_);
  nor (_04178_, _04177_, _04032_);
  or (_04179_, _04178_, _04170_);
  and (_04180_, _04179_, _04035_);
  and (_04181_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_04182_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_04183_, _04182_, _04181_);
  and (_04184_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_04185_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_04186_, _04185_, _04184_);
  and (_04187_, _04186_, _04183_);
  and (_04188_, _04187_, _04032_);
  and (_04189_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_04190_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_04191_, _04190_, _04189_);
  and (_04192_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_04193_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_04194_, _04193_, _04192_);
  and (_04195_, _04194_, _04191_);
  and (_04196_, _04195_, _04031_);
  or (_04197_, _04196_, _04035_);
  nor (_04198_, _04197_, _04188_);
  nor (_04199_, _04198_, _04180_);
  nor (_04200_, _04199_, _04086_);
  and (_04201_, _04200_, _04162_);
  nor (_04202_, _04200_, _04162_);
  nor (_04203_, _04202_, _04201_);
  and (_04204_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_04205_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_04206_, _04205_, _04204_);
  and (_04207_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_04208_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_04209_, _04208_, _04207_);
  and (_04210_, _04209_, _04206_);
  nor (_04211_, _04210_, _04031_);
  and (_04212_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_04213_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_04214_, _04213_, _04212_);
  and (_04215_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_04216_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_04217_, _04216_, _04215_);
  and (_04218_, _04217_, _04214_);
  nor (_04219_, _04218_, _04032_);
  or (_04220_, _04219_, _04211_);
  and (_04221_, _04220_, _04035_);
  and (_04222_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_04223_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_04224_, _04223_, _04222_);
  and (_04225_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_04226_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_04227_, _04226_, _04225_);
  and (_04228_, _04227_, _04224_);
  nor (_04229_, _04228_, _04031_);
  and (_04230_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_04231_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_04232_, _04231_, _04230_);
  and (_04233_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_04234_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_04235_, _04234_, _04233_);
  and (_04236_, _04235_, _04232_);
  nor (_04237_, _04236_, _04032_);
  or (_04238_, _04237_, _04229_);
  and (_04239_, _04238_, _04041_);
  nor (_04240_, _04239_, _04221_);
  nor (_04241_, _04240_, _04086_);
  nor (_04242_, _04014_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_04243_, _04242_, _04015_);
  and (_04244_, _04243_, _04241_);
  nor (_04245_, _04243_, _04241_);
  nor (_04246_, _04245_, _04244_);
  nor (_04247_, _04013_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_04248_, _04247_, _04014_);
  and (_04249_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_04250_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_04251_, _04250_, _04249_);
  and (_04252_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_04253_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_04254_, _04253_, _04252_);
  and (_04255_, _04254_, _04251_);
  and (_04256_, _04255_, _04032_);
  and (_04257_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_04258_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_04259_, _04258_, _04257_);
  and (_04260_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_04261_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_04262_, _04261_, _04260_);
  and (_04263_, _04262_, _04259_);
  and (_04264_, _04263_, _04031_);
  or (_04265_, _04264_, _04041_);
  nor (_04266_, _04265_, _04256_);
  and (_04267_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_04268_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_04269_, _04268_, _04267_);
  and (_04270_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_04271_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_04272_, _04271_, _04270_);
  and (_04273_, _04272_, _04269_);
  nor (_04274_, _04273_, _04031_);
  and (_04275_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_04276_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_04277_, _04276_, _04275_);
  and (_04278_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_04279_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_04280_, _04279_, _04278_);
  and (_04281_, _04280_, _04277_);
  nor (_04282_, _04281_, _04032_);
  or (_04283_, _04282_, _04274_);
  and (_04284_, _04283_, _04041_);
  nor (_04285_, _04284_, _04266_);
  nor (_04286_, _04285_, _04086_);
  and (_04287_, _04286_, _04248_);
  nor (_04288_, _04012_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04289_, _04288_, _04013_);
  and (_04290_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_04291_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_04292_, _04291_, _04290_);
  and (_04293_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_04294_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_04295_, _04294_, _04293_);
  and (_04296_, _04295_, _04292_);
  and (_04297_, _04296_, _04032_);
  and (_04298_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_04299_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_04300_, _04299_, _04298_);
  and (_04301_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_04302_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_04303_, _04302_, _04301_);
  and (_04304_, _04303_, _04300_);
  and (_04305_, _04304_, _04031_);
  or (_04306_, _04305_, _04041_);
  nor (_04307_, _04306_, _04297_);
  and (_04308_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_04309_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_04310_, _04309_, _04308_);
  and (_04311_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_04312_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_04313_, _04312_, _04311_);
  and (_04314_, _04313_, _04310_);
  nor (_04315_, _04314_, _04031_);
  and (_04316_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_04317_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_04318_, _04317_, _04316_);
  and (_04319_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_04320_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_04321_, _04320_, _04319_);
  and (_04322_, _04321_, _04318_);
  nor (_04323_, _04322_, _04032_);
  or (_04324_, _04323_, _04315_);
  and (_04325_, _04324_, _04041_);
  nor (_04326_, _04325_, _04307_);
  nor (_04327_, _04326_, _04086_);
  and (_04328_, _04327_, _04289_);
  not (_04329_, _04328_);
  nor (_04330_, _04327_, _04289_);
  and (_04331_, _02418_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_04332_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _02390_);
  nor (_04333_, _04332_, _04331_);
  not (_04334_, _04333_);
  not (_04335_, _04086_);
  and (_04336_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_04337_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_04338_, _04337_, _04336_);
  and (_04339_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_04340_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_04341_, _04340_, _04339_);
  and (_04342_, _04341_, _04338_);
  and (_04343_, _04342_, _04032_);
  and (_04344_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_04345_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_04346_, _04345_, _04344_);
  and (_04347_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_04348_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_04349_, _04348_, _04347_);
  and (_04350_, _04349_, _04346_);
  nand (_04351_, _04350_, _04031_);
  nand (_04352_, _04351_, _04041_);
  or (_04353_, _04352_, _04343_);
  and (_04354_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_04355_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_04356_, _04355_, _04354_);
  and (_04357_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_04358_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_04359_, _04358_, _04357_);
  and (_04360_, _04359_, _04356_);
  and (_04361_, _04360_, _04031_);
  and (_04362_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_04363_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_04364_, _04363_, _04362_);
  and (_04365_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_04366_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_04367_, _04366_, _04365_);
  and (_04368_, _04367_, _04364_);
  nand (_04369_, _04368_, _04032_);
  nand (_04370_, _04369_, _04035_);
  or (_04371_, _04370_, _04361_);
  nand (_04372_, _04371_, _04353_);
  and (_04373_, _04372_, _04335_);
  nand (_04374_, _04373_, _04334_);
  nand (_04375_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nand (_04376_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_04377_, _04376_, _04375_);
  nand (_04378_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nand (_04379_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_04380_, _04379_, _04378_);
  and (_04381_, _04380_, _04377_);
  nand (_04382_, _04381_, _04032_);
  nand (_04383_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nand (_04384_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_04385_, _04384_, _04383_);
  nand (_04386_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nand (_04387_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_04388_, _04387_, _04386_);
  and (_04389_, _04388_, _04385_);
  nand (_04390_, _04389_, _04031_);
  and (_04391_, _04390_, _04041_);
  nand (_04392_, _04391_, _04382_);
  nand (_04393_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nand (_04394_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_04395_, _04394_, _04393_);
  nand (_04396_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nand (_04397_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_04398_, _04397_, _04396_);
  and (_04399_, _04398_, _04395_);
  nand (_04400_, _04399_, _04032_);
  nand (_04401_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nand (_04402_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_04403_, _04402_, _04401_);
  nand (_04404_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nand (_04405_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_04406_, _04405_, _04404_);
  and (_04407_, _04406_, _04403_);
  nand (_04408_, _04407_, _04031_);
  and (_04409_, _04408_, _04035_);
  nand (_04410_, _04409_, _04400_);
  nand (_04411_, _04410_, _04392_);
  and (_04412_, _04411_, _04335_);
  nand (_04413_, _04412_, _02390_);
  nand (_04414_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand (_04415_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_04416_, _04415_, _04414_);
  and (_04417_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_04418_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_04419_, _04418_, _04417_);
  and (_04420_, _04419_, _04416_);
  nand (_04421_, _04420_, _04032_);
  nand (_04422_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nand (_04423_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_04424_, _04423_, _04422_);
  nand (_04425_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand (_04426_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_04427_, _04426_, _04425_);
  and (_04428_, _04427_, _04424_);
  nand (_04429_, _04428_, _04031_);
  and (_04430_, _04429_, _04035_);
  nand (_04431_, _04430_, _04421_);
  and (_04432_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_04433_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_04434_, _04433_, _04432_);
  and (_04435_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_04436_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_04437_, _04436_, _04435_);
  and (_04438_, _04437_, _04434_);
  nand (_04439_, _04438_, _04032_);
  nand (_04440_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nand (_04441_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_04442_, _04441_, _04440_);
  nand (_04443_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nand (_04444_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_04445_, _04444_, _04443_);
  and (_04446_, _04445_, _04442_);
  nand (_04447_, _04446_, _04031_);
  and (_04448_, _04447_, _04041_);
  nand (_04449_, _04448_, _04439_);
  and (_04450_, _04449_, _04431_);
  or (_04451_, _04450_, _04086_);
  or (_04452_, _04451_, _04009_);
  or (_04453_, _04412_, _02390_);
  nand (_04454_, _04453_, _04413_);
  or (_04455_, _04454_, _04452_);
  and (_04456_, _04455_, _04413_);
  not (_04457_, _04456_);
  or (_04458_, _04373_, _04334_);
  and (_04459_, _04458_, _04374_);
  nand (_04460_, _04459_, _04457_);
  and (_04461_, _04460_, _04374_);
  or (_04462_, _04461_, _04330_);
  nand (_04463_, _04462_, _04329_);
  nor (_04464_, _04286_, _04248_);
  nor (_04465_, _04464_, _04287_);
  and (_04466_, _04465_, _04463_);
  or (_04467_, _04466_, _04287_);
  and (_04468_, _04467_, _04246_);
  or (_04469_, _04468_, _04244_);
  and (_04470_, _04469_, _04203_);
  nor (_04471_, _04470_, _04201_);
  nor (_04472_, _04471_, _04160_);
  or (_04473_, _04472_, _04159_);
  nor (_04474_, _04151_, _04125_);
  nor (_04475_, _04474_, _04152_);
  nand (_04476_, _04475_, _04473_);
  or (_04477_, _04476_, _04156_);
  nand (_04478_, _04477_, _04153_);
  nand (_04479_, _04478_, _04146_);
  or (_04480_, _04479_, _04144_);
  nand (_04481_, _04480_, _04140_);
  nor (_04482_, _04131_, _04125_);
  nor (_04483_, _04482_, _04132_);
  nand (_04484_, _04483_, _04481_);
  nand (_04485_, _04484_, _04133_);
  nor (_04486_, _04485_, _04129_);
  and (_04487_, _04485_, _04129_);
  nor (_04488_, _04487_, _04486_);
  and (_04489_, _04488_, cy_reg);
  nor (_04490_, _04489_, _04026_);
  nor (_04491_, _04490_, _01810_);
  and (_04492_, _04490_, _01810_);
  nor (_04493_, _04135_, cy_reg);
  and (_04494_, _04478_, _04146_);
  nor (_04495_, _04494_, _04139_);
  nand (_04496_, _04495_, _04144_);
  or (_04497_, _04495_, _04144_);
  nand (_04498_, _04497_, _04496_);
  and (_04499_, _04498_, cy_reg);
  or (_04500_, _04499_, _04493_);
  nor (_04501_, _04500_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_04502_, _04500_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not (_04503_, cy_reg);
  and (_04504_, _04148_, _04503_);
  and (_04505_, _04475_, _04473_);
  nor (_04506_, _04505_, _04152_);
  nand (_04507_, _04506_, _04155_);
  or (_04508_, _04506_, _04155_);
  nand (_04509_, _04508_, _04507_);
  and (_04510_, _04509_, cy_reg);
  nor (_04511_, _04510_, _04504_);
  nor (_04512_, _04511_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_04513_, _04511_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_04514_, _04151_, _04503_);
  or (_04515_, _04475_, _04473_);
  and (_04516_, _04515_, _04476_);
  and (_04517_, _04516_, cy_reg);
  nor (_04518_, _04517_, _04514_);
  nor (_04519_, _04518_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_04520_, _04518_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_04521_, _04158_, cy_reg);
  nor (_04522_, _04159_, _04160_);
  and (_04523_, _04522_, _04471_);
  nor (_04524_, _04522_, _04471_);
  nor (_04525_, _04524_, _04523_);
  and (_04526_, _04525_, cy_reg);
  nor (_04527_, _04526_, _04521_);
  nor (_04528_, _04527_, _02403_);
  and (_04529_, _04527_, _02403_);
  and (_04530_, _04162_, _04503_);
  nor (_04531_, _04469_, _04203_);
  nor (_04532_, _04531_, _04470_);
  and (_04533_, _04532_, cy_reg);
  or (_04534_, _04533_, _04530_);
  nor (_04535_, _04534_, _08551_);
  and (_04536_, _04534_, _08551_);
  and (_04537_, _04243_, _04503_);
  nor (_04538_, _04467_, _04246_);
  nor (_04539_, _04538_, _04468_);
  and (_04540_, _04539_, cy_reg);
  or (_04541_, _04540_, _04537_);
  nor (_04542_, _04541_, _01968_);
  and (_04543_, _04541_, _01968_);
  and (_04544_, _04248_, _04503_);
  nor (_04545_, _04465_, _04463_);
  nor (_04546_, _04545_, _04466_);
  and (_04547_, _04546_, cy_reg);
  or (_04548_, _04547_, _04544_);
  nor (_04549_, _04548_, _02425_);
  and (_04550_, _04548_, _02425_);
  nor (_04551_, _04289_, cy_reg);
  nor (_04552_, _04330_, _04328_);
  or (_04553_, _04552_, _04461_);
  nand (_04554_, _04552_, _04461_);
  and (_04555_, _04554_, _04553_);
  and (_04556_, _04555_, cy_reg);
  or (_04557_, _04556_, _04551_);
  nor (_04558_, _04557_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04559_, _04557_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_04560_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_04561_, _04454_, _04452_);
  not (_04562_, _04561_);
  and (_04563_, _04455_, cy_reg);
  and (_04564_, _04563_, _04562_);
  nor (_04565_, _04564_, _04560_);
  nor (_04566_, _04565_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_04567_, _04451_, _04503_);
  not (_04568_, _04567_);
  nor (_04569_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04570_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04571_, _04570_, _04569_);
  nor (_04572_, _04571_, _04568_);
  and (_04573_, _04571_, _04568_);
  or (_04574_, _04573_, _04572_);
  and (_04575_, _04565_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_04576_, _04575_, _04574_);
  or (_04577_, _04576_, _04566_);
  nor (_04578_, _04333_, cy_reg);
  or (_04579_, _04459_, _04457_);
  and (_04580_, _04579_, _04460_);
  and (_04581_, _04580_, cy_reg);
  nor (_04582_, _04581_, _04578_);
  nor (_04583_, _04582_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04584_, _04582_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_04585_, _04584_, _04583_);
  or (_04586_, _04585_, _04577_);
  or (_04587_, _04586_, _04559_);
  or (_04588_, _04587_, _04558_);
  or (_04589_, _04588_, _04550_);
  or (_04590_, _04589_, _04549_);
  or (_04591_, _04590_, _04543_);
  or (_04592_, _04591_, _04542_);
  or (_04593_, _04592_, _04536_);
  or (_04594_, _04593_, _04535_);
  or (_04595_, _04594_, _04529_);
  or (_04596_, _04595_, _04528_);
  or (_04597_, _04596_, _04520_);
  or (_04598_, _04597_, _04519_);
  or (_04599_, _04598_, _04513_);
  or (_04600_, _04599_, _04512_);
  and (_04601_, _04138_, _04503_);
  or (_04602_, _04478_, _04146_);
  and (_04603_, _04602_, _04479_);
  and (_04604_, _04603_, cy_reg);
  or (_04605_, _04604_, _04601_);
  nor (_04606_, _04605_, _02399_);
  and (_04607_, _04605_, _02399_);
  or (_04608_, _04607_, _04606_);
  or (_04609_, _04608_, _04600_);
  or (_04610_, _04609_, _04502_);
  or (_04611_, _04610_, _04501_);
  and (_04612_, _04131_, _04503_);
  or (_04613_, _04483_, _04481_);
  and (_04614_, _04613_, _04484_);
  and (_04615_, _04614_, cy_reg);
  or (_04616_, _04615_, _04612_);
  nor (_04617_, _04616_, _13154_);
  and (_04618_, _04616_, _13154_);
  or (_04619_, _04618_, _04617_);
  or (_04620_, _04619_, _04611_);
  or (_04621_, _04620_, _04492_);
  or (_04622_, _04621_, _04491_);
  and (_04623_, _04023_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04624_, _04023_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04625_, _04624_, _04623_);
  and (_04626_, _04625_, _04503_);
  or (_04627_, _04484_, _04129_);
  and (_04628_, _04132_, _13116_);
  nor (_04629_, _04628_, _04126_);
  nand (_04630_, _04629_, _04627_);
  and (_04631_, _04625_, _04125_);
  nor (_04632_, _04625_, _04125_);
  nor (_04633_, _04632_, _04631_);
  nand (_04634_, _04633_, _04630_);
  or (_04635_, _04633_, _04630_);
  and (_04636_, _04635_, _04634_);
  and (_04637_, _04636_, cy_reg);
  nor (_04638_, _04637_, _04626_);
  nor (_04639_, _04638_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_04640_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand (_04641_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_04642_, _04641_, _04640_);
  or (_04643_, _04642_, _04623_);
  nand (_04644_, _04642_, _04623_);
  and (_04645_, _04644_, _04643_);
  not (_04646_, _04645_);
  and (_04647_, _04630_, _04125_);
  not (_04648_, _04625_);
  nor (_04649_, _04630_, _04648_);
  or (_04650_, _04632_, _04503_);
  or (_04651_, _04650_, _04649_);
  or (_04652_, _04651_, _04647_);
  nand (_04653_, _04652_, _04646_);
  or (_04654_, _04652_, _04646_);
  and (_04655_, _04654_, _04653_);
  and (_04656_, _04638_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_04657_, _04656_, _04655_);
  or (_04658_, _04657_, _04639_);
  or (_04659_, _04658_, _04622_);
  nor (_04660_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_04661_, _04660_, _13036_);
  nor (_04662_, _04661_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04663_, _04661_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_04664_, _04663_, _04662_);
  or (_04665_, _00677_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_04666_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_04667_, _04666_, _04665_);
  or (_04668_, _04667_, _04664_);
  and (_04669_, _04660_, _13036_);
  nor (_04670_, _04669_, _04661_);
  not (_04671_, _04670_);
  or (_04672_, _00677_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_04673_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_04674_, _04673_, _04672_);
  nand (_04675_, _04674_, _04664_);
  and (_04676_, _04675_, _04671_);
  and (_04677_, _04676_, _04668_);
  and (_04678_, _04664_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_04679_, _02407_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_04680_, _04679_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_04681_, _04680_, _04678_);
  and (_04682_, _04664_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_04683_, _02407_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_04684_, _04683_, _00677_);
  or (_04685_, _04684_, _04682_);
  and (_04686_, _04685_, _04670_);
  and (_04687_, _04686_, _04681_);
  or (_04688_, _04687_, _04677_);
  and (_04689_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04690_, _04689_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_04691_, _04689_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_04692_, _04691_, _04690_);
  not (_04693_, _04692_);
  nor (_04694_, _04690_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04695_, _04690_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_04696_, _04695_, _04694_);
  nand (_04697_, _04696_, _07691_);
  or (_04698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_04699_, _04698_, _04697_);
  or (_04700_, _04699_, _04693_);
  nor (_04701_, _04696_, _04067_);
  and (_04702_, _04696_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_04703_, _04702_, _04701_);
  or (_04704_, _04703_, _04692_);
  and (_04705_, _04704_, _04700_);
  or (_04706_, _04705_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04707_, _04696_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_04708_, _04696_, _07686_);
  or (_04709_, _04708_, _04707_);
  and (_04710_, _04709_, _04693_);
  nand (_04711_, _04696_, _07696_);
  or (_04712_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_04713_, _04712_, _04692_);
  and (_04714_, _04713_, _04711_);
  or (_04715_, _04714_, _00677_);
  or (_04716_, _04715_, _04710_);
  and (_04717_, _02407_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_04718_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [15]);
  or (_04719_, _04718_, _04717_);
  and (_04720_, _04719_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_04721_, _02407_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_04722_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_04723_, _04722_, _13036_);
  and (_04724_, _04723_, _04721_);
  or (_04725_, _04724_, _04720_);
  and (_04726_, _04725_, _04689_);
  and (_04727_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], _00677_);
  or (_04728_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_04729_, _02407_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_04730_, _04729_, _04728_);
  or (_04731_, _04730_, _13036_);
  or (_04732_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_04733_, _02407_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_04734_, _04733_, _04732_);
  or (_04735_, _04734_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04736_, _04735_, _04731_);
  and (_04737_, _04736_, _04727_);
  or (_04738_, _04737_, _04726_);
  and (_04739_, _04725_, _00677_);
  and (_04740_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04741_, _04740_, _04730_);
  or (_04742_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_04743_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_04744_, _02407_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_04745_, _04744_, _04743_);
  and (_04746_, _04745_, _04742_);
  or (_04747_, _04746_, _04741_);
  or (_04748_, _04747_, _04739_);
  and (_04749_, _04748_, _04738_);
  and (_04750_, _04749_, _04716_);
  and (_04751_, _04750_, _04706_);
  and (_04752_, _04751_, _04688_);
  and (_04753_, _04664_, \oc8051_symbolic_cxrom1.regvalid [15]);
  or (_04754_, _04717_, _04671_);
  or (_04755_, _04754_, _04753_);
  and (_04756_, _04755_, _00677_);
  nand (_04757_, _04664_, _08257_);
  or (_04758_, _04664_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_04759_, _04758_, _04757_);
  or (_04760_, _04759_, _04670_);
  and (_04761_, _04760_, _04756_);
  or (_04762_, _04761_, _04747_);
  and (_04763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_04764_, _02407_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_04765_, _04764_, _04763_);
  and (_04766_, _04765_, _13036_);
  and (_04767_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_04768_, _04767_, _04679_);
  and (_04769_, _04768_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_04770_, _04769_, _04766_);
  and (_04771_, _04770_, _00677_);
  nand (_04772_, _04696_, _07614_);
  and (_04773_, _04728_, _04692_);
  and (_04774_, _04773_, _04772_);
  nand (_04775_, _04696_, _07661_);
  or (_04776_, _04696_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_04777_, _04776_, _04693_);
  and (_04778_, _04777_, _04775_);
  or (_04779_, _04778_, _04774_);
  and (_04780_, _04779_, _04771_);
  not (_04781_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand (_04782_, _04696_, _04781_);
  or (_04783_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_04784_, _04783_, _04692_);
  and (_04785_, _04784_, _04782_);
  or (_04786_, _04696_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand (_04787_, _04696_, _08257_);
  and (_04788_, _04787_, _04693_);
  and (_04789_, _04788_, _04786_);
  or (_04790_, _04789_, _04785_);
  and (_04791_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_04792_, _04683_, _13036_);
  or (_04793_, _04792_, _04791_);
  or (_04794_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_04795_, _02407_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_04796_, _04795_, _04794_);
  or (_04797_, _04796_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04798_, _04797_, _04793_);
  and (_04799_, _04798_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04800_, _04768_, _04740_);
  or (_04801_, _02407_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_04802_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_04803_, _04802_, _04743_);
  and (_04804_, _04803_, _04801_);
  or (_04805_, _04804_, _04800_);
  and (_04806_, _04805_, _04799_);
  and (_04807_, _04806_, _04790_);
  or (_04808_, _04807_, _04780_);
  or (_04809_, _04805_, _04798_);
  and (_04810_, _04809_, _02411_);
  and (_04811_, _04810_, _04808_);
  and (_04812_, _04811_, _04762_);
  or (_04813_, _04812_, _04752_);
  nor (_04814_, _04048_, _02418_);
  and (_04815_, _04048_, _02418_);
  nor (_04816_, _04815_, _04814_);
  nor (_04817_, _04814_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04818_, _04814_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04819_, _04818_, _04817_);
  nand (_04820_, _04819_, _07691_);
  or (_04821_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_04822_, _04821_, _04027_);
  and (_04823_, _04822_, _04820_);
  nand (_04824_, _04819_, _07696_);
  or (_04825_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_04826_, _04825_, _04061_);
  and (_04827_, _04826_, _04824_);
  or (_04828_, _04827_, _04823_);
  nand (_04829_, _04819_, _04781_);
  or (_04830_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_04831_, _04830_, _04048_);
  and (_04832_, _04831_, _04829_);
  nand (_04833_, _04819_, _07614_);
  or (_04834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_04835_, _04834_, _04073_);
  and (_04836_, _04835_, _04833_);
  or (_04837_, _04836_, _04832_);
  or (_04838_, _04837_, _04828_);
  and (_04839_, _04838_, _04816_);
  and (_04840_, _04819_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_04841_, _04819_, _04067_);
  or (_04842_, _04841_, _04840_);
  and (_04843_, _04842_, _04027_);
  and (_04844_, _04819_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_04845_, _04819_, _07686_);
  or (_04846_, _04845_, _04844_);
  and (_04847_, _04846_, _04061_);
  or (_04848_, _04847_, _04843_);
  and (_04849_, _04819_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_04850_, _04819_, _07645_);
  or (_04851_, _04850_, _04849_);
  and (_04852_, _04851_, _04048_);
  and (_04853_, _04819_, \oc8051_symbolic_cxrom1.regvalid [9]);
  not (_04854_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_04855_, _04819_, _04854_);
  or (_04856_, _04855_, _04853_);
  and (_04857_, _04856_, _04073_);
  or (_04858_, _04857_, _04852_);
  nor (_04859_, _04858_, _04848_);
  nor (_04860_, _04859_, _04816_);
  or (_04861_, _04860_, _04839_);
  or (_04862_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand (_04863_, _04862_, _04048_);
  and (_04864_, _04863_, _02418_);
  or (_04865_, \oc8051_symbolic_cxrom1.regarray[3] [3], \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand (_04866_, _04865_, _04027_);
  or (_04867_, \oc8051_symbolic_cxrom1.regarray[1] [3], \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand (_04868_, _04867_, _04061_);
  and (_04869_, _04868_, _04866_);
  or (_04870_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nand (_04871_, _04870_, _04073_);
  or (_04872_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nand (_04873_, _04872_, _04048_);
  and (_04874_, _04873_, _04871_);
  and (_04875_, _04874_, _04869_);
  and (_04876_, _04875_, _04864_);
  nand (_04877_, _04061_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  or (_04878_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nand (_04879_, _04878_, _04073_);
  and (_04880_, _04879_, _04877_);
  or (_04881_, \oc8051_symbolic_cxrom1.regarray[3] [5], \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nand (_04882_, _04881_, _04027_);
  or (_04883_, \oc8051_symbolic_cxrom1.regarray[1] [5], \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nand (_04884_, _04883_, _04061_);
  and (_04885_, _04884_, _04882_);
  and (_04886_, _04885_, _04880_);
  nand (_04887_, _04073_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  or (_04888_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nand (_04889_, _04888_, _04048_);
  and (_04890_, _04889_, _04887_);
  nand (_04891_, _04027_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_04892_, _04048_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_04893_, _04892_, _04891_);
  and (_04894_, _04893_, _04890_);
  and (_04895_, _04894_, _04886_);
  and (_04896_, _04048_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_04897_, _04061_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or (_04898_, _04897_, _04896_);
  and (_04899_, _04073_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_04900_, _04027_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  or (_04901_, _04900_, _04899_);
  or (_04902_, _04901_, _04898_);
  or (_04903_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand (_04904_, _04903_, _04073_);
  or (_04905_, \oc8051_symbolic_cxrom1.regarray[3] [1], \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand (_04906_, _04905_, _04027_);
  or (_04907_, \oc8051_symbolic_cxrom1.regarray[1] [1], \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand (_04908_, _04907_, _04061_);
  and (_04909_, _04908_, _04906_);
  and (_04910_, _04909_, _04904_);
  and (_04911_, _04910_, _04902_);
  and (_04912_, _04911_, _04895_);
  and (_04913_, _04912_, _04876_);
  or (_04914_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nand (_04915_, _04914_, _04073_);
  and (_04916_, _04915_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_04917_, \oc8051_symbolic_cxrom1.regarray[7] [5], \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nand (_04918_, _04917_, _04027_);
  or (_04919_, \oc8051_symbolic_cxrom1.regarray[5] [5], \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nand (_04920_, _04919_, _04061_);
  and (_04921_, _04920_, _04918_);
  or (_04922_, \oc8051_symbolic_cxrom1.regarray[7] [1], \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nand (_04923_, _04922_, _04027_);
  or (_04924_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand (_04925_, _04924_, _04073_);
  and (_04926_, _04925_, _04923_);
  and (_04927_, _04926_, _04921_);
  and (_04928_, _04927_, _04916_);
  or (_04929_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand (_04930_, _04929_, _04048_);
  or (_04931_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand (_04932_, _04931_, _04073_);
  and (_04933_, _04932_, _04930_);
  or (_04934_, \oc8051_symbolic_cxrom1.regarray[7] [3], \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand (_04935_, _04934_, _04027_);
  or (_04936_, \oc8051_symbolic_cxrom1.regarray[5] [3], \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand (_04937_, _04936_, _04061_);
  and (_04938_, _04937_, _04935_);
  and (_04939_, _04938_, _04933_);
  nand (_04940_, _04073_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  or (_04941_, \oc8051_symbolic_cxrom1.regarray[5] [1], \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand (_04942_, _04941_, _04061_);
  and (_04943_, _04942_, _04940_);
  nand (_04944_, _04027_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_04945_, _04048_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_04946_, _04945_, _04944_);
  and (_04947_, _04946_, _04943_);
  and (_04948_, _04947_, _04939_);
  and (_04949_, _04061_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_04950_, _04048_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or (_04951_, _04950_, _04949_);
  and (_04952_, _04027_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_04953_, _04073_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  or (_04954_, _04953_, _04952_);
  or (_04955_, _04954_, _04951_);
  or (_04956_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand (_04957_, _04956_, _04048_);
  nand (_04958_, _04061_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  or (_04959_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nand (_04960_, _04959_, _04048_);
  and (_04961_, _04960_, _04958_);
  and (_04962_, _04961_, _04957_);
  and (_04963_, _04962_, _04955_);
  and (_04964_, _04963_, _04948_);
  and (_04965_, _04964_, _04928_);
  or (_04966_, _04965_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_04967_, _04966_, _04913_);
  nor (_04968_, _02383_, first_instr);
  and (_04969_, _04968_, _04967_);
  nor (_04970_, \oc8051_symbolic_cxrom1.regarray[13] [1], \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_04971_, \oc8051_symbolic_cxrom1.regarray[13] [3], \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand (_04972_, _04971_, _04970_);
  nand (_04973_, _04972_, _04061_);
  nor (_04974_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_04975_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand (_04976_, _04975_, _04974_);
  nand (_04977_, _04976_, _04073_);
  not (_04978_, _04027_);
  nor (_04979_, \oc8051_symbolic_cxrom1.regarray[15] [3], \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_04980_, \oc8051_symbolic_cxrom1.regarray[15] [1], \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_04981_, _04980_, _04979_);
  or (_04982_, _04981_, _04978_);
  and (_04983_, _04982_, _04977_);
  and (_04984_, _04983_, _04973_);
  nand (_04985_, _04027_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_04986_, _04048_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_04987_, _04986_, _04985_);
  nand (_04988_, _04061_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  or (_04989_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nand (_04990_, _04989_, _04073_);
  and (_04991_, _04990_, _04988_);
  and (_04992_, _04991_, _04987_);
  not (_04993_, _04048_);
  nor (_04994_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_04995_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_04996_, _04995_, _04994_);
  or (_04997_, _04996_, _04993_);
  nand (_04998_, _04073_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_04999_, _04998_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05000_, _04999_, _04997_);
  and (_05001_, _05000_, _04992_);
  and (_05002_, _04027_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_05003_, _04073_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or (_05004_, _05003_, _05002_);
  and (_05005_, _04061_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_05006_, _04048_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or (_05007_, _05006_, _05005_);
  or (_05008_, _05007_, _05004_);
  or (_05009_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nand (_05010_, _05009_, _04048_);
  or (_05011_, \oc8051_symbolic_cxrom1.regarray[15] [5], \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nand (_05012_, _05011_, _04027_);
  or (_05013_, \oc8051_symbolic_cxrom1.regarray[13] [5], \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nand (_05014_, _05013_, _04061_);
  and (_05015_, _05014_, _05012_);
  and (_05016_, _05015_, _05010_);
  and (_05017_, _05016_, _05008_);
  and (_05018_, _05017_, _05001_);
  and (_05019_, _05018_, _04984_);
  nor (_05020_, \oc8051_symbolic_cxrom1.regarray[11] [3], \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_05021_, \oc8051_symbolic_cxrom1.regarray[11] [1], \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_05022_, _05021_, _05020_);
  or (_05023_, _05022_, _04978_);
  nor (_05024_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_05025_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_05026_, _05025_, _05024_);
  or (_05027_, _05026_, _04993_);
  nor (_05028_, \oc8051_symbolic_cxrom1.regarray[9] [1], \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_05029_, \oc8051_symbolic_cxrom1.regarray[9] [3], \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand (_05030_, _05029_, _05028_);
  nand (_05031_, _05030_, _04061_);
  and (_05032_, _05031_, _05027_);
  and (_05033_, _05032_, _05023_);
  or (_05034_, \oc8051_symbolic_cxrom1.regarray[9] [5], \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nand (_05035_, _05034_, _04061_);
  or (_05036_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nand (_05037_, _05036_, _04073_);
  and (_05038_, _05037_, _05035_);
  nand (_05039_, _04073_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nand (_05040_, _04073_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_05041_, _05040_, _05039_);
  and (_05042_, _05041_, _05038_);
  or (_05043_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nand (_05044_, _05043_, _04073_);
  and (_05045_, _05044_, _02418_);
  or (_05046_, \oc8051_symbolic_cxrom1.regarray[11] [5], \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nand (_05047_, _05046_, _04027_);
  or (_05048_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nand (_05049_, _05048_, _04048_);
  and (_05050_, _05049_, _05047_);
  and (_05051_, _05050_, _05045_);
  and (_05052_, _05051_, _05042_);
  nand (_05053_, _04073_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_05054_, _04061_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_05055_, _05054_, _05053_);
  nand (_05056_, _04027_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_05057_, _04048_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_05058_, _05057_, _05056_);
  and (_05059_, _05058_, _05055_);
  and (_05060_, _04027_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_05061_, _04073_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  or (_05062_, _05061_, _05060_);
  and (_05063_, _04048_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_05064_, _04061_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or (_05065_, _05064_, _05063_);
  or (_05066_, _05065_, _05062_);
  and (_05067_, _05066_, _05059_);
  and (_05068_, _05067_, _05052_);
  and (_05069_, _05068_, _05033_);
  or (_05070_, _05069_, _07607_);
  or (_05071_, _05070_, _05019_);
  or (_05072_, _07607_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_05073_, _04821_, _05072_);
  or (_05074_, _05073_, _02418_);
  or (_05075_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_05076_, _07607_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05077_, _05076_, _05075_);
  or (_05078_, _05077_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05079_, _05078_, _05074_);
  and (_05080_, _05079_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_05081_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_05082_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05083_, _07607_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05084_, _05083_, _05082_);
  and (_05085_, _05084_, _05081_);
  or (_05086_, _07607_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_05087_, _05086_, _04825_);
  and (_05088_, _05087_, _04332_);
  or (_05089_, _05088_, _05085_);
  or (_05090_, _05089_, _05080_);
  and (_05091_, _05079_, _02390_);
  and (_05092_, _05087_, _04331_);
  or (_05093_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05094_, _07607_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05095_, _05094_, _04012_);
  and (_05096_, _05095_, _05093_);
  or (_05097_, _05096_, _05092_);
  or (_05098_, _05097_, _05091_);
  and (_05099_, _05098_, _04009_);
  and (_05100_, _05099_, _05090_);
  or (_05101_, _07607_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_05102_, _04830_, _05101_);
  or (_05103_, _05102_, _02418_);
  or (_05104_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_05105_, _07607_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05106_, _05105_, _05104_);
  or (_05107_, _05106_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05108_, _05107_, _05103_);
  and (_05109_, _05108_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_05110_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05111_, _07607_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05112_, _05111_, _05110_);
  and (_05113_, _05112_, _05081_);
  or (_05114_, _07607_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_05115_, _05114_, _04834_);
  and (_05116_, _05115_, _04332_);
  or (_05117_, _05116_, _05113_);
  or (_05118_, _05117_, _05109_);
  and (_05119_, _05108_, _02390_);
  and (_05120_, _05115_, _04331_);
  or (_05121_, _07607_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05122_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05123_, _05122_, _04012_);
  and (_05124_, _05123_, _05121_);
  or (_05125_, _05124_, _05120_);
  or (_05126_, _05125_, _05119_);
  and (_05127_, _05126_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05128_, _05127_, _05118_);
  or (_05129_, _05128_, _05100_);
  and (_05130_, _05129_, _05071_);
  and (_05131_, _05130_, _04969_);
  and (_05133_, _05131_, _04861_);
  and (_05134_, _05133_, _04335_);
  and (_05135_, _05134_, _04813_);
  and (property_invalid_jc, _05135_, _04659_);
  or (_05136_, pc_log_change_r, _04503_);
  nand (_05137_, pc_log_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_00000_, _05137_, _05136_);
  and (_05138_, _02383_, first_instr);
  or (_00001_, _05138_, rst);
  dff (cy_reg, _00000_);
  dff (pc_log_change_r, pc_log_change);
  dff (first_instr, _00001_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _08867_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _08870_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _08873_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _08877_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _08879_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _08882_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _08887_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _06058_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _08770_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _08775_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _08777_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _08781_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _08785_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _08788_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _08792_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _08796_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _13483_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _13484_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _13485_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _08679_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _13486_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _13487_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _13488_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _13489_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _13475_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _13476_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _13477_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _13478_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _13479_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _13480_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _13481_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _13482_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _08486_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _08490_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _08493_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _08495_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _08498_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _08502_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _08506_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _08510_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _08400_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _08403_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _08407_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _08410_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _08413_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _08416_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _08419_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _08421_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _08310_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _08314_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _08317_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _08321_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _08325_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _08329_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _08331_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _08335_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _13495_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _08219_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _08224_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _08229_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _08234_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _08236_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _08240_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _08244_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _08120_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _08123_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _13490_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _13491_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _13492_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _13493_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _13494_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _08141_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _08042_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _08045_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _08048_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _08051_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _08053_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _08056_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _08058_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _08060_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _07953_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _07957_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _07961_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _07965_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _07969_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _07971_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _07974_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _07976_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _07553_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _07558_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _07562_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _07565_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _07569_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _07573_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _07575_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _07578_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _07443_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _07449_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _07454_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _07460_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _07465_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _07470_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _07475_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _07477_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _07755_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _07760_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _07762_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _07764_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _07767_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _07770_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _07775_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _07778_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _07655_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _07660_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _07664_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _07667_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _07672_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _07677_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _07682_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _07687_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _07863_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _07866_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _07869_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _07873_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _07876_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _07879_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _07881_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _07885_);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _06079_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _06108_);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _06149_);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _06196_);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _06252_);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _06294_);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _06359_);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _06435_);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _06513_);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _06609_);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _06704_);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _06794_);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _06887_);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _06971_);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _07082_);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _06029_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _05726_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _05729_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _05732_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _05735_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _05738_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _05741_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _05744_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _05596_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _10940_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _10986_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _12116_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _12113_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _12104_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _05756_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _12082_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _05599_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _05760_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _12791_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _05764_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _05767_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _05770_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _12656_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _12109_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _03035_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _11697_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _11719_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _06984_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _08889_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _05304_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _11658_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _05369_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _11638_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _02768_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _05558_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _09689_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _09833_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _09859_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _09855_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _09862_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _11677_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _00855_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _03039_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _11679_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _03080_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _05235_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _03150_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _03152_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05238_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _03195_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _03198_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05251_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _03316_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _05340_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _03634_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _03637_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _03698_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _01783_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _03806_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _05502_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _05451_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _03849_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _03910_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _13174_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _11890_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _05139_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _03936_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _00349_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _02876_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _08473_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _02698_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _02137_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _07122_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _04141_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _01027_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _03049_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _02871_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _03622_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _02780_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _05140_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _03779_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _02888_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _03745_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _02194_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _02863_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _06673_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _06443_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _06424_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _06258_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _06405_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _06712_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _03920_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _03995_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _03300_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _08821_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _00486_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _02915_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _00457_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _05468_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _01578_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _02935_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _07680_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _12536_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _03623_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _11360_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _02660_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _07670_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _03372_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _02925_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _13260_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _07247_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _10437_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _01842_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _09109_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _07658_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _01927_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _04083_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _00002_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _01183_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _06783_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _00302_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _12994_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _12316_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _12641_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _12620_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _01890_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _01564_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _01467_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _01451_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _10557_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _02738_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _13067_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _10800_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _02734_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _02771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _02067_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _03319_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _02730_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _01582_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _02103_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _02726_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _02806_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _02701_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _01756_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _02723_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _13030_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _04103_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _02715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _02760_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _05932_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _03601_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _02713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _07446_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _03854_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _02710_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _02759_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _02797_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _02804_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _11239_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _11104_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _02705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _13021_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _11979_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _10750_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _10890_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _01733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _12623_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _03884_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _01824_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _11995_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _06232_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _08991_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _01626_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _07749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _02840_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _11987_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _10747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _03871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _03888_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _03886_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _03882_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _03876_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _12016_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _04059_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _03998_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _03997_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _03933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _03912_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _12008_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _10742_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _10887_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _10943_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _03795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _03033_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _02832_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _02999_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _03045_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _03021_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _03011_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _03006_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _12076_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _03183_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _10555_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _03031_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _10656_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _10936_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _00706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _00684_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _00670_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _00660_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _00657_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _12157_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _00826_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _00807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _00788_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _00778_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _12146_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _10715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _00387_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _00357_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _10647_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _12218_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _00147_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _00209_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _00172_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _00158_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _12212_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _10698_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _11034_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _11077_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _11068_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _11063_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _12227_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _13411_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _13436_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _13431_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _10640_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _02830_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _10388_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _10340_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _12738_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _12018_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _12013_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _11993_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _11975_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _11968_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _12734_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _10382_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _11632_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _11616_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _10377_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _10510_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _11346_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _11335_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _11323_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _11319_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _12661_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _12648_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _12767_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _10503_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _10494_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _10476_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _11229_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _11523_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _11515_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _10458_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _11645_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _11641_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _11107_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _11221_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _11263_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _11666_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _11664_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _11100_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _11675_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _11670_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _11098_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _11217_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _11688_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _11682_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _11703_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _11695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _11094_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _11214_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _11259_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _11310_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11389_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _11376_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _11163_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _11416_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _11409_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _11161_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _11236_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _11363_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _11356_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _11166_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _11281_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _02828_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _10251_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _10245_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _03037_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _11921_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _11030_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _11300_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _11947_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _10319_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _00911_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _03835_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _03700_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _03731_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _00666_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _03643_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _03709_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _03688_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _03716_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _03728_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _03983_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _03979_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _03993_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _03989_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _01025_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _12630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _07160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _06507_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _03193_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _07061_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _03305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _03180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _06503_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _05329_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _13367_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _13352_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _02397_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _13387_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _13380_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _02394_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _13332_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _03923_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _05720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _05717_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _05714_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _05707_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _05690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _05687_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _05698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _02221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _05790_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _05783_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _01188_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _10236_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _05793_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _05780_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _01207_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _01651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _09119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _01389_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _01479_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _01473_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00980_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _01500_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _01484_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00978_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _03087_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _01503_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _07816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _10115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _01392_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _01459_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _10191_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _01516_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _01511_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _07981_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _01523_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _01540_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _07616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _08859_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _07277_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _07206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _01005_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _01395_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _01465_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _10153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _01545_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _01543_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00899_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _01553_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _01548_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00890_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _01032_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _10239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _01758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _01585_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _01764_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _01762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00853_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _01030_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _07297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _02504_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _02658_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _02526_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _02502_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _02664_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _02529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _02661_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _02824_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _02635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _02523_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _02499_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _02670_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _02525_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _02668_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _02522_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _03856_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _02501_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _02666_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _02634_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _02615_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _02613_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _02519_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _02495_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _00987_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _02493_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _02672_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _02640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _02638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _02679_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _02517_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _02677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _03119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _09173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _09170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _01779_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _09564_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _09572_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _09569_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _03139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _02431_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _12861_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _12858_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _12856_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _12854_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _02429_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _12788_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _13205_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _13207_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _00366_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _00370_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _12090_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _12098_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _12102_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _12073_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _12070_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _12067_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _12080_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _00379_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _12125_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _12119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _12122_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _12143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _12134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _12140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _12137_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _00374_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _00377_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _00376_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _12160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _12154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _12180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _12190_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _12187_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _12246_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _12242_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _00341_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _12328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _12324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _12295_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _12298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _12307_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _12311_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _12284_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _00345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _00343_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _12334_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _12337_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _12348_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _12342_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _12345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _12360_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _12353_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _00355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01883_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01921_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01917_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01888_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _11180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _05132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _12210_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _12206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _12203_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _12198_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _06991_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01886_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _12183_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _12163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _12128_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _07075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _01149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _12058_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _07095_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01853_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01874_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _07098_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _03908_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _03017_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _10570_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _10610_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _10583_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _10575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01871_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _10461_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _10499_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _10492_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _10489_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _11254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _10529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _10540_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01868_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _10347_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _10344_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _12002_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _10417_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _10412_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _10409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _10406_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01860_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _03178_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _03175_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _03172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _03170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _03168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _03143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _03141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _03136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _03134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _03132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _03123_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _03818_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _07457_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _07493_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _10072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _02973_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _01681_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _06960_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _03090_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _03899_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _08477_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _08312_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _03603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _03894_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _09143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _04037_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _03904_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _03098_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _03074_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _02987_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _02897_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _03890_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _03816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _03777_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _03713_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _03523_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _06717_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _06903_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _06817_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _03519_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _08210_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _07165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _07038_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _08682_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _08517_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _10068_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _08691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _10792_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _10718_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _10871_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _03160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _06966_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _11700_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _11526_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _12085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _11717_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _06962_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _12406_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _03126_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _07027_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _12815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _12722_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _06957_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _13390_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _12925_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _07024_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _03067_);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [0], ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [1], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [2], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [3], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [4], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [5], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [6], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [7], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [8], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [9], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [10], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [11], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [12], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [13], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [14], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [15], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [16], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [0], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [1], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [2], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [3], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [4], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [5], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [6], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [7], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [0], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [1], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [2], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [3], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [4], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [5], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [6], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [7], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.mulOv , ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [0], ABINPUT000000[1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [1], ABINPUT000000[2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [2], ABINPUT000000[3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [3], ABINPUT000000[4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [4], ABINPUT000000[5]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [5], ABINPUT000000[6]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [6], ABINPUT000000[7]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [7], ABINPUT000000[8]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [0], ABINPUT000000[9]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [1], ABINPUT000000[10]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], ABINPUT000000[11]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], ABINPUT000000[12]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], ABINPUT000000[13]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], ABINPUT000000[14]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], ABINPUT000000[15]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], ABINPUT000000[16]);
  buf(\oc8051_top_1.oc8051_alu1.divOv , ABINPUT000000[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [0], ABINPUT000000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [1], ABINPUT000000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [2], ABINPUT000000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [3], ABINPUT000000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [4], ABINPUT000000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [5], ABINPUT000000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [6], ABINPUT000000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [7], ABINPUT000000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [8], ABINPUT000000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [9], ABINPUT000000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [10], ABINPUT000000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [11], ABINPUT000000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [12], ABINPUT000000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [13], ABINPUT000000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [14], ABINPUT000000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [15], ABINPUT000000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [16], ABINPUT000000[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.ABINPUT000 [0], ABINPUT000[0]);
  buf(\oc8051_top_1.ABINPUT000 [1], ABINPUT000[1]);
  buf(\oc8051_top_1.ABINPUT000 [2], ABINPUT000[2]);
  buf(\oc8051_top_1.ABINPUT000 [3], ABINPUT000[3]);
  buf(\oc8051_top_1.ABINPUT000 [4], ABINPUT000[4]);
  buf(\oc8051_top_1.ABINPUT000 [5], ABINPUT000[5]);
  buf(\oc8051_top_1.ABINPUT000 [6], ABINPUT000[6]);
  buf(\oc8051_top_1.ABINPUT000 [7], ABINPUT000[7]);
  buf(\oc8051_top_1.ABINPUT000 [8], ABINPUT000[8]);
  buf(\oc8051_top_1.ABINPUT000 [9], ABINPUT000[9]);
  buf(\oc8051_top_1.ABINPUT000 [10], ABINPUT000[10]);
  buf(\oc8051_top_1.ABINPUT000 [11], ABINPUT000[11]);
  buf(\oc8051_top_1.ABINPUT000 [12], ABINPUT000[12]);
  buf(\oc8051_top_1.ABINPUT000 [13], ABINPUT000[13]);
  buf(\oc8051_top_1.ABINPUT000 [14], ABINPUT000[14]);
  buf(\oc8051_top_1.ABINPUT000 [15], ABINPUT000[15]);
  buf(\oc8051_top_1.ABINPUT000 [16], ABINPUT000[16]);
  buf(\oc8051_top_1.ABINPUT000000 [0], ABINPUT000000[0]);
  buf(\oc8051_top_1.ABINPUT000000 [1], ABINPUT000000[1]);
  buf(\oc8051_top_1.ABINPUT000000 [2], ABINPUT000000[2]);
  buf(\oc8051_top_1.ABINPUT000000 [3], ABINPUT000000[3]);
  buf(\oc8051_top_1.ABINPUT000000 [4], ABINPUT000000[4]);
  buf(\oc8051_top_1.ABINPUT000000 [5], ABINPUT000000[5]);
  buf(\oc8051_top_1.ABINPUT000000 [6], ABINPUT000000[6]);
  buf(\oc8051_top_1.ABINPUT000000 [7], ABINPUT000000[7]);
  buf(\oc8051_top_1.ABINPUT000000 [8], ABINPUT000000[8]);
  buf(\oc8051_top_1.ABINPUT000000 [9], ABINPUT000000[9]);
  buf(\oc8051_top_1.ABINPUT000000 [10], ABINPUT000000[10]);
  buf(\oc8051_top_1.ABINPUT000000 [11], ABINPUT000000[11]);
  buf(\oc8051_top_1.ABINPUT000000 [12], ABINPUT000000[12]);
  buf(\oc8051_top_1.ABINPUT000000 [13], ABINPUT000000[13]);
  buf(\oc8051_top_1.ABINPUT000000 [14], ABINPUT000000[14]);
  buf(\oc8051_top_1.ABINPUT000000 [15], ABINPUT000000[15]);
  buf(\oc8051_top_1.ABINPUT000000 [16], ABINPUT000000[16]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
