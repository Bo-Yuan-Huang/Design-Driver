
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire [15:0] _26842_;
  wire [7:0] _26843_;
  wire [7:0] _26844_;
  wire [7:0] _26845_;
  wire [7:0] _26846_;
  wire [7:0] _26847_;
  wire [7:0] _26848_;
  wire [7:0] _26849_;
  wire [7:0] _26850_;
  wire [7:0] _26851_;
  wire [7:0] _26852_;
  wire [7:0] _26853_;
  wire [7:0] _26854_;
  wire [7:0] _26855_;
  wire [7:0] _26856_;
  wire [7:0] _26857_;
  wire [7:0] _26858_;
  wire _26859_;
  wire [7:0] _26860_;
  wire [2:0] _26861_;
  wire [2:0] _26862_;
  wire [1:0] _26863_;
  wire [7:0] _26864_;
  wire _26865_;
  wire [1:0] _26866_;
  wire [1:0] _26867_;
  wire [2:0] _26868_;
  wire [2:0] _26869_;
  wire [1:0] _26870_;
  wire [3:0] _26871_;
  wire [1:0] _26872_;
  wire _26873_;
  wire [7:0] _26874_;
  wire [7:0] _26875_;
  wire [7:0] _26876_;
  wire [7:0] _26877_;
  wire [7:0] _26878_;
  wire [7:0] _26879_;
  wire [7:0] _26880_;
  wire [7:0] _26881_;
  wire [15:0] _26882_;
  wire [15:0] _26883_;
  wire _26884_;
  wire [4:0] _26885_;
  wire [7:0] _26886_;
  wire [7:0] _26887_;
  wire _26888_;
  wire _26889_;
  wire [15:0] _26890_;
  wire [15:0] _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire [7:0] _26895_;
  wire [2:0] _26896_;
  wire [7:0] _26897_;
  wire _26898_;
  wire [7:0] _26899_;
  wire _26900_;
  wire _26901_;
  wire [3:0] _26902_;
  wire [31:0] _26903_;
  wire [31:0] _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire [15:0] _26908_;
  wire _26909_;
  wire _26910_;
  wire [7:0] _26911_;
  wire _26912_;
  wire [2:0] _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire [3:0] _27304_;
  wire _27305_;
  wire _27306_;
  wire [7:0] _27307_;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not (_22762_, rst);
  not (_22763_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  nor (_22764_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_22765_, _22764_, _22763_);
  not (_22766_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_22767_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_22768_, _22767_, _22766_);
  and (_22769_, _22768_, _22765_);
  and (_22770_, _22769_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_22771_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_22772_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_22773_, _22770_, _22772_);
  or (_22775_, _22773_, _22771_);
  and (_26882_[0], _22775_, _22762_);
  and (_22777_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_22778_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_22780_, _22770_, _22778_);
  or (_22781_, _22780_, _22777_);
  and (_26882_[1], _22781_, _22762_);
  and (_22782_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_22783_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_22784_, _22770_, _22783_);
  or (_22785_, _22784_, _22782_);
  and (_26882_[2], _22785_, _22762_);
  and (_22786_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_22788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_22789_, _22770_, _22788_);
  or (_22791_, _22789_, _22786_);
  and (_26882_[3], _22791_, _22762_);
  and (_22793_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_22794_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_22795_, _22770_, _22794_);
  or (_22796_, _22795_, _22793_);
  and (_26882_[4], _22796_, _22762_);
  and (_22797_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_22798_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_22799_, _22770_, _22798_);
  or (_22800_, _22799_, _22797_);
  and (_26882_[5], _22800_, _22762_);
  and (_22801_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_22802_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_22803_, _22770_, _22802_);
  or (_22804_, _22803_, _22801_);
  and (_26882_[6], _22804_, _22762_);
  and (_22805_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_22806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_22807_, _22770_, _22806_);
  or (_22808_, _22807_, _22805_);
  and (_26882_[7], _22808_, _22762_);
  and (_22809_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_22810_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_22811_, _22770_, _22810_);
  or (_22812_, _22811_, _22809_);
  and (_26882_[8], _22812_, _22762_);
  and (_22813_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not (_22814_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_22815_, _22770_, _22814_);
  or (_22816_, _22815_, _22813_);
  and (_26882_[9], _22816_, _22762_);
  and (_22817_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_22819_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_22820_, _22770_, _22819_);
  or (_22821_, _22820_, _22817_);
  and (_26882_[10], _22821_, _22762_);
  and (_22822_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_22823_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_22824_, _22770_, _22823_);
  or (_22825_, _22824_, _22822_);
  and (_26882_[11], _22825_, _22762_);
  and (_22826_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_22827_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_22828_, _22770_, _22827_);
  or (_22829_, _22828_, _22826_);
  and (_26882_[12], _22829_, _22762_);
  and (_22830_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_22832_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_22833_, _22770_, _22832_);
  or (_22834_, _22833_, _22830_);
  and (_26882_[13], _22834_, _22762_);
  and (_22836_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_22837_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_22838_, _22770_, _22837_);
  or (_22839_, _22838_, _22836_);
  and (_26882_[14], _22839_, _22762_);
  and (_22840_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_22841_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22842_, _22770_, _22841_);
  or (_22843_, _22842_, _22840_);
  and (_26883_[0], _22843_, _22762_);
  and (_22844_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_22845_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_22846_, _22770_, _22845_);
  or (_22847_, _22846_, _22844_);
  and (_26883_[1], _22847_, _22762_);
  and (_22848_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_22849_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_22850_, _22770_, _22849_);
  or (_22852_, _22850_, _22848_);
  and (_26883_[2], _22852_, _22762_);
  and (_22853_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_22854_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22855_, _22770_, _22854_);
  or (_22857_, _22855_, _22853_);
  and (_26883_[3], _22857_, _22762_);
  or (_22859_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nand (_22860_, _22770_, _22794_);
  and (_22861_, _22860_, _22762_);
  and (_26883_[4], _22861_, _22859_);
  and (_22862_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_22864_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_22865_, _22770_, _22864_);
  or (_22867_, _22865_, _22862_);
  and (_26883_[5], _22867_, _22762_);
  and (_22868_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_22869_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_22870_, _22770_, _22869_);
  or (_22871_, _22870_, _22868_);
  and (_26883_[6], _22871_, _22762_);
  and (_22872_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_22874_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_22875_, _22770_, _22874_);
  or (_22876_, _22875_, _22872_);
  and (_26883_[7], _22876_, _22762_);
  or (_22877_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nand (_22878_, _22770_, _22810_);
  and (_22879_, _22878_, _22762_);
  and (_26883_[8], _22879_, _22877_);
  and (_22881_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not (_22882_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_22883_, _22770_, _22882_);
  or (_22884_, _22883_, _22881_);
  and (_26883_[9], _22884_, _22762_);
  and (_22885_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  not (_22886_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_22887_, _22770_, _22886_);
  or (_22888_, _22887_, _22885_);
  and (_26883_[10], _22888_, _22762_);
  and (_22889_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not (_22890_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_22891_, _22770_, _22890_);
  or (_22892_, _22891_, _22889_);
  and (_26883_[11], _22892_, _22762_);
  or (_22893_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nand (_22894_, _22770_, _22827_);
  and (_22895_, _22894_, _22762_);
  and (_26883_[12], _22895_, _22893_);
  and (_22896_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_22897_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_22899_, _22770_, _22897_);
  or (_22900_, _22899_, _22896_);
  and (_26883_[13], _22900_, _22762_);
  or (_22901_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nand (_22903_, _22770_, _22837_);
  and (_22904_, _22903_, _22762_);
  and (_26883_[14], _22904_, _22901_);
  and (_22905_, \oc8051_top_1.oc8051_decoder1.wr , _22766_);
  not (_22906_, _22905_);
  not (_22907_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22908_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _22766_);
  and (_22909_, _22908_, _22907_);
  and (_22910_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_22912_, _22910_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_22913_, _22912_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_22914_, _22913_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_22915_, _22914_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_22917_, _22915_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_22918_, _22917_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  not (_22919_, _22918_);
  and (_22920_, _22909_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  or (_22921_, _22917_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and (_22922_, _22921_, _22920_);
  and (_22923_, _22922_, _22919_);
  not (_22924_, _22923_);
  and (_22926_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22927_, _22926_, _22908_);
  not (_22928_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_22929_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _22766_);
  and (_22930_, _22929_, _22928_);
  and (_22931_, _22930_, _22907_);
  and (_22932_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_22934_, _22932_, _22927_);
  nor (_22935_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22937_, _22935_, _22908_);
  and (_22938_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_22939_, _22930_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22940_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_22941_, _22940_, _22938_);
  and (_22942_, _22941_, _22934_);
  nand (_22943_, _22942_, _22924_);
  not (_22944_, _22943_);
  nor (_22945_, _22944_, _22909_);
  nor (_22946_, _22945_, _22906_);
  not (_22947_, _22946_);
  not (_22948_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_22949_, _22943_, _22948_);
  nor (_22950_, _22913_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_22951_, _22950_);
  not (_22952_, _22920_);
  nor (_22953_, _22952_, _22914_);
  and (_22954_, _22953_, _22951_);
  not (_22956_, _22954_);
  and (_22957_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor (_22958_, _22957_, _22927_);
  and (_22960_, _22935_, _22928_);
  or (_22961_, _22960_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_22962_, _22961_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_22963_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_22964_, _22963_, _22962_);
  and (_22966_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not (_22967_, _22966_);
  and (_22968_, _22967_, _22964_);
  and (_22969_, _22968_, _22958_);
  and (_22970_, _22969_, _22956_);
  not (_22971_, _22970_);
  and (_22972_, _22971_, _22949_);
  nor (_22973_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_22974_, _22973_, _22910_);
  and (_22975_, _22974_, _22920_);
  and (_22976_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_22977_, _22976_, _22975_);
  and (_22978_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_22979_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_22980_, _22961_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_22981_, _22980_, _22979_);
  nor (_22982_, _22981_, _22978_);
  and (_22983_, _22982_, _22977_);
  nor (_22984_, _22983_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_22985_, _22984_, _22972_);
  nor (_22986_, _22985_, _22947_);
  nor (_22987_, _22912_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_22989_, _22987_, _22913_);
  and (_22990_, _22989_, _22920_);
  not (_22991_, _22990_);
  and (_22992_, _22961_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_22994_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_22995_, _22994_, _22992_);
  and (_22996_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_22997_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_22999_, _22997_, _22996_);
  and (_23000_, _22999_, _22995_);
  and (_23002_, _23000_, _22991_);
  not (_23003_, _23002_);
  and (_23004_, _23003_, _22949_);
  and (_23005_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_23006_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_23008_, _23006_, _23005_);
  and (_23009_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not (_23011_, _23009_);
  not (_23012_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_23014_, _22920_, _23012_);
  and (_23015_, _22961_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_23016_, _23015_, _23014_);
  and (_23017_, _23016_, _23011_);
  and (_23018_, _23017_, _23008_);
  nor (_23019_, _23018_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23020_, _23019_, _23004_);
  and (_23021_, _23020_, _22986_);
  nor (_23022_, _22915_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_23023_, _23022_);
  nor (_23024_, _22952_, _22917_);
  and (_23025_, _23024_, _23023_);
  not (_23026_, _23025_);
  and (_23027_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_23028_, _23027_, _22927_);
  and (_23029_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_23030_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor (_23031_, _23030_, _23029_);
  and (_23033_, _23031_, _23028_);
  and (_23034_, _23033_, _23026_);
  not (_23035_, _23034_);
  and (_23036_, _23035_, _22949_);
  nor (_23038_, _23002_, _22949_);
  nor (_23039_, _23038_, _23036_);
  nor (_23040_, _23039_, _22947_);
  nor (_23041_, _22914_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_23042_, _23041_);
  nor (_23043_, _22952_, _22915_);
  and (_23044_, _23043_, _23042_);
  not (_23045_, _23044_);
  and (_23046_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_23047_, _23046_, _22927_);
  and (_23048_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_23049_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor (_23050_, _23049_, _23048_);
  and (_23051_, _23050_, _23047_);
  and (_23052_, _23051_, _23045_);
  not (_23053_, _23052_);
  and (_23054_, _23053_, _22949_);
  nor (_23055_, _22910_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_23056_, _23055_, _22912_);
  and (_23057_, _23056_, _22920_);
  and (_23058_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_23059_, _23058_, _23057_);
  and (_23060_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_23061_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_23062_, _22961_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_23063_, _23062_, _23061_);
  nor (_23064_, _23063_, _23060_);
  and (_23065_, _23064_, _23059_);
  nor (_23066_, _23065_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23067_, _23066_, _23054_);
  and (_23068_, _23067_, _23040_);
  and (_23069_, _23068_, _23021_);
  nor (_23070_, _22970_, _22949_);
  and (_23071_, _23070_, _22946_);
  and (_23072_, _23071_, _23053_);
  nor (_23073_, _23035_, _22943_);
  nor (_23074_, _23073_, _22949_);
  not (_23075_, _23074_);
  and (_23076_, _23075_, _23072_);
  and (_23077_, _23076_, _23069_);
  nor (_23078_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23079_, \oc8051_top_1.oc8051_ram_top1.bit_select [2], \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_23080_, _23079_, _23078_);
  and (_23081_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _22766_);
  and (_23082_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _22766_);
  nor (_23083_, _23082_, _23081_);
  not (_23084_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23085_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _22766_);
  and (_23086_, _23085_, _23084_);
  and (_23087_, _23086_, _23083_);
  not (_23088_, _23087_);
  not (_23089_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_23090_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_23091_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_23092_, _23091_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_23093_, _23092_, _23090_);
  or (_23094_, _23093_, _23089_);
  not (_23095_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_23096_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand (_23097_, _23096_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_23098_, _23097_, _23095_);
  and (_23099_, _23098_, _23094_);
  not (_23100_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  or (_23101_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_23102_, _23101_, _23091_);
  or (_23103_, _23102_, _23100_);
  not (_23104_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  or (_23105_, _23092_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_23106_, _23105_, _23104_);
  and (_23107_, _23106_, _23103_);
  and (_23108_, _23107_, _23099_);
  or (_23109_, _23101_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  not (_23110_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_23111_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23110_);
  or (_23112_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_23113_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23114_, _23113_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and (_23115_, _23114_, _23112_);
  or (_23116_, _23115_, _23111_);
  nand (_23117_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23110_);
  or (_23118_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_23120_, _23118_, _23116_);
  or (_23121_, _23120_, _23109_);
  and (_23122_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_23123_, _23122_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_23124_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  not (_23126_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand (_23127_, _23122_, _23090_);
  or (_23128_, _23127_, _23126_);
  and (_23129_, _23128_, _23124_);
  and (_23130_, _23129_, _23121_);
  and (_23131_, _23130_, _23108_);
  or (_23132_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_23133_, _23132_, _23120_);
  and (_23134_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_23135_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not (_23137_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_23138_, _23137_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nor (_23139_, _23138_, _23126_);
  nor (_23140_, _23139_, _23135_);
  and (_23141_, _23140_, _23133_);
  not (_23142_, _23141_);
  and (_23143_, _23142_, _23131_);
  nor (_23144_, _23141_, _23131_);
  and (_23145_, _23141_, _23131_);
  nor (_23146_, _23145_, _23144_);
  not (_23147_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_23148_, _23093_, _23147_);
  not (_23149_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_23150_, _23097_, _23149_);
  and (_23151_, _23150_, _23148_);
  not (_23152_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or (_23153_, _23102_, _23152_);
  not (_23154_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or (_23155_, _23105_, _23154_);
  and (_23156_, _23155_, _23153_);
  and (_23157_, _23156_, _23151_);
  or (_23158_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or (_23159_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _23113_);
  and (_23160_, _23159_, _23158_);
  or (_23161_, _23160_, _23111_);
  or (_23163_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_23164_, _23163_, _23161_);
  or (_23165_, _23164_, _23109_);
  not (_23166_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_23167_, _23127_, _23166_);
  nand (_23168_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_23169_, _23168_, _23167_);
  and (_23170_, _23169_, _23165_);
  and (_23171_, _23170_, _23157_);
  or (_23172_, _23164_, _23132_);
  nand (_23173_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or (_23174_, _23138_, _23166_);
  and (_23175_, _23174_, _23173_);
  nand (_23177_, _23175_, _23172_);
  nor (_23178_, _23177_, _23171_);
  not (_23179_, _23177_);
  nor (_23180_, _23179_, _23171_);
  and (_23181_, _23179_, _23171_);
  nor (_23182_, _23181_, _23180_);
  not (_23183_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_23184_, _23093_, _23183_);
  not (_23185_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_23186_, _23097_, _23185_);
  and (_23187_, _23186_, _23184_);
  not (_23188_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  or (_23190_, _23102_, _23188_);
  not (_23191_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or (_23192_, _23105_, _23191_);
  and (_23193_, _23192_, _23190_);
  and (_23194_, _23193_, _23187_);
  or (_23195_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or (_23196_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _23113_);
  and (_23197_, _23196_, _23195_);
  or (_23198_, _23197_, _23111_);
  or (_23199_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_23200_, _23199_, _23198_);
  or (_23201_, _23200_, _23109_);
  not (_23202_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_23203_, _23127_, _23202_);
  nand (_23204_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_23205_, _23204_, _23203_);
  and (_23206_, _23205_, _23201_);
  nand (_23208_, _23206_, _23194_);
  or (_23209_, _23200_, _23132_);
  nand (_23211_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or (_23212_, _23138_, _23202_);
  and (_23213_, _23212_, _23211_);
  and (_23214_, _23213_, _23209_);
  and (_23215_, _23214_, _23208_);
  nand (_23216_, _23213_, _23209_);
  and (_23217_, _23216_, _23208_);
  nor (_23218_, _23216_, _23208_);
  nor (_23219_, _23218_, _23217_);
  not (_23220_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_23221_, _23093_, _23220_);
  not (_23222_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_23223_, _23097_, _23222_);
  and (_23224_, _23223_, _23221_);
  not (_23225_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  or (_23226_, _23102_, _23225_);
  not (_23227_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or (_23228_, _23105_, _23227_);
  and (_23229_, _23228_, _23226_);
  and (_23230_, _23229_, _23224_);
  or (_23231_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or (_23232_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _23113_);
  and (_23233_, _23232_, _23231_);
  or (_23235_, _23233_, _23111_);
  or (_23236_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_23237_, _23236_, _23235_);
  or (_23238_, _23237_, _23109_);
  not (_23239_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_23240_, _23127_, _23239_);
  nand (_23241_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_23242_, _23241_, _23240_);
  and (_23243_, _23242_, _23238_);
  and (_23244_, _23243_, _23230_);
  or (_23245_, _23237_, _23132_);
  nand (_23246_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or (_23247_, _23138_, _23239_);
  and (_23249_, _23247_, _23246_);
  nand (_23250_, _23249_, _23245_);
  and (_23251_, _23250_, _23244_);
  nor (_23252_, _23251_, _23219_);
  nor (_23253_, _23252_, _23215_);
  nor (_23254_, _23253_, _23182_);
  nor (_23256_, _23254_, _23178_);
  and (_23257_, _23253_, _23182_);
  nor (_23258_, _23257_, _23254_);
  not (_23259_, _23258_);
  and (_23260_, _23251_, _23219_);
  nor (_23261_, _23260_, _23252_);
  not (_23262_, _23261_);
  and (_23263_, _23249_, _23245_);
  nor (_23264_, _23263_, _23244_);
  and (_23265_, _23263_, _23244_);
  nor (_23266_, _23265_, _23264_);
  not (_23267_, _23266_);
  not (_23268_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_23269_, _23093_, _23268_);
  not (_23270_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_23271_, _23097_, _23270_);
  and (_23272_, _23271_, _23269_);
  not (_23273_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or (_23274_, _23102_, _23273_);
  not (_23275_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or (_23276_, _23105_, _23275_);
  and (_23277_, _23276_, _23274_);
  and (_23278_, _23277_, _23272_);
  or (_23279_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_23280_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _23113_);
  and (_23281_, _23280_, _23279_);
  or (_23282_, _23281_, _23111_);
  or (_23283_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_23284_, _23283_, _23282_);
  or (_23285_, _23284_, _23109_);
  nand (_23286_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not (_23287_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_23288_, _23127_, _23287_);
  and (_23289_, _23288_, _23286_);
  and (_23290_, _23289_, _23285_);
  and (_23291_, _23290_, _23278_);
  or (_23292_, _23284_, _23132_);
  nand (_23293_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or (_23294_, _23138_, _23287_);
  and (_23295_, _23294_, _23293_);
  and (_23296_, _23295_, _23292_);
  and (_23298_, _23296_, _23291_);
  nor (_23299_, _23296_, _23291_);
  nor (_23301_, _23299_, _23298_);
  not (_23302_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  or (_23303_, _23102_, _23302_);
  not (_23304_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_23305_, _23127_, _23304_);
  and (_23306_, _23305_, _23303_);
  not (_23307_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_23308_, _23093_, _23307_);
  not (_23309_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_23310_, _23097_, _23309_);
  and (_23311_, _23310_, _23308_);
  and (_23312_, _23311_, _23306_);
  or (_23313_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or (_23314_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _23113_);
  and (_23315_, _23314_, _23313_);
  or (_23316_, _23315_, _23111_);
  or (_23317_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_23318_, _23317_, _23316_);
  or (_23320_, _23318_, _23109_);
  nand (_23321_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  not (_23322_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_23323_, _23105_, _23322_);
  and (_23324_, _23323_, _23321_);
  and (_23325_, _23324_, _23320_);
  nand (_23326_, _23325_, _23312_);
  or (_23327_, _23318_, _23132_);
  nand (_23329_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_23330_, _23138_, _23304_);
  and (_23331_, _23330_, _23329_);
  nand (_23332_, _23331_, _23327_);
  and (_23333_, _23332_, _23326_);
  nor (_23334_, _23332_, _23326_);
  nor (_23335_, _23334_, _23333_);
  not (_23336_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_23337_, _23093_, _23336_);
  not (_23338_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_23339_, _23097_, _23338_);
  and (_23340_, _23339_, _23337_);
  not (_23341_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  or (_23342_, _23102_, _23341_);
  not (_23343_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_23344_, _23105_, _23343_);
  and (_23345_, _23344_, _23342_);
  and (_23346_, _23345_, _23340_);
  or (_23347_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or (_23348_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _23113_);
  and (_23349_, _23348_, _23347_);
  or (_23350_, _23349_, _23111_);
  or (_23351_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_23352_, _23351_, _23350_);
  or (_23353_, _23352_, _23109_);
  nand (_23354_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  not (_23355_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_23356_, _23127_, _23355_);
  and (_23357_, _23356_, _23354_);
  and (_23358_, _23357_, _23353_);
  nand (_23359_, _23358_, _23346_);
  or (_23360_, _23352_, _23132_);
  nand (_23361_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_23362_, _23138_, _23355_);
  and (_23363_, _23362_, _23361_);
  nand (_23364_, _23363_, _23360_);
  and (_23365_, _23364_, _23359_);
  nor (_23366_, _23364_, _23359_);
  nor (_23367_, _23366_, _23365_);
  not (_23368_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_23369_, _23093_, _23368_);
  not (_23370_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_23371_, _23097_, _23370_);
  nor (_23372_, _23371_, _23369_);
  not (_23373_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor (_23374_, _23102_, _23373_);
  not (_23375_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_23376_, _23105_, _23375_);
  nor (_23377_, _23376_, _23374_);
  and (_23378_, _23377_, _23372_);
  or (_23379_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or (_23380_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _23113_);
  and (_23381_, _23380_, _23379_);
  or (_23382_, _23381_, _23111_);
  or (_23383_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_23384_, _23383_, _23382_);
  or (_23385_, _23384_, _23109_);
  and (_23386_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  not (_23387_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_23389_, _23127_, _23387_);
  nor (_23390_, _23389_, _23386_);
  and (_23391_, _23390_, _23385_);
  and (_23392_, _23391_, _23378_);
  or (_23393_, _23384_, _23132_);
  nand (_23394_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or (_23395_, _23138_, _23387_);
  and (_23396_, _23395_, _23394_);
  nand (_23397_, _23396_, _23393_);
  and (_23398_, _23397_, _23392_);
  nor (_23399_, _23398_, _23367_);
  and (_23400_, _23363_, _23360_);
  and (_23401_, _23400_, _23359_);
  nor (_23402_, _23401_, _23399_);
  nor (_23403_, _23402_, _23335_);
  and (_23404_, _23331_, _23327_);
  and (_23405_, _23404_, _23326_);
  nor (_23407_, _23405_, _23403_);
  nor (_23408_, _23407_, _23301_);
  and (_23409_, _23407_, _23301_);
  nor (_23411_, _23409_, _23408_);
  and (_23412_, _23402_, _23335_);
  nor (_23413_, _23412_, _23403_);
  not (_23414_, _23413_);
  and (_23415_, _23398_, _23367_);
  nor (_23416_, _23415_, _23399_);
  not (_23417_, _23416_);
  and (_23418_, _23396_, _23393_);
  nor (_23419_, _23418_, _23392_);
  and (_23420_, _23418_, _23392_);
  nor (_23421_, _23420_, _23419_);
  not (_23422_, _23421_);
  nor (_23423_, _23117_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_23424_, _23423_);
  not (_23425_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_23427_, _23425_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_23428_, _23427_, _23160_);
  and (_23429_, _23428_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23430_, _23233_, _23078_);
  and (_23431_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_23432_, _23431_, _23115_);
  not (_23433_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23434_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _23433_);
  nand (_23435_, _23434_, _23197_);
  and (_23436_, _23435_, _23432_);
  and (_23437_, _23436_, _23430_);
  nand (_23438_, _23437_, _23429_);
  not (_23439_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23440_, _23427_, _23315_);
  and (_23441_, _23440_, _23439_);
  nand (_23442_, _23434_, _23349_);
  nand (_23443_, _23431_, _23281_);
  nand (_23444_, _23381_, _23078_);
  and (_23445_, _23444_, _23443_);
  and (_23446_, _23445_, _23442_);
  nand (_23447_, _23446_, _23441_);
  nand (_23448_, _23447_, _23438_);
  nand (_23449_, _23448_, _23117_);
  and (_23450_, _23449_, _23424_);
  and (_23451_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_23452_, _23451_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_23453_, _23452_);
  and (_23454_, _23453_, _23450_);
  and (_23455_, _23453_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_23456_, _23455_, _23454_);
  and (_23457_, _23456_, _23422_);
  and (_23458_, _23457_, _23417_);
  and (_23459_, _23458_, _23414_);
  not (_23460_, _23459_);
  nor (_23461_, _23460_, _23411_);
  nand (_23462_, _23295_, _23292_);
  or (_23463_, _23462_, _23291_);
  and (_23464_, _23462_, _23291_);
  or (_23465_, _23407_, _23464_);
  and (_23466_, _23465_, _23463_);
  or (_23467_, _23466_, _23461_);
  and (_23468_, _23467_, _23267_);
  and (_23469_, _23468_, _23262_);
  and (_23470_, _23469_, _23259_);
  nor (_23471_, _23470_, _23256_);
  nor (_23472_, _23471_, _23146_);
  nor (_23473_, _23472_, _23143_);
  nor (_23474_, _23473_, _23088_);
  not (_23475_, _23474_);
  not (_23476_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_23478_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _22766_);
  and (_23479_, _23478_, _23476_);
  and (_23480_, _23479_, _23083_);
  not (_23481_, _23480_);
  not (_23482_, _23144_);
  not (_23483_, _23146_);
  not (_23484_, _23335_);
  and (_23485_, _23419_, _23367_);
  nor (_23486_, _23485_, _23365_);
  nor (_23487_, _23486_, _23484_);
  nor (_23488_, _23487_, _23333_);
  nor (_23489_, _23488_, _23301_);
  and (_23490_, _23488_, _23301_);
  nor (_23491_, _23490_, _23489_);
  and (_23492_, _23456_, _23421_);
  and (_23493_, _23492_, _23367_);
  and (_23494_, _23486_, _23484_);
  nor (_23495_, _23494_, _23487_);
  and (_23496_, _23495_, _23493_);
  not (_23497_, _23496_);
  nor (_23498_, _23497_, _23491_);
  nor (_23499_, _23488_, _23298_);
  or (_23500_, _23499_, _23299_);
  or (_23501_, _23500_, _23498_);
  and (_23502_, _23501_, _23266_);
  and (_23503_, _23502_, _23219_);
  not (_23505_, _23182_);
  and (_23506_, _23264_, _23219_);
  nor (_23508_, _23506_, _23217_);
  nor (_23509_, _23508_, _23505_);
  and (_23510_, _23508_, _23505_);
  nor (_23511_, _23510_, _23509_);
  and (_23512_, _23511_, _23503_);
  not (_23514_, _23512_);
  nor (_23515_, _23509_, _23180_);
  and (_23516_, _23515_, _23514_);
  or (_23518_, _23516_, _23483_);
  and (_23519_, _23518_, _23482_);
  nor (_23520_, _23519_, _23481_);
  nor (_23521_, _23455_, _23454_);
  not (_23522_, _23208_);
  and (_23523_, _23522_, _23171_);
  not (_23524_, _23523_);
  not (_23525_, _23244_);
  not (_23526_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_23527_, _23082_, _23526_);
  and (_23528_, _23527_, _23479_);
  nor (_23529_, _23359_, _23326_);
  nor (_23530_, _23529_, _23291_);
  and (_23531_, _23530_, _23528_);
  and (_23532_, _23531_, _23525_);
  nor (_23533_, _23532_, _23524_);
  nand (_23534_, _23533_, _23521_);
  not (_23535_, _23533_);
  not (_23536_, _23131_);
  and (_23537_, _23456_, _23536_);
  and (_23538_, _23537_, _23535_);
  not (_23539_, _23528_);
  and (_23540_, _23521_, _23131_);
  or (_23541_, _23540_, _23539_);
  nor (_23542_, _23541_, _23538_);
  and (_23543_, _23542_, _23534_);
  not (_23544_, _23543_);
  nor (_23545_, _23455_, _23450_);
  not (_23546_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_23547_, _23081_, _23546_);
  and (_23548_, _23547_, _23479_);
  nor (_23549_, _23478_, _23085_);
  and (_23550_, _23549_, _23547_);
  not (_23551_, _23550_);
  nor (_23552_, _23551_, _23454_);
  nor (_23553_, _23552_, _23548_);
  nor (_23555_, _23553_, _23545_);
  not (_23556_, _23555_);
  and (_23557_, _23527_, _23086_);
  and (_23558_, _23557_, _23521_);
  not (_23559_, _23558_);
  not (_23560_, _23531_);
  not (_23561_, _23450_);
  and (_23562_, _23081_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_23563_, _23562_, _23549_);
  and (_23564_, _23563_, _23455_);
  and (_23565_, _23564_, _23561_);
  not (_23567_, _23392_);
  and (_23568_, _23562_, _23479_);
  and (_23569_, _23568_, _23567_);
  and (_23570_, _23085_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23571_, _23570_, _23547_);
  and (_23572_, _23571_, _23536_);
  nor (_23574_, _23572_, _23569_);
  not (_23575_, _23574_);
  nor (_23576_, _23575_, _23565_);
  and (_23577_, _23576_, _23560_);
  and (_23578_, _23577_, _23559_);
  and (_23579_, _23549_, _23083_);
  and (_23580_, _23579_, _23456_);
  and (_23581_, _23452_, _23450_);
  and (_23582_, _23547_, _23086_);
  and (_23583_, _23570_, _23527_);
  and (_23584_, _23583_, _23450_);
  nor (_23585_, _23584_, _23582_);
  nor (_23587_, _23585_, _23581_);
  nor (_23588_, _23587_, _23580_);
  and (_23589_, _23588_, _23578_);
  and (_23590_, _23589_, _23556_);
  and (_23591_, _23590_, _23544_);
  not (_23592_, _23591_);
  nor (_23593_, _23592_, _23520_);
  and (_23594_, _23593_, _23475_);
  nor (_23595_, _23594_, _23080_);
  and (_23596_, _23570_, _23083_);
  not (_23597_, _23596_);
  and (_23598_, _23479_, _23526_);
  and (_23599_, _23549_, _23527_);
  nor (_23600_, _23599_, _23598_);
  and (_23601_, _23600_, _23597_);
  and (_23602_, _23562_, _23476_);
  not (_23603_, _23602_);
  and (_23604_, _23547_, _23085_);
  nor (_23605_, _23604_, _23579_);
  and (_23606_, _23605_, _23603_);
  and (_23607_, _23606_, _23601_);
  nor (_23608_, _23607_, _23244_);
  and (_23609_, _23562_, _23086_);
  not (_23610_, _23326_);
  and (_23611_, _23610_, _23291_);
  not (_23612_, _23359_);
  and (_23613_, _23392_, _23612_);
  and (_23614_, _23613_, _23611_);
  or (_23615_, _23614_, _23521_);
  not (_23616_, _23291_);
  and (_23617_, _23567_, _23359_);
  and (_23618_, _23617_, _23326_);
  and (_23619_, _23618_, _23616_);
  or (_23621_, _23619_, _23456_);
  and (_23622_, _23621_, _23615_);
  or (_23623_, _23622_, _23525_);
  nand (_23624_, _23622_, _23525_);
  and (_23625_, _23624_, _23623_);
  and (_23626_, _23625_, _23609_);
  and (_23627_, _23570_, _23562_);
  or (_23628_, _23521_, _23263_);
  or (_23629_, _23456_, _23244_);
  nand (_23630_, _23629_, _23628_);
  nand (_23631_, _23630_, _23627_);
  and (_23632_, _23550_, _23266_);
  and (_23633_, _23583_, _23264_);
  not (_23634_, _23548_);
  nor (_23635_, _23634_, _23265_);
  and (_23636_, _23557_, _23244_);
  or (_23637_, _23636_, _23635_);
  or (_23638_, _23637_, _23633_);
  nor (_23639_, _23638_, _23632_);
  nand (_23640_, _23639_, _23631_);
  or (_23641_, _23640_, _23626_);
  or (_23642_, _23641_, _23608_);
  and (_23643_, _23642_, _22948_);
  and (_23644_, _23078_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23645_, _23233_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23646_, _23645_, _23644_);
  or (_23647_, _23646_, _23643_);
  or (_23648_, _23647_, _23595_);
  and (_23649_, _23648_, _22946_);
  and (_23651_, _23649_, _23077_);
  not (_23652_, _23077_);
  and (_23653_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or (_02714_, _23653_, _23651_);
  nor (_23654_, _23067_, _22947_);
  and (_23655_, _23654_, _23039_);
  and (_23656_, _23655_, _23021_);
  nor (_23657_, _23053_, _22949_);
  not (_23658_, _23657_);
  and (_23660_, _23658_, _22946_);
  nor (_23661_, _23660_, _23071_);
  and (_23662_, _23035_, _22943_);
  and (_23663_, _23662_, _22946_);
  and (_23664_, _23663_, _23661_);
  and (_23665_, _23664_, _23656_);
  nand (_23666_, _23431_, _23079_);
  nor (_23667_, _23666_, _23594_);
  nand (_23668_, _23431_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_23669_, _23115_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23670_, _23669_, _23668_);
  nor (_23671_, _23607_, _23131_);
  not (_23672_, _23671_);
  and (_23673_, _23614_, _23244_);
  and (_23674_, _23673_, _23523_);
  nor (_23675_, _23674_, _23521_);
  nand (_23676_, _23619_, _23525_);
  or (_23677_, _23676_, _23522_);
  or (_23678_, _23677_, _23171_);
  and (_23679_, _23678_, _23521_);
  nor (_23680_, _23679_, _23675_);
  or (_23681_, _23680_, _23131_);
  nand (_23682_, _23680_, _23131_);
  nand (_23683_, _23682_, _23681_);
  nand (_23684_, _23683_, _23609_);
  and (_23686_, _23456_, _23141_);
  not (_23687_, _23686_);
  not (_23688_, _23627_);
  nor (_23689_, _23688_, _23540_);
  and (_23690_, _23689_, _23687_);
  and (_23691_, _23550_, _23146_);
  and (_23692_, _23583_, _23144_);
  nor (_23693_, _23634_, _23145_);
  and (_23694_, _23557_, _23131_);
  or (_23695_, _23694_, _23693_);
  or (_23696_, _23695_, _23692_);
  nor (_23697_, _23696_, _23691_);
  not (_23699_, _23697_);
  nor (_23700_, _23699_, _23690_);
  and (_23701_, _23700_, _23684_);
  and (_23702_, _23701_, _23672_);
  nor (_23704_, _23702_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  or (_23705_, _23704_, _23670_);
  or (_23706_, _23705_, _23667_);
  and (_23707_, _23706_, _22946_);
  and (_23708_, _23707_, _23665_);
  not (_23709_, _23665_);
  and (_23710_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or (_27079_, _23710_, _23708_);
  not (_23711_, _23594_);
  and (_23712_, _23439_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23713_, _23712_, _23431_);
  and (_23714_, _23713_, _23711_);
  and (_23715_, _23627_, _23462_);
  nor (_23716_, _23618_, _23616_);
  or (_23717_, _23716_, _23621_);
  nand (_23718_, _23529_, _23392_);
  and (_23719_, _23718_, _23616_);
  or (_23720_, _23719_, _23614_);
  nand (_23721_, _23720_, _23456_);
  nand (_23722_, _23721_, _23717_);
  and (_23724_, _23722_, _23609_);
  nor (_23725_, _23724_, _23715_);
  nor (_23726_, _23607_, _23291_);
  not (_23727_, _23726_);
  and (_23728_, _23550_, _23301_);
  not (_23729_, _23728_);
  nor (_23730_, _23634_, _23298_);
  not (_23731_, _23730_);
  and (_23732_, _23583_, _23299_);
  and (_23733_, _23557_, _23291_);
  nor (_23734_, _23733_, _23732_);
  and (_23735_, _23734_, _23731_);
  and (_23736_, _23735_, _23729_);
  and (_23737_, _23736_, _23727_);
  nand (_23738_, _23737_, _23725_);
  and (_23739_, _23738_, _22948_);
  and (_23740_, _23712_, _23425_);
  and (_23741_, _23712_, _23433_);
  or (_23742_, _23741_, _23079_);
  or (_23743_, _23742_, _23740_);
  and (_23744_, _23743_, _23281_);
  or (_23745_, _23744_, _23739_);
  or (_23746_, _23745_, _23714_);
  and (_23747_, _23746_, _22946_);
  and (_23748_, _23747_, _23077_);
  and (_23749_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  or (_09923_, _23749_, _23748_);
  nor (_23750_, _23020_, _22947_);
  and (_23751_, _23750_, _22986_);
  and (_23752_, _23751_, _23655_);
  and (_23753_, _23034_, _22943_);
  and (_23754_, _23753_, _23072_);
  and (_23755_, _23754_, _23752_);
  and (_23756_, _23712_, _23078_);
  nand (_23757_, _23756_, _23594_);
  nor (_23758_, _23551_, _23419_);
  nor (_23759_, _23758_, _23548_);
  or (_23760_, _23759_, _23420_);
  and (_23761_, _23583_, _23419_);
  and (_23762_, _23557_, _23392_);
  nor (_23764_, _23762_, _23761_);
  and (_23765_, _23627_, _23397_);
  and (_23766_, _23609_, _23392_);
  nor (_23767_, _23766_, _23765_);
  nor (_23768_, _23607_, _23392_);
  not (_23769_, _23768_);
  and (_23770_, _23769_, _23767_);
  and (_23771_, _23770_, _23764_);
  and (_23772_, _23771_, _23760_);
  nand (_23773_, _23772_, _22948_);
  or (_23774_, _23381_, _22948_);
  and (_23775_, _23774_, _23773_);
  or (_23776_, _23775_, _23756_);
  and (_23777_, _23776_, _23757_);
  and (_23778_, _23777_, _22946_);
  and (_23779_, _23778_, _23755_);
  not (_23780_, _23755_);
  and (_23781_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or (_13798_, _23781_, _23779_);
  nor (_23782_, _23750_, _22986_);
  nor (_23783_, _23654_, _23040_);
  and (_23784_, _23783_, _23782_);
  and (_23785_, _23071_, _23052_);
  nor (_23786_, _23034_, _22949_);
  and (_23787_, _23786_, _22946_);
  and (_23788_, _23787_, _22944_);
  and (_23789_, _23788_, _23785_);
  and (_23790_, _23789_, _23784_);
  nand (_23791_, _23712_, _23427_);
  nor (_23792_, _23791_, _23594_);
  and (_23793_, _23627_, _23332_);
  not (_23794_, _23613_);
  or (_23795_, _23794_, _23521_);
  not (_23796_, _23617_);
  or (_23797_, _23796_, _23456_);
  and (_23798_, _23797_, _23795_);
  nand (_23799_, _23798_, _23610_);
  or (_23800_, _23798_, _23610_);
  and (_23801_, _23800_, _23609_);
  and (_23802_, _23801_, _23799_);
  nor (_23803_, _23802_, _23793_);
  and (_23804_, _23550_, _23335_);
  nor (_23805_, _23634_, _23334_);
  or (_23806_, _23805_, _23804_);
  not (_23807_, _23806_);
  and (_23808_, _23583_, _23333_);
  and (_23809_, _23557_, _23610_);
  nor (_23810_, _23809_, _23808_);
  and (_23811_, _23810_, _23807_);
  nor (_23812_, _23607_, _23610_);
  not (_23813_, _23812_);
  and (_23814_, _23813_, _23811_);
  nand (_23816_, _23814_, _23803_);
  and (_23817_, _23816_, _22948_);
  or (_23818_, _23713_, _23079_);
  or (_23820_, _23818_, _23741_);
  and (_23821_, _23820_, _23315_);
  or (_23822_, _23821_, _23817_);
  or (_23823_, _23822_, _23792_);
  and (_23824_, _23823_, _22946_);
  and (_23825_, _23824_, _23790_);
  not (_23827_, _23790_);
  and (_23828_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  or (_16236_, _23828_, _23825_);
  and (_23829_, _23790_, _23649_);
  and (_23830_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  or (_16455_, _23830_, _23829_);
  and (_23831_, _23790_, _23747_);
  and (_23832_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  or (_22627_, _23832_, _23831_);
  and (_23833_, _23754_, _23656_);
  and (_23834_, _23833_, _23824_);
  not (_23835_, _23833_);
  and (_23836_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_22643_, _23836_, _23834_);
  not (_23837_, _22767_);
  not (_23838_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_23839_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_23840_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_23841_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_23842_, _23841_, _23840_);
  and (_23843_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_23844_, _23841_, _23840_);
  and (_23845_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_23846_, _23841_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_23847_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_23848_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_23849_, _23848_, _23840_);
  and (_23850_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_23851_, _23850_, _23847_);
  nor (_23852_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_23853_, _23852_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_23854_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  not (_23855_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_23856_, _23855_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_23857_, _23856_, _23840_);
  and (_23858_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_23859_, _23858_, _23854_);
  nand (_23860_, _23859_, _23851_);
  or (_23861_, _23860_, _23845_);
  nor (_23862_, _23861_, _23843_);
  and (_23863_, _23862_, _23839_);
  and (_23864_, _23863_, _23838_);
  nor (_23865_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _23838_);
  nor (_23866_, _23865_, _23864_);
  or (_23867_, _23866_, _23837_);
  or (_23868_, _22767_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_23869_, _23868_, _22762_);
  and (_26864_[1], _23869_, _23867_);
  nand (_23870_, _23712_, _23434_);
  nor (_23871_, _23870_, _23594_);
  and (_23872_, _23627_, _23364_);
  nor (_23873_, _23617_, _23613_);
  nand (_23874_, _23873_, _23456_);
  or (_23875_, _23873_, _23456_);
  and (_23876_, _23875_, _23609_);
  and (_23877_, _23876_, _23874_);
  nor (_23878_, _23877_, _23872_);
  nor (_23879_, _23607_, _23612_);
  not (_23880_, _23879_);
  and (_23881_, _23550_, _23367_);
  not (_23882_, _23881_);
  nor (_23883_, _23634_, _23366_);
  not (_23884_, _23883_);
  and (_23885_, _23583_, _23365_);
  and (_23886_, _23557_, _23612_);
  nor (_23887_, _23886_, _23885_);
  and (_23888_, _23887_, _23884_);
  and (_23889_, _23888_, _23882_);
  and (_23890_, _23889_, _23880_);
  nand (_23892_, _23890_, _23878_);
  and (_23893_, _23892_, _22948_);
  or (_23894_, _23740_, _23818_);
  and (_23895_, _23894_, _23349_);
  or (_23896_, _23895_, _23893_);
  or (_23897_, _23896_, _23871_);
  and (_23898_, _23897_, _22946_);
  and (_23899_, _23898_, _23833_);
  and (_23900_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_22722_, _23900_, _23899_);
  and (_23901_, _23750_, _22985_);
  and (_23902_, _23654_, _23040_);
  and (_23903_, _23902_, _23901_);
  not (_23904_, _23070_);
  and (_23905_, _23660_, _23904_);
  and (_23906_, _23905_, _23788_);
  and (_23907_, _23906_, _23903_);
  and (_23908_, _23907_, _23747_);
  not (_23909_, _23907_);
  and (_23910_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_22746_, _23910_, _23908_);
  and (_23911_, _23783_, _23751_);
  and (_23912_, _23911_, _23789_);
  nand (_23913_, _23434_, _23079_);
  nor (_23914_, _23913_, _23594_);
  and (_23915_, _23521_, _23522_);
  and (_23916_, _23456_, _23214_);
  or (_23917_, _23916_, _23688_);
  nor (_23918_, _23917_, _23915_);
  or (_23919_, _23676_, _23456_);
  nand (_23920_, _23673_, _23456_);
  and (_23921_, _23920_, _23919_);
  and (_23922_, _23921_, _23522_);
  or (_23923_, _23921_, _23522_);
  nand (_23924_, _23923_, _23609_);
  nor (_23925_, _23924_, _23922_);
  nor (_23926_, _23925_, _23918_);
  and (_23927_, _23550_, _23219_);
  and (_23929_, _23583_, _23217_);
  nor (_23930_, _23634_, _23218_);
  and (_23932_, _23557_, _23522_);
  or (_23933_, _23932_, _23930_);
  or (_23934_, _23933_, _23929_);
  nor (_23935_, _23934_, _23927_);
  nor (_23936_, _23607_, _23522_);
  not (_23937_, _23936_);
  and (_23938_, _23937_, _23935_);
  nand (_23939_, _23938_, _23926_);
  and (_23940_, _23939_, _22948_);
  nand (_23941_, _23434_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_23942_, _23197_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23943_, _23942_, _23941_);
  or (_23944_, _23943_, _23940_);
  or (_23945_, _23944_, _23914_);
  and (_23946_, _23945_, _22946_);
  and (_23947_, _23946_, _23912_);
  not (_23948_, _23912_);
  and (_23949_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or (_22757_, _23949_, _23947_);
  not (_23950_, _22768_);
  nor (_23951_, _23848_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_23952_, _23951_, _23950_);
  nor (_23953_, _23952_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_23954_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  not (_23955_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor (_23956_, _23953_, _23955_);
  or (_23957_, _23956_, _23954_);
  and (_26904_[31], _23957_, _22762_);
  and (_23958_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_23959_, _23958_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  or (_23960_, _23959_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_26902_[3], _23960_, _22762_);
  or (_23961_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  nand (_23962_, _23953_, _23955_);
  and (_23963_, _23962_, _22762_);
  and (_26903_[31], _23963_, _23961_);
  and (_26900_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _22762_);
  not (_23964_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_23965_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor (_23966_, _23965_, _23964_);
  and (_23967_, _23965_, _23964_);
  nor (_23968_, _23967_, _23966_);
  not (_23969_, _23968_);
  and (_23970_, _23969_, _26902_[3]);
  nor (_23971_, _23966_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_23972_, _23966_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_23973_, _23972_, _23971_);
  nor (_23974_, _23958_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_23975_, _23974_, _23959_);
  or (_23976_, _23975_, _23965_);
  and (_23977_, _23976_, _23973_);
  and (_26901_, _23977_, _23970_);
  not (_23978_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_23979_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _23978_);
  and (_23980_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_23981_, _23980_, _23979_);
  and (_26899_[7], _23981_, _22762_);
  and (_23982_, _23907_, _23898_);
  and (_23983_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_24175_, _23983_, _23982_);
  and (_23984_, _23755_, _23649_);
  and (_23985_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or (_24247_, _23985_, _23984_);
  and (_23986_, _23751_, _23068_);
  and (_23987_, _23986_, _23906_);
  and (_23988_, _23987_, _23747_);
  not (_23989_, _23987_);
  and (_23990_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or (_24383_, _23990_, _23988_);
  and (_23991_, _23902_, _23021_);
  and (_23992_, _23991_, _23906_);
  and (_23993_, _23992_, _23778_);
  not (_23994_, _23992_);
  and (_23995_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_26943_, _23995_, _23993_);
  and (_23997_, _23946_, _23907_);
  and (_23998_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_26940_, _23998_, _23997_);
  and (_24000_, _23907_, _23707_);
  and (_24001_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_26941_, _24001_, _24000_);
  and (_24003_, _23907_, _23649_);
  and (_24004_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_26939_, _24004_, _24003_);
  and (_24005_, _23902_, _23782_);
  and (_24006_, _24005_, _23906_);
  and (_24007_, _24006_, _23707_);
  not (_24008_, _24006_);
  and (_24009_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or (_26938_, _24009_, _24007_);
  and (_24010_, _23783_, _23021_);
  and (_24011_, _24010_, _23789_);
  and (_24012_, _24011_, _23707_);
  not (_24013_, _24011_);
  and (_24014_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_27264_, _24014_, _24012_);
  nand (_24015_, _23427_, _23079_);
  nor (_24016_, _24015_, _23594_);
  nor (_24017_, _23607_, _23171_);
  and (_24018_, _23677_, _23171_);
  not (_24019_, _24018_);
  and (_24020_, _24019_, _23679_);
  and (_24021_, _23673_, _23522_);
  nor (_24022_, _24021_, _23171_);
  nor (_24023_, _24022_, _23674_);
  nor (_24024_, _24023_, _23521_);
  or (_24025_, _24024_, _24020_);
  nand (_24026_, _24025_, _23609_);
  and (_24027_, _23456_, _23177_);
  not (_24028_, _23171_);
  and (_24029_, _23521_, _24028_);
  nor (_24030_, _24029_, _24027_);
  nor (_24031_, _24030_, _23688_);
  not (_24032_, _24031_);
  and (_24033_, _23550_, _23182_);
  nor (_24034_, _23634_, _23181_);
  or (_24035_, _24034_, _24033_);
  not (_24036_, _24035_);
  and (_24037_, _23583_, _23180_);
  and (_24038_, _23557_, _23171_);
  nor (_24039_, _24038_, _24037_);
  and (_24040_, _24039_, _24036_);
  and (_24041_, _24040_, _24032_);
  nand (_24042_, _24041_, _24026_);
  or (_24043_, _24042_, _24017_);
  and (_24044_, _24043_, _22948_);
  nand (_24045_, _23427_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_24046_, _23160_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_24047_, _24046_, _24045_);
  or (_24048_, _24047_, _24044_);
  or (_24049_, _24048_, _24016_);
  and (_24050_, _24049_, _22946_);
  and (_24051_, _24050_, _24011_);
  and (_24052_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_27263_, _24052_, _24051_);
  and (_24053_, _23833_, _23649_);
  and (_24054_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_27064_, _24054_, _24053_);
  and (_24055_, _23833_, _23747_);
  and (_24056_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_27063_, _24056_, _24055_);
  and (_24057_, _23912_, _23747_);
  and (_24058_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  or (_27267_, _24058_, _24057_);
  and (_24059_, _23912_, _23824_);
  and (_24060_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  or (_27266_, _24060_, _24059_);
  and (_24061_, _23912_, _23898_);
  and (_24062_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or (_27265_, _24062_, _24061_);
  and (_24063_, _23052_, _22970_);
  and (_24064_, _24063_, _23753_);
  not (_24065_, _23018_);
  and (_24066_, _23065_, _22983_);
  and (_24067_, _24066_, _24065_);
  nor (_24068_, _22909_, _22906_);
  and (_24069_, _24068_, _22948_);
  not (_24070_, _24069_);
  nor (_24071_, _24070_, _23002_);
  and (_24072_, _24071_, _24067_);
  and (_24073_, _24072_, _24064_);
  or (_24074_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_24075_, _24074_, _22762_);
  and (_24076_, _24067_, _23003_);
  and (_24077_, _24064_, _24069_);
  and (_24078_, _24077_, _24076_);
  not (_24079_, _24078_);
  or (_24080_, _24079_, _23738_);
  and (_26382_, _24080_, _24075_);
  and (_24081_, _24010_, _23754_);
  and (_24082_, _24081_, _23824_);
  not (_24083_, _24081_);
  and (_24084_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_27052_, _24084_, _24082_);
  and (_24085_, _23901_, _23783_);
  and (_24086_, _24085_, _23789_);
  and (_24087_, _24086_, _23707_);
  not (_24088_, _24086_);
  and (_24089_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_27257_, _24089_, _24087_);
  and (_24090_, _24011_, _23898_);
  and (_24092_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_27259_, _24092_, _24090_);
  and (_24093_, _24081_, _23898_);
  and (_24094_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_27051_, _24094_, _24093_);
  nor (_24095_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_24096_, _24095_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_26907_, _24096_, _22762_);
  and (_24098_, _26900_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_26906_, _24098_, _26907_);
  and (_24100_, _24011_, _23778_);
  and (_24101_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_27258_, _24101_, _24100_);
  and (_24102_, _24081_, _23778_);
  and (_24103_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_27050_, _24103_, _24102_);
  not (_24104_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_24105_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , _24104_);
  and (_26905_, _24105_, _22762_);
  and (_24107_, _24011_, _23649_);
  and (_24108_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_27262_, _24108_, _24107_);
  and (_24109_, _24011_, _23747_);
  and (_24110_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_27261_, _24110_, _24109_);
  and (_24111_, _24011_, _23824_);
  and (_24112_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_27260_, _24112_, _24111_);
  and (_24113_, _24081_, _23946_);
  and (_24114_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_27055_, _24114_, _24113_);
  and (_24115_, _24081_, _23649_);
  and (_24116_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_27054_, _24116_, _24115_);
  nor (_24117_, _23018_, _22983_);
  and (_24118_, _24117_, _23065_);
  and (_24119_, _24118_, _24071_);
  and (_24120_, _24119_, _24064_);
  and (_24121_, _24120_, _22762_);
  and (_24122_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not (_24123_, _23065_);
  and (_24124_, _24065_, _22983_);
  and (_24125_, _24124_, _24123_);
  and (_24126_, _24125_, _24071_);
  and (_24127_, _24126_, _24064_);
  not (_24128_, _24127_);
  or (_24129_, _24128_, _23892_);
  not (_24130_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not (_24131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_24132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _24131_);
  not (_24134_, _24132_);
  not (_24135_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_24136_, t1_i);
  and (_24137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _24136_);
  nor (_24138_, _24137_, _24135_);
  not (_24139_, _24138_);
  not (_24140_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_24141_, _24140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nor (_24142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_24143_, _24142_);
  and (_24144_, _24143_, _24141_);
  and (_24145_, _24144_, _24139_);
  not (_24146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand (_24147_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_24148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_24149_, _24148_, _24147_);
  nor (_24150_, _24149_, _24146_);
  and (_24151_, _24150_, _24145_);
  and (_24152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_24153_, _24152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_24154_, _24153_, _24151_);
  nor (_24155_, _24154_, _24134_);
  not (_24156_, _24155_);
  not (_24157_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_24158_, _24151_, _24131_);
  nor (_24159_, _24158_, _24132_);
  nor (_24160_, _24159_, _24157_);
  and (_24161_, _24160_, _24156_);
  nor (_24162_, _24161_, _24130_);
  and (_24163_, _24161_, _24130_);
  or (_24164_, _24163_, _24162_);
  or (_24165_, _24164_, _24127_);
  nor (_24166_, _24120_, rst);
  and (_24167_, _24166_, _24165_);
  and (_24168_, _24167_, _24129_);
  or (_00740_, _24168_, _24122_);
  and (_24169_, _24081_, _23747_);
  and (_24170_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_27053_, _24170_, _24169_);
  not (_24171_, _24120_);
  or (_24172_, _24171_, _23642_);
  and (_24173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_24174_, _24173_, _24127_);
  nor (_24176_, _24174_, _24146_);
  not (_24177_, _24145_);
  nor (_24178_, _24149_, _24177_);
  or (_24179_, _24178_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_24180_, _24173_, _24151_);
  and (_24181_, _24180_, _24179_);
  not (_24182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_24184_, _24182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_24185_, _24184_, _24154_);
  and (_24186_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_24187_, _24186_, _24181_);
  nor (_24188_, _24187_, _24127_);
  or (_24189_, _24188_, _24176_);
  or (_24190_, _24189_, _24120_);
  and (_24191_, _24190_, _22762_);
  and (_00832_, _24191_, _24172_);
  and (_24192_, _24086_, _23946_);
  and (_24193_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_27255_, _24193_, _24192_);
  and (_24194_, _24085_, _23754_);
  and (_24195_, _24194_, _23747_);
  not (_24196_, _24194_);
  and (_24197_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_27048_, _24197_, _24195_);
  and (_24198_, _24194_, _23649_);
  and (_24199_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_27049_, _24199_, _24198_);
  and (_24201_, _23788_, _23661_);
  and (_24203_, _24201_, _23991_);
  not (_24204_, _24203_);
  and (_24206_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  and (_24207_, _24203_, _23747_);
  or (_27248_, _24207_, _24206_);
  and (_01412_, t1_i, _22762_);
  and (_24208_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  and (_24209_, _24203_, _23824_);
  or (_27247_, _24209_, _24208_);
  and (_24210_, _23824_, _23077_);
  and (_24211_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or (_27214_, _24211_, _24210_);
  and (_24212_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  and (_24213_, _24203_, _23707_);
  or (_01716_, _24213_, _24212_);
  and (_24214_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  and (_24215_, _24203_, _24050_);
  or (_27250_, _24215_, _24214_);
  and (_24216_, _24194_, _23707_);
  and (_24217_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_01953_, _24217_, _24216_);
  and (_24218_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  and (_24219_, _24203_, _23946_);
  or (_27249_, _24219_, _24218_);
  and (_24220_, _24194_, _24050_);
  and (_24221_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_02060_, _24221_, _24220_);
  and (_24222_, _24201_, _23903_);
  not (_24223_, _24222_);
  and (_24224_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  and (_24225_, _24222_, _23946_);
  or (_02437_, _24225_, _24224_);
  and (_24226_, _23784_, _23754_);
  and (_24228_, _24226_, _23707_);
  not (_24229_, _24226_);
  and (_24230_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or (_02582_, _24230_, _24228_);
  and (_24231_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_24232_, _24127_, _23702_);
  and (_24234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_24235_, _24234_, _24150_);
  and (_24236_, _24235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_24237_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_24238_, _24237_, _24236_);
  and (_24239_, _24238_, _24153_);
  and (_24240_, _24145_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_24241_, _24240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_24242_, _24241_, _24239_);
  and (_24243_, _24242_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_24244_, _24242_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_24245_, _24244_, _24132_);
  nor (_24246_, _24245_, _24243_);
  and (_24248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_24249_, _24236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_24250_, _24249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_24251_, _24250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_24252_, _24251_, _24145_);
  and (_24253_, _24252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_24254_, _24253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_24255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_24256_, _24255_);
  and (_24257_, _24253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_24258_, _24257_, _24256_);
  and (_24259_, _24258_, _24254_);
  or (_24260_, _24259_, _24248_);
  or (_24261_, _24260_, _24246_);
  or (_24262_, _24261_, _24127_);
  and (_24263_, _24262_, _24166_);
  and (_24264_, _24263_, _24232_);
  or (_02663_, _24264_, _24231_);
  and (_24265_, _24226_, _24050_);
  and (_24266_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or (_02867_, _24266_, _24265_);
  and (_24267_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  and (_24268_, _24203_, _23778_);
  or (_02903_, _24268_, _24267_);
  and (_24269_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  and (_24270_, _24222_, _23707_);
  or (_03083_, _24270_, _24269_);
  and (_24271_, _24194_, _23778_);
  and (_24272_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_03542_, _24272_, _24271_);
  and (_24273_, _24194_, _23898_);
  and (_24274_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_27046_, _24274_, _24273_);
  and (_24275_, _23902_, _23751_);
  and (_24276_, _24275_, _24201_);
  not (_24277_, _24276_);
  and (_24279_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and (_24280_, _24276_, _23824_);
  or (_03788_, _24280_, _24279_);
  and (_24282_, _23782_, _23655_);
  and (_24283_, _24282_, _23076_);
  and (_24284_, _24283_, _23824_);
  not (_24285_, _24283_);
  and (_24286_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  or (_03822_, _24286_, _24284_);
  and (_24287_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and (_24288_, _24276_, _23898_);
  or (_03855_, _24288_, _24287_);
  not (_24289_, _22983_);
  and (_24290_, _23018_, _24289_);
  and (_24291_, _24290_, _23065_);
  and (_24292_, _24291_, _24071_);
  and (_24293_, _24292_, _24064_);
  not (_24294_, _24293_);
  and (_24295_, _23018_, _22983_);
  and (_24296_, _24295_, _24123_);
  and (_24297_, _24296_, _24071_);
  and (_24299_, _24297_, _24064_);
  and (_24300_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_24301_, _24300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_24302_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_24303_, _24302_, _22762_);
  and (_24304_, _24303_, _24301_);
  not (_24305_, _24300_);
  and (_24307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_24308_, _24307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_24309_, _24308_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_24310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_24312_, _24310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_24313_, _24312_, _24309_);
  and (_24315_, _24313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_24316_, _24315_, _24305_);
  nand (_24317_, _24316_, _24304_);
  nor (_24318_, _24317_, _24299_);
  and (_04338_, _24318_, _24294_);
  and (_24319_, _24226_, _23778_);
  and (_24320_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or (_04361_, _24320_, _24319_);
  and (_24322_, _24226_, _23898_);
  and (_24323_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  or (_04416_, _24323_, _24322_);
  and (_24324_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and (_24325_, _24276_, _23946_);
  or (_04519_, _24325_, _24324_);
  and (_24326_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and (_24328_, _24276_, _23649_);
  or (_04742_, _24328_, _24326_);
  and (_24329_, _23782_, _23068_);
  and (_24331_, _24329_, _23754_);
  and (_24332_, _24331_, _23778_);
  not (_24333_, _24331_);
  and (_24334_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_04802_, _24334_, _24332_);
  and (_24335_, _23898_, _23077_);
  and (_24336_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or (_04851_, _24336_, _24335_);
  and (_24337_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not (_24338_, _24337_);
  nand (_24339_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_24340_, _24339_, _24338_);
  nand (_24341_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_24342_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_24343_, _24342_, _24341_);
  nand (_24344_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_24345_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_24346_, _24345_, _24344_);
  and (_24347_, _24346_, _24343_);
  and (_24348_, _24347_, _24340_);
  or (_24349_, _24348_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_24350_, _24349_, _23838_);
  nor (_24351_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _23838_);
  or (_24352_, _24351_, _24350_);
  nor (_26860_[3], _24352_, rst);
  and (_24353_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and (_24354_, _24276_, _23707_);
  or (_05258_, _24354_, _24353_);
  and (_24356_, _23785_, _23075_);
  and (_24358_, _24356_, _24282_);
  and (_24359_, _24358_, _23824_);
  not (_24360_, _24358_);
  and (_24361_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  or (_05587_, _24361_, _24359_);
  and (_24362_, _24226_, _23747_);
  and (_24363_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  or (_27045_, _24363_, _24362_);
  and (_24364_, _24358_, _23898_);
  and (_24365_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  or (_05673_, _24365_, _24364_);
  and (_24366_, _24226_, _23649_);
  and (_24367_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or (_05825_, _24367_, _24366_);
  and (_24368_, _24358_, _23778_);
  and (_24369_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  or (_05902_, _24369_, _24368_);
  and (_24370_, _23905_, _23075_);
  and (_24371_, _24370_, _23991_);
  and (_24372_, _24371_, _23707_);
  not (_24373_, _24371_);
  and (_24374_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_06170_, _24374_, _24372_);
  and (_24375_, _24370_, _23784_);
  and (_24376_, _24375_, _23778_);
  not (_24377_, _24375_);
  and (_24378_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_06542_, _24378_, _24376_);
  and (_24379_, _24375_, _23824_);
  and (_24380_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_06585_, _24380_, _24379_);
  and (_24381_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_24382_, _22767_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_24384_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_24385_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_24386_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_24388_, _24386_, _24385_);
  and (_24389_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_24391_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_24392_, _24391_, _24389_);
  and (_24393_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_24394_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_24396_, _24394_, _24393_);
  and (_24397_, _24396_, _24392_);
  and (_24399_, _24397_, _24388_);
  nor (_24400_, _24399_, _24384_);
  and (_24401_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  nor (_24402_, _24401_, _24400_);
  and (_24403_, _24402_, _22769_);
  not (_24404_, _24403_);
  not (_24405_, _22765_);
  nor (_24406_, _22768_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_24407_, _24406_, _24405_);
  and (_24408_, _24407_, _24404_);
  not (_24409_, _22769_);
  nor (_24411_, _23866_, _24409_);
  not (_24412_, _24411_);
  nor (_24414_, _22768_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_24415_, _24414_, _24405_);
  and (_24417_, _24415_, _24412_);
  and (_24418_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_24420_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_24421_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_24422_, _24421_, _24420_);
  and (_24424_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_24425_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_24426_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_24427_, _24426_, _24425_);
  or (_24428_, _24427_, _24424_);
  or (_24429_, _24428_, _24422_);
  or (_24430_, _24429_, _24418_);
  nand (_24431_, _24430_, _23839_);
  nand (_24432_, _24431_, _23838_);
  nor (_24434_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _23838_);
  not (_24435_, _24434_);
  and (_24436_, _24435_, _24432_);
  or (_24437_, _24436_, _24409_);
  nor (_24438_, _22768_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_24439_, _24438_, _24405_);
  and (_24440_, _24439_, _24437_);
  and (_24441_, _24352_, _22769_);
  not (_24442_, _24441_);
  nor (_24443_, _22768_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_24444_, _24443_, _24405_);
  and (_24445_, _24444_, _24442_);
  nor (_24446_, _24445_, _24440_);
  and (_24447_, _24446_, _24417_);
  and (_24448_, _24447_, _24408_);
  and (_24450_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_24451_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_24452_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_24453_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_24454_, _24453_, _24452_);
  and (_24455_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_24456_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_24457_, _24456_, _24455_);
  nand (_24458_, _24457_, _24454_);
  or (_24459_, _24458_, _24451_);
  nor (_24460_, _24459_, _24450_);
  and (_24461_, _24460_, _23839_);
  and (_24462_, _24461_, _23838_);
  nor (_24463_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _23838_);
  nor (_24464_, _24463_, _24462_);
  nor (_24466_, _24464_, _24409_);
  not (_24467_, _24466_);
  nor (_24469_, _22768_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_24470_, _24469_, _24405_);
  nand (_24471_, _24470_, _24467_);
  nand (_24472_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand (_24473_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_24474_, _24473_, _24472_);
  nand (_24475_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nand (_24476_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_24477_, _24476_, _24475_);
  and (_24478_, _24477_, _24474_);
  and (_24479_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_24480_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_24481_, _24480_, _24479_);
  and (_24482_, _24481_, _24478_);
  or (_24483_, _24482_, _24384_);
  and (_24484_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_24485_, _24484_);
  and (_24486_, _24485_, _24483_);
  nand (_24487_, _24486_, _22769_);
  nor (_24488_, _22768_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_24489_, _24488_, _24405_);
  and (_24490_, _24489_, _24487_);
  and (_24491_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_24492_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_24493_, _24492_, _24491_);
  nand (_24494_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nand (_24495_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_24497_, _24495_, _24494_);
  nand (_24498_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_24500_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_24501_, _24500_, _24498_);
  and (_24503_, _24501_, _24497_);
  and (_24504_, _24503_, _24493_);
  or (_24505_, _24504_, _24384_);
  and (_24506_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_24507_, _24506_);
  and (_24508_, _24507_, _24505_);
  nand (_24509_, _24508_, _22769_);
  nor (_24510_, _22768_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_24511_, _24510_, _24405_);
  and (_24512_, _24511_, _24509_);
  not (_24513_, _24512_);
  nor (_24514_, _24513_, _24490_);
  nor (_24515_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_24516_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_24517_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_24518_, _24517_, _24516_);
  and (_24519_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_24520_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_24521_, _24520_, _24519_);
  and (_24522_, _24521_, _24518_);
  and (_24523_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_24524_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_24525_, _24524_, _24523_);
  nand (_24526_, _24525_, _24522_);
  nand (_24527_, _24526_, _24515_);
  and (_24528_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_24529_, _24528_);
  and (_24530_, _24529_, _24527_);
  nand (_24531_, _24530_, _22769_);
  nor (_24532_, _22768_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_24533_, _24532_, _24405_);
  and (_24534_, _24533_, _24531_);
  and (_24535_, _24534_, _24514_);
  and (_24536_, _24535_, _24471_);
  and (_24537_, _24536_, _24448_);
  and (_24538_, _24470_, _24467_);
  and (_24539_, _24513_, _24490_);
  and (_24540_, _24539_, _24534_);
  and (_24541_, _24540_, _24538_);
  and (_24542_, _24541_, _24448_);
  nor (_24543_, _24542_, _24537_);
  not (_24544_, _24534_);
  and (_24545_, _24544_, _24514_);
  and (_24546_, _24545_, _24538_);
  and (_24548_, _24546_, _24448_);
  not (_24549_, _24548_);
  and (_24550_, _24549_, _24543_);
  and (_24552_, _24545_, _24471_);
  not (_24553_, _24445_);
  and (_24554_, _24553_, _24440_);
  nor (_24555_, _24417_, _24408_);
  and (_24556_, _24555_, _24554_);
  and (_24558_, _24556_, _24552_);
  and (_24559_, _24556_, _24536_);
  nor (_24560_, _24559_, _24558_);
  and (_24561_, _24560_, _24550_);
  nor (_24562_, _24561_, _24382_);
  not (_24563_, _24562_);
  not (_24564_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_24565_, \oc8051_top_1.oc8051_decoder1.state [1], _22766_);
  and (_24566_, _24565_, _24564_);
  and (_24567_, _24555_, _24446_);
  and (_24568_, _24567_, _24539_);
  and (_24569_, _24568_, _24566_);
  nor (_24570_, _24560_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_24572_, _24570_, _23837_);
  nor (_24573_, _24572_, _24569_);
  and (_24574_, _24573_, _24563_);
  nor (_24575_, _24574_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_24576_, _24575_, _24381_);
  not (_24577_, _24576_);
  and (_24578_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_24579_, _24578_);
  and (_24581_, _24554_, _24417_);
  and (_24582_, _24544_, _24490_);
  and (_24584_, _24582_, _24512_);
  and (_24585_, _24584_, _24581_);
  and (_24586_, _24581_, _24546_);
  or (_24587_, _24586_, _24585_);
  and (_24588_, _24539_, _24544_);
  and (_24589_, _24588_, _24538_);
  and (_24591_, _24581_, _24589_);
  nor (_24592_, _24512_, _24490_);
  and (_24593_, _24592_, _24534_);
  and (_24594_, _24593_, _24581_);
  or (_24595_, _24594_, _24591_);
  and (_24596_, _24581_, _24471_);
  and (_24597_, _24534_, _24490_);
  and (_24598_, _24597_, _24512_);
  or (_24599_, _24598_, _24588_);
  and (_24600_, _24599_, _24596_);
  or (_24601_, _24600_, _24595_);
  nor (_24602_, _24601_, _24587_);
  and (_24604_, _24540_, _24471_);
  and (_24605_, _24581_, _24604_);
  and (_24606_, _24535_, _24538_);
  and (_24607_, _24606_, _24581_);
  and (_24608_, _24581_, _24552_);
  or (_24610_, _24608_, _24607_);
  nor (_24611_, _24610_, _24605_);
  not (_24612_, _24408_);
  and (_24613_, _24447_, _24612_);
  and (_24614_, _24613_, _24593_);
  not (_24615_, _24614_);
  and (_24616_, _24592_, _24544_);
  and (_24617_, _24616_, _24581_);
  and (_24618_, _24584_, _24538_);
  and (_24619_, _24618_, _24567_);
  nor (_24620_, _24619_, _24617_);
  and (_24621_, _24620_, _24615_);
  and (_24622_, _24621_, _24611_);
  and (_24623_, _24622_, _24602_);
  and (_24624_, _24623_, _24550_);
  nor (_24625_, _24624_, _24382_);
  and (_24626_, \oc8051_top_1.oc8051_decoder1.state [0], _22766_);
  and (_24627_, _24626_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_24628_, _24614_, _24627_);
  and (_24629_, _24566_, _24540_);
  and (_24630_, _24629_, _24567_);
  or (_24631_, _24630_, _24628_);
  or (_24632_, _24631_, _24625_);
  nand (_24633_, _24632_, _22766_);
  and (_24634_, _24633_, _24579_);
  nor (_24635_, _24634_, _24577_);
  and (_26909_, _24635_, _22762_);
  and (_24636_, _24375_, _23747_);
  and (_24637_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_27175_, _24637_, _24636_);
  and (_24639_, _24356_, _24005_);
  and (_24640_, _24639_, _24050_);
  not (_24641_, _24639_);
  and (_24642_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_27170_, _24642_, _24640_);
  and (_24643_, _23053_, _23034_);
  nor (_24644_, _23002_, _22970_);
  and (_24645_, _24068_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_24646_, _24645_, _22943_);
  and (_24647_, _24646_, _24644_);
  and (_24648_, _24647_, _24643_);
  and (_24649_, _24648_, _24118_);
  nand (_24650_, _24649_, _23594_);
  or (_24651_, _24649_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_24652_, _24069_, _23002_);
  nor (_24653_, _23065_, _22983_);
  and (_24654_, _24653_, _24065_);
  and (_24655_, _24654_, _24652_);
  nor (_24656_, _23052_, _22970_);
  and (_24657_, _24656_, _23753_);
  and (_24658_, _24657_, _24655_);
  not (_24659_, _24658_);
  and (_24660_, _24659_, _24651_);
  and (_24661_, _24660_, _24650_);
  and (_24662_, _24658_, _23738_);
  or (_24663_, _24662_, _24661_);
  and (_06844_, _24663_, _22762_);
  and (_24664_, _24648_, _24291_);
  nand (_24665_, _24664_, _23594_);
  or (_24666_, _24664_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_24667_, _24666_, _24659_);
  and (_24668_, _24667_, _24665_);
  and (_24669_, _24658_, _23816_);
  or (_24670_, _24669_, _24668_);
  and (_06893_, _24670_, _22762_);
  and (_24671_, _24648_, _24067_);
  nand (_24672_, _24671_, _23594_);
  or (_24673_, _24671_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24674_, _24673_, _24659_);
  and (_24675_, _24674_, _24672_);
  and (_24676_, _24658_, _23892_);
  or (_24677_, _24676_, _24675_);
  and (_06909_, _24677_, _22762_);
  and (_24678_, _24066_, _23018_);
  and (_24679_, _24678_, _24648_);
  nand (_24680_, _24679_, _23594_);
  or (_24682_, _24679_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_24683_, _24682_, _24659_);
  and (_24684_, _24683_, _24680_);
  not (_24685_, _23772_);
  and (_24686_, _24658_, _24685_);
  or (_24687_, _24686_, _24684_);
  and (_06934_, _24687_, _22762_);
  and (_24688_, _24356_, _23903_);
  and (_24689_, _24688_, _23898_);
  not (_24690_, _24688_);
  and (_24691_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or (_06977_, _24691_, _24689_);
  and (_24692_, _24201_, _23656_);
  not (_24693_, _24692_);
  and (_24694_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and (_24695_, _24692_, _23898_);
  or (_07011_, _24695_, _24694_);
  and (_24696_, _24688_, _23747_);
  and (_24698_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  or (_07034_, _24698_, _24696_);
  and (_24699_, _24370_, _24329_);
  and (_24700_, _24699_, _23824_);
  not (_24701_, _24699_);
  and (_24702_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or (_07185_, _24702_, _24700_);
  and (_24703_, _24688_, _23946_);
  and (_24704_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or (_07208_, _24704_, _24703_);
  and (_24705_, _24653_, _23018_);
  and (_24706_, _24705_, _24648_);
  nand (_24707_, _24706_, _23594_);
  or (_24708_, _24706_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_24709_, _24708_, _24659_);
  and (_24710_, _24709_, _24707_);
  and (_24711_, _24658_, _24043_);
  or (_24712_, _24711_, _24710_);
  and (_07234_, _24712_, _22762_);
  and (_24713_, _24688_, _23707_);
  and (_24714_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or (_27171_, _24714_, _24713_);
  and (_24715_, _24648_, _24125_);
  nand (_24716_, _24715_, _23594_);
  or (_24717_, _24715_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_24718_, _24717_, _24659_);
  and (_24719_, _24718_, _24716_);
  and (_24720_, _24658_, _23939_);
  or (_24721_, _24720_, _24719_);
  and (_07281_, _24721_, _22762_);
  and (_24722_, _24356_, _23991_);
  and (_24723_, _24722_, _23778_);
  not (_24724_, _24722_);
  and (_24725_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or (_27173_, _24725_, _24723_);
  and (_24726_, _24722_, _23898_);
  and (_24727_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  or (_07490_, _24727_, _24726_);
  and (_24728_, _23003_, _22970_);
  and (_24729_, _24728_, _24646_);
  and (_24730_, _24729_, _24643_);
  and (_24731_, _24730_, _24067_);
  nand (_24732_, _24731_, _23594_);
  and (_24733_, _23053_, _22970_);
  and (_24734_, _24733_, _23753_);
  and (_24735_, _24678_, _24071_);
  and (_24736_, _24735_, _24734_);
  not (_24737_, _24736_);
  or (_24738_, _24731_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_24739_, _24738_, _24737_);
  and (_24740_, _24739_, _24732_);
  and (_24741_, _24736_, _23892_);
  or (_24742_, _24741_, _24740_);
  and (_07512_, _24742_, _22762_);
  and (_24743_, _24722_, _23649_);
  and (_24744_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  or (_07528_, _24744_, _24743_);
  and (_24745_, _24296_, _23711_);
  nor (_24746_, _24295_, _24123_);
  and (_24747_, _24746_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_24748_, _24747_, _24745_);
  and (_24749_, _24748_, _24730_);
  not (_24750_, _24730_);
  nor (_24751_, _24295_, _23065_);
  or (_24752_, _24751_, _24678_);
  or (_24753_, _24752_, _24750_);
  and (_24754_, _24753_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_24755_, _24754_, _24736_);
  or (_24756_, _24755_, _24749_);
  or (_24757_, _24737_, _23642_);
  and (_24758_, _24757_, _22762_);
  and (_07548_, _24758_, _24756_);
  and (_24759_, _24730_, _24118_);
  nand (_24760_, _24759_, _23594_);
  or (_24761_, _24759_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_24762_, _24761_, _24737_);
  and (_24763_, _24762_, _24760_);
  and (_24764_, _24736_, _23738_);
  or (_24765_, _24764_, _24763_);
  and (_07595_, _24765_, _22762_);
  and (_24766_, _23905_, _23753_);
  and (_24767_, _24766_, _24275_);
  not (_24768_, _24767_);
  and (_24769_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_24770_, _24767_, _23747_);
  or (_07629_, _24770_, _24769_);
  and (_24771_, _24730_, _24291_);
  nand (_24772_, _24771_, _23594_);
  or (_24773_, _24771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_24774_, _24773_, _24737_);
  and (_24775_, _24774_, _24772_);
  and (_24776_, _24736_, _23816_);
  or (_24777_, _24776_, _24775_);
  and (_07661_, _24777_, _22762_);
  and (_24778_, _24730_, _24678_);
  nand (_24779_, _24778_, _23594_);
  or (_24780_, _24778_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_24781_, _24780_, _24737_);
  and (_24782_, _24781_, _24779_);
  and (_24783_, _24736_, _24685_);
  or (_24784_, _24783_, _24782_);
  and (_07683_, _24784_, _22762_);
  and (_24785_, _24722_, _23946_);
  and (_24786_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  or (_07737_, _24786_, _24785_);
  and (_24787_, _24722_, _23707_);
  and (_24788_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or (_07894_, _24788_, _24787_);
  and (_24789_, _24356_, _24275_);
  and (_24790_, _24789_, _23778_);
  not (_24791_, _24789_);
  and (_24792_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_07925_, _24792_, _24790_);
  and (_24793_, _24789_, _23747_);
  and (_24794_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_07944_, _24794_, _24793_);
  and (_24795_, _24730_, _24705_);
  nand (_24796_, _24795_, _23594_);
  or (_24797_, _24795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_24798_, _24797_, _24737_);
  and (_24799_, _24798_, _24796_);
  and (_24800_, _24736_, _24043_);
  or (_24801_, _24800_, _24799_);
  and (_07995_, _24801_, _22762_);
  and (_24802_, _24789_, _23649_);
  and (_24803_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_08032_, _24803_, _24802_);
  and (_24804_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_24805_, _24767_, _23824_);
  or (_08049_, _24805_, _24804_);
  and (_24806_, _24789_, _24050_);
  and (_24807_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_08086_, _24807_, _24806_);
  and (_24808_, _24789_, _23707_);
  and (_24809_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_08131_, _24809_, _24808_);
  and (_24810_, _24375_, _24050_);
  and (_24811_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_08161_, _24811_, _24810_);
  and (_24812_, _23052_, _23034_);
  and (_24813_, _24812_, _24729_);
  and (_24814_, _24813_, _24296_);
  or (_24815_, _24814_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_24816_, _24735_, _24064_);
  not (_24817_, _24816_);
  and (_24818_, _24817_, _24815_);
  nand (_24819_, _24814_, _23594_);
  and (_24820_, _24819_, _24818_);
  and (_24821_, _24816_, _23642_);
  or (_24822_, _24821_, _24820_);
  and (_08221_, _24822_, _22762_);
  and (_24823_, _24813_, _24291_);
  nand (_24824_, _24823_, _23594_);
  or (_24825_, _24823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_24826_, _24825_, _24817_);
  and (_24827_, _24826_, _24824_);
  and (_24828_, _24816_, _23816_);
  or (_24829_, _24828_, _24827_);
  and (_08240_, _24829_, _22762_);
  and (_24830_, _24813_, _24678_);
  or (_24831_, _24830_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_24832_, _24831_, _24817_);
  nand (_24833_, _24830_, _23594_);
  and (_24834_, _24833_, _24832_);
  and (_24835_, _24816_, _24685_);
  or (_24836_, _24835_, _24834_);
  and (_08258_, _24836_, _22762_);
  and (_24837_, _24375_, _23707_);
  and (_24838_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_27176_, _24838_, _24837_);
  and (_24839_, _24370_, _24085_);
  and (_24840_, _24839_, _23898_);
  not (_24841_, _24839_);
  and (_24842_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or (_08365_, _24842_, _24840_);
  and (_24843_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_24844_, _24767_, _23898_);
  or (_08380_, _24844_, _24843_);
  or (_24845_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_24846_, _24845_, _22762_);
  or (_24847_, _24079_, _23642_);
  and (_08395_, _24847_, _24846_);
  and (_24848_, _24839_, _23824_);
  and (_24849_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  or (_08416_, _24849_, _24848_);
  and (_24850_, _24839_, _23946_);
  and (_24851_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  or (_08466_, _24851_, _24850_);
  and (_24852_, _23911_, _23076_);
  and (_24853_, _24852_, _23649_);
  not (_24854_, _24852_);
  and (_24855_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  or (_08496_, _24855_, _24853_);
  and (_24856_, _24839_, _24050_);
  and (_24857_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or (_08544_, _24857_, _24856_);
  and (_24858_, _24370_, _24010_);
  and (_24859_, _24858_, _23778_);
  not (_24860_, _24858_);
  and (_24861_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or (_08572_, _24861_, _24859_);
  and (_24862_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_24863_, _24862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_24864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_24865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_24866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _24865_);
  and (_24867_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_24868_, _24867_, _24866_);
  and (_24869_, _24868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_24870_, _24869_, _24864_);
  not (_24871_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_24872_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_24873_, _24872_, _24871_);
  nand (_24874_, _24873_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_24875_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_24876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_24877_, _24876_, _24875_);
  and (_24878_, _24877_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_24879_, _24878_);
  and (_24880_, _24879_, _24874_);
  and (_24881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_24882_, _24881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_24883_, _24882_);
  and (_24884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_24885_, _24884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_24887_, _24886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_24888_, _24887_, _24885_);
  and (_24889_, _24888_, _24883_);
  and (_24890_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_24891_, _24890_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_24892_, _24891_);
  and (_24893_, _24892_, _24889_);
  and (_24894_, _24893_, _24880_);
  nor (_24895_, _24894_, _24870_);
  and (_24896_, _24864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not (_24897_, _24896_);
  not (_24898_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_24899_, _24873_, _24898_);
  not (_24900_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_24901_, _24877_, _24900_);
  nor (_24902_, _24901_, _24899_);
  not (_24903_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_24904_, _24890_, _24903_);
  not (_24905_, _24904_);
  not (_24906_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_24907_, _24881_, _24906_);
  not (_24908_, _24907_);
  not (_24909_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24910_, _24884_, _24909_);
  not (_24911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_24912_, _24886_, _24911_);
  nor (_24913_, _24912_, _24910_);
  and (_24914_, _24913_, _24908_);
  and (_24915_, _24914_, _24905_);
  and (_24916_, _24915_, _24902_);
  or (_24917_, _24916_, _24897_);
  nor (_24918_, _24917_, _24895_);
  nand (_24919_, _24918_, _24863_);
  and (_24920_, _24895_, _24863_);
  or (_24921_, _24920_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and (_24922_, _24921_, _22762_);
  and (_08672_, _24922_, _24919_);
  and (_24923_, _24858_, _23898_);
  and (_24924_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  or (_27177_, _24924_, _24923_);
  and (_24925_, _24858_, _23649_);
  and (_24926_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or (_27178_, _24926_, _24925_);
  and (_24927_, _24858_, _24050_);
  and (_24928_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  or (_08777_, _24928_, _24927_);
  nand (_24929_, _24530_, _22767_);
  or (_24930_, _22767_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_24931_, _24930_, _22762_);
  and (_26864_[5], _24931_, _24929_);
  and (_24932_, _24370_, _23911_);
  and (_24933_, _24932_, _23898_);
  not (_24934_, _24932_);
  and (_24935_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_08852_, _24935_, _24933_);
  and (_24936_, _24932_, _23747_);
  and (_24937_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_08908_, _24937_, _24936_);
  nor (_24938_, _24862_, _24865_);
  nand (_24939_, _24938_, _24918_);
  and (_24940_, _24938_, _24895_);
  or (_24941_, _24940_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and (_24942_, _24941_, _22762_);
  and (_08926_, _24942_, _24939_);
  and (_24943_, _24932_, _23946_);
  and (_24944_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_09009_, _24944_, _24943_);
  and (_24945_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_24946_, _24767_, _23946_);
  or (_09056_, _24946_, _24945_);
  and (_24947_, _24932_, _23707_);
  and (_24948_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_09081_, _24948_, _24947_);
  not (_24949_, _24917_);
  nor (_24950_, _24949_, _24895_);
  nor (_24951_, _24950_, _24862_);
  not (_24952_, _24951_);
  and (_24953_, _24952_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_24954_, _24862_);
  nor (_24955_, _24874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_24956_, _24955_, _24891_);
  not (_24957_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_24958_, _24878_, _24865_);
  or (_24959_, _24958_, _24957_);
  nand (_24960_, _24959_, _24956_);
  and (_24961_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_24962_, _24961_, _24892_);
  and (_24963_, _24962_, _24960_);
  or (_24964_, _24963_, _24887_);
  not (_24965_, _24885_);
  not (_24966_, _24887_);
  or (_24967_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _24865_);
  or (_24968_, _24967_, _24966_);
  and (_24969_, _24968_, _24965_);
  and (_24970_, _24969_, _24964_);
  and (_24971_, _24961_, _24885_);
  or (_24972_, _24971_, _24882_);
  or (_24973_, _24972_, _24970_);
  or (_24974_, _24967_, _24883_);
  and (_24975_, _24974_, _24895_);
  and (_24976_, _24975_, _24973_);
  or (_24977_, _24967_, _24908_);
  and (_24978_, _24899_, _24865_);
  nor (_24979_, _24978_, _24904_);
  and (_24980_, _24901_, _24865_);
  or (_24981_, _24980_, _24957_);
  nand (_24982_, _24981_, _24979_);
  or (_24983_, _24961_, _24905_);
  and (_24984_, _24983_, _24982_);
  or (_24985_, _24984_, _24912_);
  not (_24986_, _24910_);
  not (_24987_, _24912_);
  or (_24988_, _24967_, _24987_);
  and (_24989_, _24988_, _24986_);
  and (_24990_, _24989_, _24985_);
  and (_24991_, _24961_, _24910_);
  or (_24992_, _24991_, _24907_);
  or (_24993_, _24992_, _24990_);
  and (_24994_, _24993_, _24918_);
  and (_24995_, _24994_, _24977_);
  or (_24996_, _24995_, _24976_);
  and (_24997_, _24996_, _24954_);
  or (_24998_, _24997_, _24953_);
  and (_09127_, _24998_, _22762_);
  and (_24999_, _24370_, _24282_);
  and (_25000_, _24999_, _23778_);
  not (_25001_, _24999_);
  and (_25002_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_09156_, _25002_, _25000_);
  nand (_25003_, _24950_, _24863_);
  nor (_25004_, _24895_, _24862_);
  or (_25005_, _25004_, _24865_);
  and (_25006_, _25005_, _22762_);
  and (_09190_, _25006_, _25003_);
  and (_25007_, _24999_, _23747_);
  and (_25008_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_27183_, _25008_, _25007_);
  and (_25009_, _24999_, _23946_);
  and (_25010_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_09277_, _25010_, _25009_);
  and (_25011_, _24999_, _23707_);
  and (_25012_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_09338_, _25012_, _25011_);
  and (_25013_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_25014_, _24236_, _24145_);
  nand (_25015_, _25014_, _24153_);
  and (_25016_, _25015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  not (_25017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_25018_, _25014_, _24256_);
  or (_25019_, _25018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_25020_, _25019_, _25017_);
  or (_25021_, _25020_, _25016_);
  nor (_25022_, _24153_, _24182_);
  or (_25023_, _25022_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_25024_, _25023_);
  and (_25025_, _24235_, _24145_);
  and (_25026_, _25025_, _25024_);
  or (_25027_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand (_25028_, _25027_, _25021_);
  nor (_25029_, _25028_, _24127_);
  and (_25030_, _24127_, _23816_);
  or (_25031_, _25030_, _25029_);
  and (_25032_, _25031_, _24166_);
  or (_09365_, _25032_, _25013_);
  and (_25033_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_25034_, _24767_, _24050_);
  or (_09393_, _25034_, _25033_);
  not (_25035_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor (_25036_, _24951_, _25035_);
  or (_25037_, _24892_, _24887_);
  and (_25038_, _25037_, _24965_);
  and (_25039_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _24865_);
  or (_25040_, _25039_, _25038_);
  and (_25041_, _24878_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_25042_, _25041_, _25035_);
  nor (_25043_, _24874_, _24865_);
  nor (_25044_, _25043_, _24891_);
  nand (_25045_, _25044_, _24888_);
  or (_25046_, _25045_, _25042_);
  and (_25047_, _25046_, _25040_);
  or (_25048_, _25047_, _24882_);
  or (_25049_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25050_, _24966_, _24885_);
  and (_25051_, _25050_, _24883_);
  or (_25052_, _25051_, _25049_);
  and (_25053_, _25052_, _24895_);
  and (_25054_, _25053_, _25048_);
  and (_25055_, _24899_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_25056_, _25055_, _24904_);
  and (_25057_, _24901_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25058_, _25057_, _25035_);
  nand (_25059_, _25058_, _25056_);
  or (_25060_, _25039_, _24905_);
  and (_25061_, _25060_, _25059_);
  or (_25062_, _25061_, _24912_);
  or (_25063_, _25049_, _24987_);
  and (_25064_, _25063_, _24986_);
  and (_25065_, _25064_, _25062_);
  and (_25066_, _25039_, _24910_);
  or (_25067_, _25066_, _24907_);
  or (_25068_, _25067_, _25065_);
  and (_25069_, _24918_, _24908_);
  and (_25070_, _25049_, _24918_);
  or (_25071_, _25070_, _25069_);
  and (_25072_, _25071_, _25068_);
  or (_25073_, _25072_, _25054_);
  and (_25074_, _25073_, _24954_);
  or (_25075_, _25074_, _25036_);
  and (_09413_, _25075_, _22762_);
  and (_25076_, _24852_, _23824_);
  and (_25077_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or (_09433_, _25077_, _25076_);
  and (_25078_, _23901_, _23655_);
  and (_25079_, _25078_, _24370_);
  and (_25080_, _25079_, _23778_);
  not (_25081_, _25079_);
  and (_25082_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  or (_09490_, _25082_, _25080_);
  and (_25083_, _25079_, _23824_);
  and (_25084_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or (_09519_, _25084_, _25083_);
  and (_25085_, _25079_, _23649_);
  and (_25086_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or (_27185_, _25086_, _25085_);
  and (_25087_, _25079_, _24050_);
  and (_25088_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or (_09609_, _25088_, _25087_);
  and (_25089_, _25079_, _23707_);
  and (_25090_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or (_09650_, _25090_, _25089_);
  and (_25091_, _24370_, _23656_);
  and (_25092_, _25091_, _23824_);
  not (_25093_, _25091_);
  and (_25094_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  or (_09680_, _25094_, _25092_);
  and (_25095_, _24862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_25096_, _25095_, _24951_);
  and (_09728_, _25096_, _22762_);
  nand (_25097_, _24915_, _24896_);
  or (_25098_, _25097_, _24902_);
  nor (_25099_, _25098_, _24895_);
  and (_25100_, _24862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  not (_25101_, _24870_);
  nand (_25102_, _24893_, _25101_);
  nor (_25103_, _25102_, _24880_);
  and (_25104_, _25103_, _24954_);
  or (_25105_, _25104_, _25100_);
  or (_25106_, _25105_, _25099_);
  and (_09750_, _25106_, _22762_);
  nor (_25108_, _24910_, _24907_);
  or (_25109_, _24912_, _24904_);
  and (_25110_, _24902_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_25111_, _25110_, _25109_);
  and (_25112_, _25111_, _25108_);
  and (_25113_, _25112_, _24918_);
  nor (_25114_, _24885_, _24882_);
  or (_25115_, _24891_, _24887_);
  and (_25116_, _24880_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_25117_, _25116_, _25115_);
  and (_25118_, _25117_, _25114_);
  and (_25119_, _25118_, _24895_);
  or (_25120_, _25119_, _25113_);
  or (_25121_, _25120_, _24862_);
  or (_25122_, _24954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_25123_, _25122_, _22762_);
  and (_09772_, _25123_, _25121_);
  nor (_25125_, _24901_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_25126_, _25125_, _24899_);
  or (_25127_, _25126_, _24904_);
  and (_25128_, _25127_, _24987_);
  or (_25129_, _25128_, _24910_);
  and (_25130_, _25129_, _25069_);
  or (_25131_, _24878_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_25132_, _25131_, _24874_);
  or (_25133_, _25132_, _24891_);
  and (_25134_, _25133_, _24966_);
  or (_25135_, _25134_, _24885_);
  and (_25136_, _24895_, _24883_);
  and (_25137_, _25136_, _25135_);
  or (_25138_, _25137_, _24862_);
  or (_25139_, _25138_, _25130_);
  or (_25140_, _24954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_25141_, _25140_, _22762_);
  and (_09791_, _25141_, _25139_);
  and (_25142_, _24370_, _24275_);
  and (_25143_, _25142_, _23778_);
  not (_25144_, _25142_);
  and (_25145_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  or (_27199_, _25145_, _25143_);
  and (_25146_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _22762_);
  and (_09843_, _25146_, _24862_);
  and (_25148_, _25091_, _23747_);
  and (_25150_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  or (_27187_, _25150_, _25148_);
  and (_25151_, _25091_, _23946_);
  and (_25153_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or (_09958_, _25153_, _25151_);
  and (_25154_, _25091_, _23707_);
  and (_25155_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or (_09981_, _25155_, _25154_);
  and (_25156_, _24370_, _23752_);
  and (_25157_, _25156_, _23898_);
  not (_25158_, _25156_);
  and (_25159_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_10015_, _25159_, _25157_);
  and (_25160_, _25156_, _23824_);
  and (_25161_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_10138_, _25161_, _25160_);
  nor (_25162_, _23003_, _22970_);
  and (_25163_, _25162_, _22943_);
  and (_25164_, _25163_, _24643_);
  and (_25165_, _25164_, _24118_);
  nand (_25166_, _25165_, _23594_);
  or (_25167_, _25165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_25168_, _25167_, _24645_);
  and (_25169_, _25168_, _25166_);
  and (_25170_, _23065_, _23002_);
  and (_25171_, _25170_, _24295_);
  and (_25172_, _25171_, _24656_);
  and (_25173_, _25172_, _23753_);
  not (_25174_, _25173_);
  or (_25175_, _25174_, _23738_);
  or (_25176_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_25178_, _25176_, _24069_);
  and (_25179_, _25178_, _25175_);
  not (_25181_, _24068_);
  and (_25182_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_25183_, _25182_, rst);
  or (_25184_, _25183_, _25179_);
  or (_10161_, _25184_, _25169_);
  and (_25185_, _25164_, _24291_);
  nand (_25186_, _25185_, _23594_);
  or (_25187_, _25185_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_25188_, _25187_, _24645_);
  and (_25189_, _25188_, _25186_);
  or (_25190_, _25174_, _23816_);
  or (_25191_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_25192_, _25191_, _24069_);
  and (_25193_, _25192_, _25190_);
  and (_25194_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_25195_, _25194_, rst);
  or (_25196_, _25195_, _25193_);
  or (_10186_, _25196_, _25189_);
  and (_25197_, _25164_, _24067_);
  nand (_25198_, _25197_, _23594_);
  or (_25199_, _25197_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_25200_, _25199_, _24645_);
  and (_25201_, _25200_, _25198_);
  or (_25202_, _25174_, _23892_);
  or (_25203_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_25204_, _25203_, _24069_);
  and (_25205_, _25204_, _25202_);
  and (_25206_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_25207_, _25206_, rst);
  or (_25208_, _25207_, _25205_);
  or (_10212_, _25208_, _25201_);
  and (_25209_, _25164_, _24678_);
  nand (_25210_, _25209_, _23594_);
  or (_25211_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_25212_, _25211_, _24645_);
  and (_25213_, _25212_, _25210_);
  nand (_25214_, _25173_, _23772_);
  and (_25215_, _25214_, _24069_);
  and (_25216_, _25215_, _25211_);
  not (_25217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_25218_, _24068_, _25217_);
  or (_25219_, _25218_, rst);
  or (_25220_, _25219_, _25216_);
  or (_10236_, _25220_, _25213_);
  and (_25221_, _25156_, _23649_);
  and (_25222_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_10291_, _25222_, _25221_);
  and (_25223_, _25156_, _24050_);
  and (_25224_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_27188_, _25224_, _25223_);
  and (_25225_, _25164_, _24705_);
  nand (_25226_, _25225_, _23594_);
  or (_25227_, _25225_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_25228_, _25227_, _24645_);
  and (_25229_, _25228_, _25226_);
  or (_25230_, _25174_, _24043_);
  or (_25231_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_25232_, _25231_, _24069_);
  and (_25233_, _25232_, _25230_);
  not (_25234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_25235_, _24068_, _25234_);
  or (_25236_, _25235_, rst);
  or (_25237_, _25236_, _25233_);
  or (_10409_, _25237_, _25229_);
  and (_25238_, _25164_, _24125_);
  nand (_25239_, _25238_, _23594_);
  or (_25240_, _25238_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_25241_, _25240_, _24645_);
  and (_25242_, _25241_, _25239_);
  or (_25243_, _25174_, _23939_);
  or (_25244_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_25245_, _25244_, _24069_);
  and (_25246_, _25245_, _25243_);
  and (_25247_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_25248_, _25247_, rst);
  or (_25249_, _25248_, _25246_);
  or (_10540_, _25249_, _25242_);
  and (_25250_, _24358_, _23649_);
  and (_25251_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or (_10604_, _25251_, _25250_);
  and (_25252_, _24766_, _23991_);
  not (_25253_, _25252_);
  and (_25254_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  and (_25255_, _25252_, _24050_);
  or (_10628_, _25255_, _25254_);
  and (_25256_, _24358_, _23747_);
  and (_25257_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or (_10652_, _25257_, _25256_);
  and (_25258_, _23002_, _22970_);
  and (_25259_, _25258_, _22943_);
  and (_25260_, _25259_, _24643_);
  and (_25261_, _25260_, _24067_);
  nand (_25262_, _25261_, _23594_);
  or (_25263_, _25261_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_25264_, _25263_, _24645_);
  and (_25265_, _25264_, _25262_);
  and (_25266_, _25171_, _24734_);
  not (_25267_, _25266_);
  or (_25268_, _25267_, _23892_);
  or (_25269_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_25270_, _25269_, _24069_);
  and (_25271_, _25270_, _25268_);
  and (_25272_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_25273_, _25272_, rst);
  or (_25274_, _25273_, _25271_);
  or (_10718_, _25274_, _25265_);
  and (_25275_, _25260_, _24125_);
  nand (_25276_, _25275_, _23594_);
  or (_25277_, _25275_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_25278_, _25277_, _24645_);
  and (_25279_, _25278_, _25276_);
  or (_25280_, _25267_, _23939_);
  or (_25281_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_25282_, _25281_, _24069_);
  and (_25283_, _25282_, _25280_);
  and (_25284_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_25286_, _25284_, rst);
  or (_25287_, _25286_, _25283_);
  or (_10757_, _25287_, _25279_);
  and (_25289_, _25260_, _24296_);
  nand (_25290_, _25289_, _23594_);
  or (_25291_, _25289_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_25292_, _25291_, _24645_);
  and (_25293_, _25292_, _25290_);
  or (_25294_, _25267_, _23642_);
  or (_25296_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_25297_, _25296_, _24069_);
  and (_25299_, _25297_, _25294_);
  not (_25300_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_25301_, _24068_, _25300_);
  or (_25302_, _25301_, rst);
  or (_25303_, _25302_, _25299_);
  or (_10779_, _25303_, _25293_);
  and (_25304_, _25260_, _24118_);
  nand (_25305_, _25304_, _23594_);
  or (_25306_, _25304_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_25307_, _25306_, _24645_);
  and (_25308_, _25307_, _25305_);
  or (_25309_, _25267_, _23738_);
  or (_25310_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_25311_, _25310_, _24069_);
  and (_25312_, _25311_, _25309_);
  and (_25313_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_25314_, _25313_, rst);
  or (_25315_, _25314_, _25312_);
  or (_10829_, _25315_, _25308_);
  and (_25316_, _25260_, _24291_);
  nand (_25317_, _25316_, _23594_);
  or (_25318_, _25316_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_25319_, _25318_, _24645_);
  and (_25320_, _25319_, _25317_);
  or (_25321_, _25267_, _23816_);
  or (_25322_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_25323_, _25322_, _24069_);
  and (_25324_, _25323_, _25321_);
  and (_25325_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_25326_, _25325_, rst);
  or (_25327_, _25326_, _25324_);
  or (_10855_, _25327_, _25320_);
  and (_25328_, _25260_, _24678_);
  nand (_25329_, _25328_, _23594_);
  or (_25330_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_25331_, _25330_, _24645_);
  and (_25332_, _25331_, _25329_);
  nand (_25333_, _25266_, _23772_);
  and (_25334_, _25333_, _24069_);
  and (_25335_, _25334_, _25330_);
  not (_25336_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_25337_, _24068_, _25336_);
  or (_25338_, _25337_, rst);
  or (_25339_, _25338_, _25335_);
  or (_10891_, _25339_, _25332_);
  and (_25340_, _24356_, _23911_);
  and (_25341_, _25340_, _23649_);
  not (_25342_, _25340_);
  and (_25343_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  or (_27081_, _25343_, _25341_);
  and (_25345_, _25340_, _23747_);
  and (_25346_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  or (_11051_, _25346_, _25345_);
  and (_25348_, _25340_, _23824_);
  and (_25349_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or (_11091_, _25349_, _25348_);
  and (_25350_, _25163_, _24812_);
  and (_25352_, _25350_, _24118_);
  nand (_25353_, _25352_, _23594_);
  or (_25354_, _25352_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_25355_, _25354_, _24645_);
  and (_25356_, _25355_, _25353_);
  and (_25358_, _25350_, _24678_);
  not (_25359_, _25358_);
  or (_25360_, _25359_, _23738_);
  or (_25361_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_25362_, _25361_, _24069_);
  and (_25363_, _25362_, _25360_);
  and (_25364_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_25365_, _25364_, rst);
  or (_25367_, _25365_, _25363_);
  or (_11413_, _25367_, _25356_);
  and (_25368_, _25350_, _24291_);
  nand (_25369_, _25368_, _23594_);
  or (_25370_, _25368_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_25371_, _25370_, _24645_);
  and (_25372_, _25371_, _25369_);
  or (_25373_, _25359_, _23816_);
  or (_25374_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_25375_, _25374_, _24069_);
  and (_25376_, _25375_, _25373_);
  and (_25377_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_25378_, _25377_, rst);
  or (_25379_, _25378_, _25376_);
  or (_11482_, _25379_, _25372_);
  and (_25380_, _25350_, _24067_);
  nand (_25381_, _25380_, _23594_);
  or (_25382_, _25380_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_25383_, _25382_, _24645_);
  and (_25384_, _25383_, _25381_);
  or (_25385_, _25359_, _23892_);
  or (_25386_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_25387_, _25386_, _24069_);
  and (_25388_, _25387_, _25385_);
  and (_25389_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_25390_, _25389_, rst);
  or (_25391_, _25390_, _25388_);
  or (_11558_, _25391_, _25384_);
  nand (_25393_, _25358_, _23594_);
  or (_25394_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_25395_, _25394_, _24645_);
  and (_25396_, _25395_, _25393_);
  nand (_25397_, _25358_, _23772_);
  and (_25398_, _25397_, _24069_);
  and (_25399_, _25398_, _25394_);
  not (_25400_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_25401_, _24068_, _25400_);
  or (_25402_, _25401_, rst);
  or (_25403_, _25402_, _25399_);
  or (_11583_, _25403_, _25396_);
  and (_25404_, _25340_, _23707_);
  and (_25405_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or (_11681_, _25405_, _25404_);
  and (_25406_, _25340_, _24050_);
  and (_25407_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  or (_11792_, _25407_, _25406_);
  and (_25408_, _25350_, _24705_);
  nand (_25409_, _25408_, _23594_);
  or (_25410_, _25408_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_25411_, _25410_, _24645_);
  and (_25412_, _25411_, _25409_);
  or (_25414_, _25359_, _24043_);
  or (_25415_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_25416_, _25415_, _24069_);
  and (_25417_, _25416_, _25414_);
  not (_25418_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_25419_, _24068_, _25418_);
  or (_25420_, _25419_, rst);
  or (_25421_, _25420_, _25417_);
  or (_11878_, _25421_, _25412_);
  and (_25422_, _25350_, _24125_);
  nand (_25423_, _25422_, _23594_);
  or (_25425_, _25422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_25426_, _25425_, _24645_);
  and (_25427_, _25426_, _25423_);
  or (_25429_, _25359_, _23939_);
  or (_25430_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_25431_, _25430_, _24069_);
  and (_25432_, _25431_, _25429_);
  and (_25433_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_25434_, _25433_, rst);
  or (_25435_, _25434_, _25432_);
  or (_11954_, _25435_, _25427_);
  and (_25437_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  and (_25438_, _25252_, _23898_);
  or (_11987_, _25438_, _25437_);
  and (_25439_, _25259_, _24812_);
  and (_25441_, _25439_, _24291_);
  nand (_25442_, _25441_, _23594_);
  or (_25443_, _25441_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_25444_, _25443_, _24645_);
  and (_25445_, _25444_, _25442_);
  and (_25446_, _25171_, _24064_);
  not (_25447_, _25446_);
  or (_25448_, _25447_, _23816_);
  or (_25449_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_25450_, _25449_, _24069_);
  and (_25451_, _25450_, _25448_);
  and (_25453_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_25455_, _25453_, rst);
  or (_25456_, _25455_, _25451_);
  or (_12139_, _25456_, _25445_);
  and (_25459_, _25439_, _24067_);
  nand (_25460_, _25459_, _23594_);
  or (_25461_, _25459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_25462_, _25461_, _24645_);
  and (_25464_, _25462_, _25460_);
  or (_25466_, _25447_, _23892_);
  or (_25467_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_25468_, _25467_, _24069_);
  and (_25469_, _25468_, _25466_);
  and (_25470_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_25472_, _25470_, rst);
  or (_25473_, _25472_, _25469_);
  or (_12170_, _25473_, _25464_);
  and (_25474_, _25439_, _24678_);
  nand (_25475_, _25474_, _23594_);
  or (_25476_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_25477_, _25476_, _24645_);
  and (_25479_, _25477_, _25475_);
  nand (_25480_, _25446_, _23772_);
  and (_25481_, _25476_, _24069_);
  and (_25482_, _25481_, _25480_);
  not (_25483_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_25484_, _24068_, _25483_);
  or (_25485_, _25484_, rst);
  or (_25486_, _25485_, _25482_);
  or (_12192_, _25486_, _25479_);
  and (_25488_, _24356_, _24010_);
  and (_25489_, _25488_, _24050_);
  not (_25490_, _25488_);
  and (_25491_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_12223_, _25491_, _25489_);
  and (_25493_, _25488_, _23946_);
  and (_25494_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_12344_, _25494_, _25493_);
  and (_25495_, _25439_, _24125_);
  nand (_25496_, _25495_, _23594_);
  or (_25497_, _25495_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_25498_, _25497_, _24645_);
  and (_25499_, _25498_, _25496_);
  or (_25500_, _25447_, _23939_);
  or (_25501_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_25502_, _25501_, _24069_);
  and (_25503_, _25502_, _25500_);
  and (_25504_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_25505_, _25504_, rst);
  or (_25506_, _25505_, _25503_);
  or (_12395_, _25506_, _25499_);
  and (_25507_, _25439_, _24705_);
  nand (_25508_, _25507_, _23594_);
  or (_25509_, _25507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_25510_, _25509_, _24645_);
  and (_25511_, _25510_, _25508_);
  or (_25512_, _25447_, _24043_);
  or (_25514_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_25515_, _25514_, _24069_);
  and (_25516_, _25515_, _25512_);
  not (_25517_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_25518_, _24068_, _25517_);
  or (_25519_, _25518_, rst);
  or (_25520_, _25519_, _25516_);
  or (_12507_, _25520_, _25511_);
  and (_25521_, _25439_, _24296_);
  nand (_25523_, _25521_, _23594_);
  or (_25524_, _25521_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_25525_, _25524_, _24645_);
  and (_25526_, _25525_, _25523_);
  or (_25527_, _25447_, _23642_);
  or (_25528_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_25529_, _25528_, _24069_);
  and (_25530_, _25529_, _25527_);
  not (_25531_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_25532_, _24068_, _25531_);
  or (_25533_, _25532_, rst);
  or (_25534_, _25533_, _25530_);
  or (_12529_, _25534_, _25526_);
  and (_25536_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  and (_25537_, _25252_, _23747_);
  or (_27043_, _25537_, _25536_);
  and (_25538_, _25340_, _23778_);
  and (_25539_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or (_27080_, _25539_, _25538_);
  and (_25540_, _25488_, _23707_);
  and (_25541_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_12805_, _25541_, _25540_);
  and (_25542_, _24766_, _23903_);
  not (_25543_, _25542_);
  and (_25544_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and (_25545_, _25542_, _23946_);
  or (_12920_, _25545_, _25544_);
  and (_25546_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  and (_25547_, _25542_, _24050_);
  or (_12950_, _25547_, _25546_);
  and (_25548_, _25488_, _23898_);
  and (_25549_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_14450_, _25549_, _25548_);
  nor (_25550_, _22768_, _23373_);
  and (_25551_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_25552_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_25553_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_25554_, _25553_, _25552_);
  and (_25555_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_25556_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_25557_, _25556_, _25555_);
  or (_25558_, _25557_, _25554_);
  and (_25559_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_25560_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_25561_, _25560_, _25559_);
  or (_25562_, _25561_, _25558_);
  and (_25563_, _25562_, _23839_);
  or (_25564_, _25563_, _25551_);
  and (_25565_, _25564_, _22768_);
  nor (_25566_, _25565_, _25550_);
  nor (_26897_[0], _25566_, rst);
  and (_25568_, _25488_, _23778_);
  and (_25570_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_14601_, _25570_, _25568_);
  and (_25571_, _24356_, _24085_);
  and (_25572_, _25571_, _23707_);
  not (_25573_, _25571_);
  and (_25574_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_14938_, _25574_, _25572_);
  or (_25576_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_25577_, _25576_, _22762_);
  or (_25579_, _24079_, _23939_);
  and (_15132_, _25579_, _25577_);
  and (_25581_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_25582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand (_25583_, _25582_, _24152_);
  nor (_25584_, _25583_, _24149_);
  and (_25586_, _24234_, _25584_);
  and (_25587_, _25586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_25588_, _25587_, _24145_);
  nand (_25590_, _25588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_25591_, _25588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_25592_, _25591_, _24132_);
  and (_25593_, _25592_, _25590_);
  and (_25594_, _25019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_25595_, _24256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_25596_, _25595_, _25014_);
  or (_25597_, _25596_, _25594_);
  nor (_25598_, _25597_, _25593_);
  nor (_25599_, _25598_, _24127_);
  and (_25601_, _24127_, _23738_);
  or (_25602_, _25601_, _25599_);
  and (_25603_, _25602_, _24166_);
  or (_15153_, _25603_, _25581_);
  and (_25604_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  and (_25605_, _25542_, _23707_);
  or (_15784_, _25605_, _25604_);
  and (_25607_, _25488_, _23747_);
  and (_25608_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_17267_, _25608_, _25607_);
  or (_25609_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_25610_, _25609_, _22762_);
  or (_25611_, _24079_, _24043_);
  and (_17294_, _25611_, _25610_);
  and (_25612_, _25488_, _23824_);
  and (_25613_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_17417_, _25613_, _25612_);
  and (_25615_, _23755_, _23747_);
  and (_25616_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  or (_17600_, _25616_, _25615_);
  and (_25618_, \oc8051_top_1.oc8051_sfr1.wait_data , _22762_);
  and (_25619_, _25618_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_25620_, _24567_, _24552_);
  and (_25621_, _24584_, _24471_);
  and (_25622_, _25621_, _24448_);
  or (_25623_, _25622_, _25620_);
  or (_25624_, _25623_, _24568_);
  and (_25625_, _24593_, _24471_);
  and (_25626_, _25625_, _24567_);
  and (_25627_, _24592_, _24538_);
  and (_25629_, _25627_, _24567_);
  nor (_25630_, _25629_, _25626_);
  and (_25631_, _25621_, _24613_);
  and (_25633_, _24618_, _24447_);
  nor (_25634_, _25633_, _25631_);
  nand (_25635_, _25634_, _25630_);
  and (_25636_, _24552_, _24448_);
  and (_25638_, _24598_, _24471_);
  and (_25639_, _25638_, _24556_);
  or (_25640_, _25639_, _25636_);
  or (_25641_, _25640_, _25635_);
  or (_25642_, _25641_, _25624_);
  and (_25644_, _22768_, _22762_);
  and (_25645_, _25644_, _25642_);
  or (_26865_, _25645_, _25619_);
  and (_25646_, _25571_, _23778_);
  and (_25647_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_17981_, _25647_, _25646_);
  and (_25649_, _24010_, _23076_);
  and (_25650_, _25649_, _23649_);
  not (_25651_, _25649_);
  and (_25652_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_18188_, _25652_, _25650_);
  and (_25653_, _25571_, _23898_);
  and (_25654_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_18303_, _25654_, _25653_);
  and (_25656_, _24370_, _23069_);
  and (_25657_, _25656_, _23946_);
  not (_25659_, _25656_);
  and (_25660_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_18519_, _25660_, _25657_);
  not (_25661_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_25662_, _24626_, _25661_);
  not (_25663_, _24560_);
  and (_25664_, _25663_, _25662_);
  nand (_25665_, _24415_, _24412_);
  and (_25666_, _25665_, _24408_);
  and (_25667_, _25666_, _24554_);
  and (_25668_, _25667_, _24552_);
  and (_25669_, _25668_, _22767_);
  or (_25671_, _25669_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_25672_, _25671_, _25664_);
  or (_25674_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _22766_);
  and (_25675_, _25674_, _22762_);
  and (_26868_[2], _25675_, _25672_);
  and (_25676_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_25677_, _24128_, _23939_);
  not (_25678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_25679_, _24252_, _24256_);
  and (_25680_, _24145_, _24131_);
  and (_25681_, _24239_, _25680_);
  nand (_25682_, _25681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_25683_, _25682_, _24256_);
  nor (_25684_, _25683_, _25679_);
  nor (_25685_, _25684_, _25678_);
  and (_25686_, _25683_, _25681_);
  and (_25687_, _25014_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_25688_, _25687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_25689_, _25688_, _25679_);
  or (_25690_, _25689_, _25686_);
  or (_25691_, _25690_, _25685_);
  or (_25692_, _25691_, _24127_);
  and (_25693_, _25692_, _24166_);
  and (_25694_, _25693_, _25677_);
  or (_18600_, _25694_, _25676_);
  and (_25695_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and (_25696_, _25542_, _23778_);
  or (_27042_, _25696_, _25695_);
  nor (_25697_, _22768_, _23100_);
  and (_25698_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_25699_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_25700_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_25701_, _25700_, _25699_);
  and (_25702_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_25703_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_25704_, _25703_, _25702_);
  and (_25705_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_25706_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_25707_, _25706_, _25705_);
  and (_25708_, _25707_, _25704_);
  and (_25709_, _25708_, _25701_);
  nor (_25710_, _25709_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_25711_, _25710_, _25698_);
  nor (_25712_, _25711_, _23950_);
  nor (_25713_, _25712_, _25697_);
  nor (_26897_[7], _25713_, rst);
  and (_25714_, _25571_, _23747_);
  and (_25715_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_19421_, _25715_, _25714_);
  nor (_25716_, _22768_, _23227_);
  and (_25717_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_25718_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_25719_, _25718_, _25717_);
  and (_25720_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_25721_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_25722_, _25721_, _25720_);
  and (_25723_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_25724_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_25725_, _25724_, _25723_);
  and (_25726_, _25725_, _25722_);
  and (_25727_, _25726_, _25719_);
  and (_25728_, _22768_, _23839_);
  not (_25729_, _25728_);
  nor (_25730_, _25729_, _25727_);
  nor (_25731_, _25730_, _25716_);
  nor (_26887_[4], _25731_, rst);
  and (_25733_, _23986_, _23076_);
  and (_25734_, _25733_, _23649_);
  not (_25735_, _25733_);
  and (_25736_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_19920_, _25736_, _25734_);
  and (_25737_, _23946_, _23755_);
  and (_25738_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  or (_19941_, _25738_, _25737_);
  and (_25739_, _23903_, _23754_);
  and (_25740_, _25739_, _23946_);
  not (_25741_, _25739_);
  and (_25742_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or (_19972_, _25742_, _25740_);
  and (_25743_, _25571_, _23649_);
  and (_25744_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_20043_, _25744_, _25743_);
  and (_25745_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  and (_25746_, _25542_, _23824_);
  or (_20570_, _25746_, _25745_);
  and (_25748_, _23784_, _23664_);
  and (_25749_, _25748_, _23898_);
  not (_25750_, _25748_);
  and (_25751_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_27069_, _25751_, _25749_);
  and (_25752_, _24050_, _23790_);
  and (_25753_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  or (_27253_, _25753_, _25752_);
  and (_25754_, _24356_, _23784_);
  and (_25755_, _25754_, _23898_);
  not (_25756_, _25754_);
  and (_25757_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or (_21247_, _25757_, _25755_);
  and (_25759_, _25754_, _23747_);
  and (_25760_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  or (_21348_, _25760_, _25759_);
  and (_25761_, _25754_, _23824_);
  and (_25762_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  or (_21419_, _25762_, _25761_);
  and (_26860_[4], _24464_, _22762_);
  and (_25763_, _24766_, _24005_);
  not (_25764_, _25763_);
  and (_25765_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_25766_, _25763_, _23946_);
  or (_21820_, _25766_, _25765_);
  and (_26885_[0], _24408_, _22762_);
  and (_26885_[1], _24417_, _22762_);
  and (_26885_[2], _24440_, _22762_);
  and (_25769_, _23052_, _22971_);
  and (_25770_, _25171_, _24069_);
  and (_25772_, _25770_, _25769_);
  and (_25773_, _25772_, _23662_);
  not (_25774_, _25773_);
  and (_25775_, _25774_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_25776_, _25769_, _23662_);
  and (_25777_, _25776_, _25770_);
  and (_25779_, _25777_, _23738_);
  nor (_25780_, _25779_, _25775_);
  nor (_26885_[3], _25780_, rst);
  or (_25782_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  not (_25783_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nand (_25784_, _23953_, _25783_);
  and (_25785_, _25784_, _22762_);
  and (_26903_[0], _25785_, _25782_);
  or (_25787_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  not (_25788_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand (_25789_, _23953_, _25788_);
  and (_25790_, _25789_, _22762_);
  and (_26903_[1], _25790_, _25787_);
  or (_25791_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  not (_25793_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand (_25794_, _23953_, _25793_);
  and (_25795_, _25794_, _22762_);
  and (_26903_[2], _25795_, _25791_);
  or (_25797_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  not (_25798_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand (_25799_, _23953_, _25798_);
  and (_25801_, _25799_, _22762_);
  and (_26903_[3], _25801_, _25797_);
  or (_25802_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  not (_25803_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand (_25804_, _23953_, _25803_);
  and (_25805_, _25804_, _22762_);
  and (_26903_[4], _25805_, _25802_);
  or (_25806_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  not (_25807_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand (_25808_, _23953_, _25807_);
  and (_25809_, _25808_, _22762_);
  and (_26903_[5], _25809_, _25806_);
  or (_25810_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  not (_25811_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand (_25812_, _23953_, _25811_);
  and (_25813_, _25812_, _22762_);
  and (_26903_[6], _25813_, _25810_);
  or (_25816_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  not (_25817_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nand (_25818_, _23953_, _25817_);
  and (_25820_, _25818_, _22762_);
  and (_26903_[7], _25820_, _25816_);
  or (_25821_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not (_25822_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_25823_, _23953_, _25822_);
  and (_25824_, _25823_, _22762_);
  and (_26903_[8], _25824_, _25821_);
  or (_25825_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  not (_25826_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_25827_, _23953_, _25826_);
  and (_25828_, _25827_, _22762_);
  and (_26903_[9], _25828_, _25825_);
  or (_25829_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  not (_25830_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_25831_, _23953_, _25830_);
  and (_25832_, _25831_, _22762_);
  and (_26903_[10], _25832_, _25829_);
  or (_25833_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  not (_25834_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_25835_, _23953_, _25834_);
  and (_25836_, _25835_, _22762_);
  and (_26903_[11], _25836_, _25833_);
  or (_25837_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  not (_25838_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand (_25839_, _23953_, _25838_);
  and (_25840_, _25839_, _22762_);
  and (_26903_[12], _25840_, _25837_);
  or (_25841_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  not (_25842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_25843_, _23953_, _25842_);
  and (_25844_, _25843_, _22762_);
  and (_26903_[13], _25844_, _25841_);
  or (_25845_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  not (_25846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_25847_, _23953_, _25846_);
  and (_25848_, _25847_, _22762_);
  and (_26903_[14], _25848_, _25845_);
  or (_25849_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  not (_25850_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_25851_, _23953_, _25850_);
  and (_25852_, _25851_, _22762_);
  and (_26903_[15], _25852_, _25849_);
  or (_25853_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  not (_25854_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_25855_, _23953_, _25854_);
  and (_25856_, _25855_, _22762_);
  and (_26903_[16], _25856_, _25853_);
  or (_25857_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  not (_25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_25859_, _23953_, _25858_);
  and (_25860_, _25859_, _22762_);
  and (_26903_[17], _25860_, _25857_);
  or (_25861_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  not (_25862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_25863_, _23953_, _25862_);
  and (_25864_, _25863_, _22762_);
  and (_26903_[18], _25864_, _25861_);
  or (_25865_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  not (_25866_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_25867_, _23953_, _25866_);
  and (_25868_, _25867_, _22762_);
  and (_26903_[19], _25868_, _25865_);
  or (_25869_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  not (_25870_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand (_25871_, _23953_, _25870_);
  and (_25873_, _25871_, _22762_);
  and (_26903_[20], _25873_, _25869_);
  or (_25875_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  not (_25876_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_25877_, _23953_, _25876_);
  and (_25878_, _25877_, _22762_);
  and (_26903_[21], _25878_, _25875_);
  or (_25879_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  not (_25880_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_25881_, _23953_, _25880_);
  and (_25882_, _25881_, _22762_);
  and (_26903_[22], _25882_, _25879_);
  or (_25883_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  not (_25884_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand (_25885_, _23953_, _25884_);
  and (_25886_, _25885_, _22762_);
  and (_26903_[23], _25886_, _25883_);
  and (_25887_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  not (_25888_, _23953_);
  and (_25889_, _25888_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or (_25890_, _25889_, _25887_);
  and (_26903_[24], _25890_, _22762_);
  or (_25891_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  not (_25892_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_25893_, _23953_, _25892_);
  and (_25894_, _25893_, _22762_);
  and (_26903_[25], _25894_, _25891_);
  or (_25895_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  not (_25896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_25897_, _23953_, _25896_);
  and (_25898_, _25897_, _22762_);
  and (_26903_[26], _25898_, _25895_);
  or (_25899_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  not (_25900_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_25901_, _23953_, _25900_);
  and (_25902_, _25901_, _22762_);
  and (_26903_[27], _25902_, _25899_);
  or (_25903_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  not (_25904_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand (_25905_, _23953_, _25904_);
  and (_25906_, _25905_, _22762_);
  and (_26903_[28], _25906_, _25903_);
  or (_25907_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  not (_25908_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_25909_, _23953_, _25908_);
  and (_25910_, _25909_, _22762_);
  and (_26903_[29], _25910_, _25907_);
  or (_25911_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  not (_25912_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand (_25913_, _23953_, _25912_);
  and (_25914_, _25913_, _22762_);
  and (_26903_[30], _25914_, _25911_);
  and (_25915_, _25754_, _24050_);
  and (_25916_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or (_22542_, _25916_, _25915_);
  and (_25917_, _25774_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_25918_, _25777_, _23642_);
  nor (_25919_, _25918_, _25917_);
  nor (_25920_, _25919_, _22971_);
  and (_25921_, _25919_, _22971_);
  nor (_25922_, _25921_, _25920_);
  nor (_25923_, _24408_, _23018_);
  and (_25924_, _24408_, _23018_);
  nor (_25925_, _25924_, _25923_);
  and (_25926_, _22905_, _22948_);
  and (_25927_, _25926_, _23052_);
  and (_25928_, _25927_, _24066_);
  and (_25929_, _25928_, _23073_);
  and (_25930_, _25929_, _25925_);
  and (_25931_, _25780_, _23003_);
  nor (_25932_, _25780_, _23003_);
  nor (_25933_, _25932_, _25931_);
  and (_25934_, _25933_, _25930_);
  and (_25935_, _25934_, _25922_);
  and (_25936_, _25780_, _24408_);
  and (_25937_, _25936_, _25919_);
  and (_25938_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_25939_, _25780_, _24612_);
  and (_25940_, _25939_, _25919_);
  and (_25941_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_25942_, _25941_, _25938_);
  nor (_25943_, _25780_, _24612_);
  and (_25945_, _25943_, _25919_);
  and (_25946_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_25947_, _25780_, _24408_);
  and (_25948_, _25947_, _25919_);
  and (_25949_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_25950_, _25949_, _25946_);
  and (_25952_, _25950_, _25942_);
  not (_25953_, _25919_);
  and (_25954_, _25947_, _25953_);
  and (_25955_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_25956_, _25943_, _25953_);
  and (_25957_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_25958_, _25957_, _25955_);
  and (_25959_, _25939_, _25953_);
  and (_25960_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_25961_, _25936_, _25953_);
  and (_25962_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_25963_, _25962_, _25960_);
  and (_25964_, _25963_, _25958_);
  and (_25965_, _25964_, _25952_);
  nor (_25966_, _25965_, _25935_);
  and (_25967_, _25935_, _24685_);
  nor (_25968_, _25967_, _25966_);
  nor (_26886_[0], _25968_, rst);
  and (_25969_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_25970_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_25971_, _25970_, _25969_);
  and (_25973_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_25974_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_25975_, _25974_, _25973_);
  and (_25976_, _25975_, _25971_);
  and (_25977_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_25978_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_25979_, _25978_, _25977_);
  and (_25980_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_25981_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_25982_, _25981_, _25980_);
  and (_25983_, _25982_, _25979_);
  and (_25984_, _25983_, _25976_);
  nor (_25985_, _25984_, _25935_);
  and (_25986_, _25935_, _23892_);
  nor (_25987_, _25986_, _25985_);
  nor (_26886_[1], _25987_, rst);
  and (_25988_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_25989_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_25990_, _25989_, _25988_);
  and (_25991_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_25992_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_25993_, _25992_, _25991_);
  and (_25994_, _25993_, _25990_);
  and (_25995_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_25996_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_25997_, _25996_, _25995_);
  and (_25998_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_26000_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_26001_, _26000_, _25998_);
  and (_26002_, _26001_, _25997_);
  and (_26003_, _26002_, _25994_);
  nor (_26004_, _26003_, _25935_);
  and (_26005_, _25935_, _23816_);
  nor (_26006_, _26005_, _26004_);
  nor (_26886_[2], _26006_, rst);
  and (_26007_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_26008_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_26009_, _26008_, _26007_);
  and (_26010_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_26011_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_26012_, _26011_, _26010_);
  and (_26013_, _26012_, _26009_);
  and (_26014_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_26015_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_26016_, _26015_, _26014_);
  and (_26017_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_26018_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_26019_, _26018_, _26017_);
  and (_26020_, _26019_, _26016_);
  and (_26021_, _26020_, _26013_);
  nor (_26022_, _26021_, _25935_);
  and (_26023_, _25935_, _23738_);
  nor (_26024_, _26023_, _26022_);
  nor (_26886_[3], _26024_, rst);
  and (_26026_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_26027_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_26028_, _26027_, _26026_);
  and (_26029_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_26030_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_26031_, _26030_, _26029_);
  and (_26032_, _26031_, _26028_);
  and (_26033_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_26034_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_26035_, _26034_, _26033_);
  and (_26036_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_26037_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_26038_, _26037_, _26036_);
  and (_26039_, _26038_, _26035_);
  and (_26040_, _26039_, _26032_);
  nor (_26041_, _26040_, _25935_);
  and (_26042_, _25935_, _23642_);
  nor (_26043_, _26042_, _26041_);
  nor (_26886_[4], _26043_, rst);
  and (_26044_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_26045_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor (_26046_, _26045_, _26044_);
  and (_26047_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_26048_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_26049_, _26048_, _26047_);
  and (_26051_, _26049_, _26046_);
  and (_26052_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_26053_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_26055_, _26053_, _26052_);
  and (_26056_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_26058_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_26060_, _26058_, _26056_);
  and (_26061_, _26060_, _26055_);
  and (_26062_, _26061_, _26051_);
  nor (_26063_, _26062_, _25935_);
  and (_26064_, _25935_, _23939_);
  nor (_26065_, _26064_, _26063_);
  nor (_26886_[5], _26065_, rst);
  and (_26067_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_26069_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_26070_, _26069_, _26067_);
  and (_26072_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_26073_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_26074_, _26073_, _26072_);
  and (_26075_, _26074_, _26070_);
  and (_26076_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_26077_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nor (_26078_, _26077_, _26076_);
  and (_26079_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_26080_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_26082_, _26080_, _26079_);
  and (_26083_, _26082_, _26078_);
  and (_26084_, _26083_, _26075_);
  nor (_26085_, _26084_, _25935_);
  and (_26086_, _25935_, _24043_);
  nor (_26088_, _26086_, _26085_);
  nor (_26886_[6], _26088_, rst);
  and (_26089_, _23824_, _23755_);
  and (_26090_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or (_22628_, _26090_, _26089_);
  and (_26091_, _25754_, _23946_);
  and (_26092_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or (_22629_, _26092_, _26091_);
  and (_26094_, _25754_, _23649_);
  and (_26095_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  or (_27034_, _26095_, _26094_);
  nand (_26096_, _24293_, _23702_);
  nor (_26097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not (_26098_, _26097_);
  not (_26099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_26100_, _26099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_26101_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not (_26102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_26103_, t0_i);
  and (_26104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _26103_);
  nor (_26105_, _26104_, _26102_);
  not (_26106_, _26105_);
  not (_26107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_26108_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_26109_, _26108_, _26107_);
  and (_26110_, _26109_, _26106_);
  and (_26111_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_26112_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_26113_, _26112_, _26111_);
  and (_26114_, _26113_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_26115_, _26114_, _26110_);
  and (_26116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_26117_, _26116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_26118_, _26117_, _26115_);
  nor (_26119_, _26118_, _26097_);
  nor (_26120_, _26119_, _26101_);
  nand (_26121_, _26120_, _26098_);
  or (_26122_, _26121_, _24299_);
  and (_26123_, _26122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_26124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand (_26125_, _26124_, _26115_);
  or (_26126_, _26125_, _26120_);
  nor (_26127_, _26126_, _24299_);
  or (_26128_, _26127_, _26123_);
  or (_26129_, _26128_, _24293_);
  and (_26130_, _26129_, _22762_);
  and (_22630_, _26130_, _26096_);
  nor (_26131_, _22768_, _23275_);
  and (_26133_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_26134_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_26135_, _26134_, _26133_);
  and (_26136_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_26137_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_26138_, _26137_, _26136_);
  and (_26139_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_26140_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_26141_, _26140_, _26139_);
  and (_26142_, _26141_, _26138_);
  and (_26143_, _26142_, _26135_);
  nor (_26144_, _26143_, _25729_);
  nor (_26145_, _26144_, _26131_);
  nor (_26887_[3], _26145_, rst);
  nor (_26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_26147_, _26146_, _23392_);
  nor (_26148_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_26149_, _26148_, _26147_);
  and (_26150_, _23397_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_26151_, _26150_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26152_, _23179_, _23141_);
  nor (_26153_, _26152_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_26154_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_26155_, _23462_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26157_, _23216_, _26156_);
  nand (_26158_, _26157_, _26155_);
  or (_26159_, _23250_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26160_, _23177_, _26156_);
  nand (_26161_, _26160_, _26159_);
  and (_26162_, _26161_, _26158_);
  or (_26163_, _23332_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26164_, _23250_, _26156_);
  nand (_26165_, _26164_, _26163_);
  or (_26166_, _23216_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_26167_, _23141_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_26168_, _26167_, _26166_);
  and (_26169_, _26168_, _26165_);
  nand (_26170_, _26169_, _26162_);
  and (_26171_, _26170_, _26154_);
  nor (_26172_, _26171_, _26153_);
  or (_26173_, _23364_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26174_, _23462_, _26156_);
  nand (_26175_, _26174_, _26173_);
  and (_26176_, _26175_, _26154_);
  and (_26177_, _26168_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_26178_, _26177_, _26176_);
  not (_26179_, _26178_);
  nor (_26180_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_26181_, _26180_);
  nand (_26182_, _26146_, _23131_);
  and (_26183_, _26182_, _26181_);
  not (_26184_, _26183_);
  or (_26185_, _23397_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26186_, _23332_, _26156_);
  and (_26187_, _26186_, _26185_);
  or (_26188_, _26187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26189_, _26161_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26190_, _26189_, _26188_);
  or (_26191_, _26190_, _26184_);
  and (_26192_, _23364_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26193_, _26192_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26194_, _26158_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26195_, _26194_, _26193_);
  nor (_26196_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_26197_, _26196_);
  nand (_26198_, _26146_, _23171_);
  and (_26199_, _26198_, _26197_);
  not (_26200_, _26199_);
  or (_26201_, _26200_, _26195_);
  nand (_26202_, _26189_, _26188_);
  or (_26203_, _26202_, _26183_);
  and (_26204_, _26203_, _26191_);
  not (_26205_, _26204_);
  or (_26206_, _26205_, _26201_);
  and (_26207_, _26206_, _26191_);
  nand (_26208_, _26194_, _26193_);
  or (_26209_, _26199_, _26208_);
  and (_26210_, _26209_, _26201_);
  and (_26211_, _26210_, _26204_);
  nor (_26212_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_26213_, _26212_);
  not (_26214_, _26146_);
  or (_26215_, _26214_, _23208_);
  nand (_26216_, _26215_, _26213_);
  or (_26217_, _26150_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26218_, _26165_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26219_, _26218_, _26217_);
  or (_26220_, _26219_, _26216_);
  nor (_26221_, _26175_, _26154_);
  nand (_26222_, _26146_, _23244_);
  nor (_26223_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_26224_, _26223_);
  and (_26225_, _26224_, _26222_);
  not (_26226_, _26225_);
  or (_26227_, _26226_, _26221_);
  and (_26228_, _26215_, _26213_);
  nand (_26229_, _26218_, _26217_);
  or (_26230_, _26229_, _26228_);
  nand (_26231_, _26230_, _26220_);
  or (_26232_, _26231_, _26227_);
  nand (_26233_, _26232_, _26220_);
  nand (_26234_, _26233_, _26211_);
  and (_26235_, _26234_, _26207_);
  and (_26236_, _26187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_26237_, _26236_);
  nor (_26238_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_26239_, _26238_);
  nand (_26240_, _26146_, _23291_);
  and (_26241_, _26240_, _26239_);
  nand (_26242_, _26241_, _26237_);
  or (_26243_, _26241_, _26237_);
  nand (_26244_, _26243_, _26242_);
  nand (_26245_, _26192_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_26246_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_26247_, _26246_);
  or (_26248_, _26214_, _23326_);
  and (_26249_, _26248_, _26247_);
  nand (_26250_, _26249_, _26245_);
  nor (_26251_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_26252_, _26251_);
  or (_26253_, _26214_, _23359_);
  nand (_26254_, _26253_, _26252_);
  and (_26255_, _26254_, _26151_);
  or (_26256_, _26249_, _26245_);
  nand (_26257_, _26256_, _26250_);
  or (_26258_, _26257_, _26255_);
  and (_26259_, _26258_, _26250_);
  or (_26260_, _26259_, _26244_);
  nand (_26261_, _26260_, _26242_);
  not (_26262_, _26221_);
  or (_26263_, _26225_, _26262_);
  and (_26264_, _26263_, _26227_);
  and (_26265_, _26230_, _26220_);
  and (_26266_, _26265_, _26264_);
  and (_26267_, _26266_, _26211_);
  nand (_26268_, _26267_, _26261_);
  nand (_26269_, _26268_, _26235_);
  and (_26270_, _26179_, _26172_);
  nand (_26271_, _26270_, _26269_);
  and (_26272_, _26271_, _26184_);
  not (_26273_, _26272_);
  and (_26274_, _26270_, _26269_);
  and (_26275_, _26219_, _26216_);
  not (_26276_, _26227_);
  and (_26277_, _26264_, _26261_);
  nor (_26278_, _26277_, _26276_);
  or (_26279_, _26278_, _26275_);
  and (_26280_, _26279_, _26220_);
  not (_26281_, _26280_);
  nand (_26282_, _26281_, _26210_);
  nand (_26283_, _26282_, _26201_);
  nand (_26284_, _26283_, _26205_);
  nand (_26285_, _26284_, _26274_);
  and (_26286_, _26285_, _26273_);
  and (_26287_, _26286_, _26179_);
  nor (_26288_, _26286_, _26179_);
  or (_26289_, _26281_, _26210_);
  nand (_26290_, _26289_, _26282_);
  nand (_26291_, _26290_, _26274_);
  and (_26292_, _26271_, _26200_);
  not (_26293_, _26292_);
  and (_26294_, _26293_, _26291_);
  nand (_26295_, _26294_, _26202_);
  nor (_26296_, _26295_, _26288_);
  nor (_26297_, _26296_, _26287_);
  or (_26298_, _26288_, _26287_);
  or (_26299_, _26294_, _26202_);
  and (_26300_, _26299_, _26295_);
  not (_26301_, _26300_);
  nor (_26302_, _26301_, _26298_);
  nand (_26303_, _26231_, _26278_);
  or (_26304_, _26231_, _26278_);
  nand (_26305_, _26304_, _26303_);
  nand (_26306_, _26305_, _26274_);
  and (_26307_, _26271_, _26216_);
  not (_26308_, _26307_);
  and (_26309_, _26308_, _26306_);
  and (_26310_, _26309_, _26208_);
  nor (_26311_, _26264_, _26261_);
  or (_26312_, _26311_, _26277_);
  and (_26313_, _26312_, _26274_);
  and (_26314_, _26271_, _26226_);
  nor (_26315_, _26314_, _26313_);
  and (_26316_, _26315_, _26229_);
  not (_26317_, _26316_);
  nor (_26318_, _26309_, _26208_);
  or (_26319_, _26318_, _26310_);
  nor (_26320_, _26319_, _26317_);
  nor (_26321_, _26320_, _26310_);
  and (_26322_, _26259_, _26244_);
  not (_26323_, _26322_);
  and (_26324_, _26323_, _26260_);
  or (_26325_, _26324_, _26271_);
  or (_26326_, _26274_, _26241_);
  and (_26327_, _26326_, _26325_);
  nor (_26328_, _26327_, _26262_);
  not (_26329_, _26328_);
  not (_26330_, _26151_);
  or (_26331_, _26271_, _26330_);
  nand (_26332_, _26331_, _26254_);
  or (_26333_, _26331_, _26254_);
  and (_26334_, _26333_, _26332_);
  nand (_26335_, _26334_, _26245_);
  or (_26336_, _26334_, _26245_);
  and (_26337_, _26336_, _26335_);
  nor (_26338_, _26330_, _26149_);
  not (_26339_, _26338_);
  nand (_26340_, _26339_, _26337_);
  and (_26341_, _26340_, _26335_);
  and (_26342_, _26257_, _26255_);
  not (_26343_, _26342_);
  and (_26344_, _26343_, _26258_);
  or (_26345_, _26344_, _26271_);
  or (_26346_, _26274_, _26249_);
  and (_26347_, _26346_, _26345_);
  nand (_26348_, _26347_, _26237_);
  or (_26349_, _26347_, _26237_);
  and (_26350_, _26349_, _26348_);
  not (_26351_, _26350_);
  or (_26352_, _26351_, _26341_);
  and (_26353_, _26327_, _26262_);
  not (_26354_, _26353_);
  and (_26355_, _26354_, _26348_);
  nand (_26356_, _26355_, _26352_);
  and (_26357_, _26356_, _26329_);
  nor (_26358_, _26315_, _26229_);
  nor (_26359_, _26358_, _26316_);
  not (_26360_, _26359_);
  nor (_26361_, _26319_, _26360_);
  nand (_26362_, _26361_, _26357_);
  nand (_26363_, _26362_, _26321_);
  nand (_26364_, _26363_, _26302_);
  nand (_26365_, _26364_, _26297_);
  and (_26366_, _26365_, _26172_);
  nand (_26367_, _26366_, _26151_);
  and (_26368_, _26367_, _26149_);
  nor (_26369_, _26367_, _26149_);
  or (_26370_, _26369_, _26368_);
  nand (_26371_, _26370_, _23599_);
  nor (_26372_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_26373_, _26372_);
  and (_26374_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  not (_26375_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _26375_);
  not (_26377_, _26376_);
  or (_26378_, _26377_, _23296_);
  not (_26379_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_26380_, _26379_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_26381_, _26380_);
  or (_26383_, _26381_, _23214_);
  and (_26384_, _26383_, _26378_);
  or (_26385_, _26380_, _26376_);
  or (_26386_, _26385_, _23400_);
  and (_26387_, _26386_, _26373_);
  and (_26388_, _26387_, _26384_);
  and (_26389_, _26372_, _23141_);
  nor (_26390_, _26389_, _26388_);
  and (_26391_, _26390_, _23359_);
  or (_26392_, _26377_, _23404_);
  or (_26393_, _26381_, _23263_);
  and (_26394_, _26393_, _26392_);
  or (_26395_, _26385_, _23418_);
  and (_26396_, _26395_, _26373_);
  nand (_26397_, _26396_, _26394_);
  or (_26398_, _26373_, _23177_);
  and (_26399_, _26398_, _26397_);
  and (_26400_, _26399_, _23326_);
  nand (_26401_, _26400_, _26391_);
  and (_26402_, _26399_, _23616_);
  nand (_26403_, _26398_, _26397_);
  or (_26404_, _26403_, _23612_);
  and (_26405_, _26390_, _23326_);
  and (_26406_, _26405_, _26404_);
  nand (_26407_, _26406_, _26402_);
  nand (_26408_, _26407_, _26401_);
  or (_26409_, _26389_, _26388_);
  or (_26410_, _26409_, _23291_);
  or (_26411_, _26403_, _23244_);
  or (_26412_, _26411_, _26410_);
  nand (_26413_, _26411_, _26410_);
  and (_26414_, _26413_, _26412_);
  and (_26415_, _26414_, _26408_);
  and (_26416_, _26390_, _23525_);
  and (_26417_, _26416_, _26402_);
  or (_26418_, _26409_, _23522_);
  or (_26419_, _26418_, _26411_);
  and (_26420_, _26399_, _23208_);
  or (_26421_, _26420_, _26416_);
  and (_26422_, _26421_, _26419_);
  nand (_26423_, _26422_, _26417_);
  or (_26424_, _26422_, _26417_);
  and (_26425_, _26424_, _26423_);
  nand (_26426_, _26425_, _26415_);
  not (_26427_, _26418_);
  or (_26428_, _26419_, _23171_);
  and (_26429_, _26399_, _24028_);
  not (_26430_, _26429_);
  nand (_26431_, _26430_, _26419_);
  and (_26432_, _26431_, _26428_);
  nand (_26433_, _26432_, _26427_);
  or (_26434_, _26429_, _26427_);
  nand (_26435_, _26434_, _26433_);
  or (_26436_, _26435_, _26426_);
  or (_26437_, _26409_, _23392_);
  nor (_26438_, _26437_, _26404_);
  or (_26439_, _26400_, _26391_);
  and (_26440_, _26439_, _26401_);
  and (_26441_, _26440_, _26438_);
  or (_26442_, _26406_, _26402_);
  and (_26443_, _26442_, _26407_);
  and (_26444_, _26443_, _26441_);
  nand (_26445_, _26414_, _26408_);
  or (_26446_, _26414_, _26408_);
  and (_26447_, _26446_, _26445_);
  and (_26448_, _26447_, _26444_);
  or (_26449_, _26425_, _26415_);
  and (_26450_, _26449_, _26426_);
  nand (_26451_, _26450_, _26448_);
  not (_26452_, _26451_);
  and (_26453_, _26426_, _26423_);
  nand (_26454_, _26453_, _26435_);
  or (_26455_, _26453_, _26435_);
  and (_26456_, _26455_, _26454_);
  nand (_26457_, _26456_, _26452_);
  nand (_26458_, _26457_, _26436_);
  nor (_26459_, _26435_, _26423_);
  not (_26460_, _26428_);
  and (_26461_, _26432_, _26427_);
  or (_26462_, _26403_, _23131_);
  or (_26463_, _26409_, _23171_);
  or (_26464_, _26463_, _26462_);
  nand (_26465_, _26463_, _26462_);
  and (_26466_, _26465_, _26464_);
  nand (_26467_, _26466_, _26461_);
  or (_26468_, _26466_, _26461_);
  and (_26469_, _26468_, _26467_);
  nand (_26470_, _26469_, _26460_);
  or (_26471_, _26469_, _26460_);
  and (_26472_, _26471_, _26470_);
  nand (_26473_, _26472_, _26459_);
  or (_26474_, _26472_, _26459_);
  and (_26475_, _26474_, _26473_);
  nand (_26476_, _26475_, _26458_);
  or (_26477_, _26475_, _26458_);
  and (_26478_, _26477_, _26476_);
  nand (_26479_, _26478_, _26374_);
  or (_26480_, _26478_, _26374_);
  and (_26481_, _26480_, _26479_);
  and (_26482_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or (_26483_, _26456_, _26452_);
  and (_26484_, _26483_, _26457_);
  nand (_26485_, _26484_, _26482_);
  or (_26486_, _26484_, _26482_);
  nand (_26487_, _26486_, _26485_);
  and (_26488_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or (_26489_, _26450_, _26448_);
  and (_26490_, _26489_, _26451_);
  nand (_26491_, _26490_, _26488_);
  or (_26492_, _26490_, _26488_);
  and (_26493_, _26492_, _26491_);
  and (_26494_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nand (_26495_, _26447_, _26444_);
  or (_26496_, _26447_, _26444_);
  and (_26497_, _26496_, _26495_);
  nand (_26498_, _26497_, _26494_);
  and (_26499_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nand (_26500_, _26443_, _26441_);
  or (_26501_, _26443_, _26441_);
  and (_26502_, _26501_, _26500_);
  nand (_26503_, _26502_, _26499_);
  and (_26504_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand (_26505_, _26440_, _26438_);
  or (_26506_, _26440_, _26438_);
  and (_26507_, _26506_, _26505_);
  and (_26508_, _26507_, _26504_);
  not (_26509_, _26508_);
  or (_26510_, _26502_, _26499_);
  nand (_26511_, _26510_, _26503_);
  or (_26512_, _26511_, _26509_);
  nand (_26513_, _26512_, _26503_);
  or (_26514_, _26497_, _26494_);
  and (_26515_, _26514_, _26498_);
  nand (_26516_, _26515_, _26513_);
  nand (_26517_, _26516_, _26498_);
  nand (_26518_, _26517_, _26493_);
  and (_26519_, _26518_, _26491_);
  or (_26520_, _26519_, _26487_);
  nand (_26521_, _26520_, _26485_);
  nand (_26522_, _26521_, _26481_);
  nand (_26523_, _26522_, _26479_);
  and (_26524_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  nand (_26525_, _26476_, _26473_);
  and (_26526_, _26390_, _23536_);
  and (_26527_, _26526_, _26430_);
  and (_26528_, _26470_, _26467_);
  not (_26529_, _26528_);
  nand (_26530_, _26529_, _26527_);
  or (_26531_, _26529_, _26527_);
  and (_26532_, _26531_, _26530_);
  nand (_26533_, _26532_, _26525_);
  or (_26534_, _26532_, _26525_);
  and (_26535_, _26534_, _26533_);
  nand (_26536_, _26535_, _26524_);
  or (_26537_, _26535_, _26524_);
  and (_26538_, _26537_, _26536_);
  and (_26539_, _26538_, _26523_);
  nor (_26540_, _26538_, _26523_);
  nor (_26541_, _26540_, _26539_);
  and (_26542_, _26541_, _23596_);
  and (_26543_, _23521_, _23422_);
  nor (_26544_, _26543_, _23492_);
  and (_26545_, _26544_, _23087_);
  not (_26546_, _26545_);
  and (_26547_, _23480_, _26544_);
  and (_26548_, _23571_, _23456_);
  not (_26549_, _26548_);
  nand (_26550_, _23602_, _23359_);
  and (_26551_, _23582_, _23536_);
  and (_26552_, _23579_, _23567_);
  nor (_26553_, _26552_, _26551_);
  or (_26554_, _23539_, _23392_);
  and (_26555_, _26554_, _23767_);
  and (_26556_, _26555_, _23764_);
  and (_26557_, _26556_, _26553_);
  and (_26558_, _26557_, _26550_);
  nand (_26559_, _26558_, _26549_);
  nor (_26560_, _26559_, _26547_);
  and (_26561_, _26560_, _23760_);
  and (_26562_, _26561_, _26546_);
  not (_26563_, _26562_);
  nor (_26564_, _26563_, _26542_);
  nand (_26565_, _26564_, _26371_);
  and (_26566_, _24566_, _24542_);
  and (_26567_, _24616_, _24613_);
  and (_26568_, _25666_, _24446_);
  nor (_26569_, _26568_, _26567_);
  nor (_26570_, _26569_, _24382_);
  nor (_26571_, _26566_, _26570_);
  not (_26572_, _24382_);
  and (_26573_, _26567_, _26572_);
  not (_26574_, _26573_);
  and (_26575_, _24593_, _24567_);
  and (_26576_, _26575_, _26572_);
  nor (_26577_, _26576_, _24628_);
  and (_26578_, _26577_, _26574_);
  not (_26579_, _24566_);
  nor (_26580_, _25630_, _26579_);
  and (_26581_, _25667_, _24618_);
  and (_26582_, _24554_, _25665_);
  and (_26583_, _24606_, _26582_);
  or (_26584_, _26583_, _26581_);
  and (_26585_, _24440_, _24417_);
  and (_26586_, _24538_, _24553_);
  and (_26587_, _26586_, _26585_);
  and (_26588_, _26587_, _24535_);
  and (_26589_, _24538_, _24445_);
  and (_26590_, _26589_, _24535_);
  or (_26591_, _26590_, _26588_);
  or (_26592_, _26591_, _26584_);
  and (_26593_, _26592_, _24566_);
  nor (_26594_, _26593_, _26580_);
  nand (_26595_, _26594_, _26578_);
  and (_26596_, _26575_, _24471_);
  nor (_26597_, _26596_, _25629_);
  and (_26598_, _24606_, _24445_);
  or (_26599_, _26598_, _24607_);
  and (_26600_, _26589_, _24584_);
  nor (_26601_, _26600_, _26599_);
  nand (_26602_, _26601_, _26597_);
  nor (_26603_, _25620_, _24542_);
  not (_26604_, _26603_);
  or (_26605_, _26604_, _26584_);
  or (_26606_, _26605_, _26602_);
  and (_26607_, _26606_, _24566_);
  or (_26608_, _26576_, _24569_);
  or (_26609_, _26608_, _26607_);
  nor (_26610_, _26609_, _26595_);
  and (_26611_, _26610_, _26571_);
  or (_26612_, _26611_, _26566_);
  and (_26613_, _26612_, _26565_);
  and (_26614_, _24616_, _24471_);
  and (_26615_, _26614_, _25667_);
  and (_26616_, _24596_, _24535_);
  or (_26618_, _26616_, _26615_);
  and (_26619_, _25667_, _24606_);
  and (_26620_, _24604_, _24447_);
  and (_26621_, _24584_, _24567_);
  or (_26622_, _26621_, _26620_);
  or (_26623_, _26622_, _26619_);
  or (_26624_, _26623_, _26618_);
  and (_26625_, _24471_, _24445_);
  and (_26626_, _26625_, _24535_);
  or (_26627_, _26626_, _24614_);
  or (_26628_, _24593_, _24589_);
  and (_26629_, _25667_, _26628_);
  or (_26630_, _25638_, _24546_);
  and (_26631_, _26630_, _25667_);
  or (_26632_, _26631_, _26629_);
  or (_26633_, _26632_, _26627_);
  not (_26634_, _26597_);
  and (_26635_, _24613_, _24536_);
  and (_26636_, _25633_, _24612_);
  or (_26637_, _26636_, _26635_);
  or (_26638_, _26637_, _26634_);
  or (_26639_, _26638_, _26633_);
  or (_26640_, _26639_, _26624_);
  and (_26641_, _24606_, _24567_);
  or (_26643_, _26581_, _26641_);
  and (_26644_, _24613_, _24541_);
  and (_26645_, _24616_, _24538_);
  and (_26646_, _26645_, _25667_);
  or (_26647_, _26646_, _26644_);
  or (_26648_, _26647_, _26643_);
  and (_26650_, _24588_, _24471_);
  and (_26651_, _25667_, _26650_);
  and (_26652_, _24567_, _24536_);
  or (_26653_, _26652_, _26651_);
  and (_26654_, _26650_, _24447_);
  or (_26655_, _25621_, _24606_);
  and (_26656_, _26655_, _24613_);
  or (_26657_, _26656_, _26654_);
  or (_26658_, _26657_, _26653_);
  or (_26659_, _26658_, _26648_);
  and (_26660_, _24613_, _24552_);
  and (_26661_, _24589_, _24447_);
  or (_26662_, _26661_, _26660_);
  and (_26663_, _25667_, _24604_);
  and (_26665_, _25621_, _25667_);
  or (_26666_, _26665_, _26663_);
  and (_26668_, _24613_, _24546_);
  or (_26669_, _25668_, _26668_);
  or (_26670_, _26669_, _26666_);
  or (_26671_, _26670_, _26662_);
  or (_26672_, _26671_, _26659_);
  or (_26673_, _26672_, _26640_);
  nand (_26674_, _26673_, _26572_);
  nor (_26675_, _24628_, _24569_);
  nand (_26676_, _26675_, _26674_);
  nand (_26677_, _26676_, _22766_);
  and (_26678_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_26679_, _26678_);
  and (_26680_, _26679_, _26677_);
  nor (_26681_, _26680_, _24634_);
  and (_26682_, _26681_, _24576_);
  and (_26683_, _24067_, _23002_);
  and (_26684_, _26683_, _24077_);
  not (_26685_, _26684_);
  nor (_26686_, _26685_, _23702_);
  and (_26687_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_26688_, _26684_, _23738_);
  nor (_26689_, _26688_, _26687_);
  and (_26691_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_26692_, _26684_, _23816_);
  or (_26693_, _26692_, _26691_);
  nand (_26694_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nand (_26695_, _26684_, _23892_);
  and (_26696_, _26695_, _26694_);
  or (_26697_, _26684_, _23012_);
  nand (_26698_, _26684_, _24685_);
  and (_26699_, _26698_, _26697_);
  and (_26700_, _26699_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_26701_, _26700_, _26696_);
  not (_26702_, _26701_);
  nor (_26703_, _26702_, _26693_);
  and (_26704_, _26703_, _26689_);
  and (_26705_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_26707_, _26684_, _23642_);
  nor (_26708_, _26707_, _26705_);
  and (_26709_, _26708_, _26704_);
  and (_26710_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_26711_, _26684_, _23939_);
  nor (_26712_, _26711_, _26710_);
  and (_26713_, _26712_, _26709_);
  and (_26714_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_26715_, _26684_, _24043_);
  nor (_26716_, _26715_, _26714_);
  and (_26717_, _26716_, _26713_);
  and (_26718_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and (_26719_, _26718_, _26717_);
  nor (_26721_, _26718_, _26717_);
  or (_26722_, _26721_, _22920_);
  or (_26723_, _26722_, _26719_);
  and (_26724_, _26723_, _22924_);
  nor (_26725_, _26724_, _26684_);
  or (_26727_, _26725_, _26686_);
  nand (_26728_, _26727_, _26682_);
  not (_26729_, _24634_);
  and (_26730_, _26680_, _26729_);
  and (_26732_, _26730_, _24576_);
  nand (_26733_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand (_26734_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_26735_, _26734_, _26733_);
  nand (_26736_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand (_26737_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_26738_, _26737_, _26736_);
  and (_26739_, _26738_, _26735_);
  nand (_26740_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand (_26741_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_26742_, _26741_, _26740_);
  nand (_26743_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nand (_26744_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_26745_, _26744_, _26743_);
  and (_26746_, _26745_, _26742_);
  and (_26747_, _26746_, _26739_);
  nor (_26749_, _26747_, _25935_);
  not (_26750_, _23702_);
  and (_26751_, _25935_, _26750_);
  or (_26752_, _26751_, _26749_);
  nand (_26753_, _26752_, _26732_);
  nor (_26754_, _26680_, _26729_);
  nor (_26755_, _22768_, _23104_);
  and (_26756_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_26757_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_26758_, _26757_, _26756_);
  and (_26759_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_26760_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_26761_, _26760_, _26759_);
  and (_26762_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_26763_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_26765_, _26763_, _26762_);
  and (_26766_, _26765_, _26761_);
  and (_26767_, _26766_, _26758_);
  nor (_26768_, _26767_, _25729_);
  nor (_26770_, _26768_, _26755_);
  not (_26772_, _26770_);
  nand (_26773_, _26772_, _26754_);
  and (_26775_, _26773_, _24576_);
  and (_26776_, _26775_, _26753_);
  nand (_26777_, _26776_, _26728_);
  and (_26778_, _26777_, _22943_);
  nor (_26779_, _26777_, _22943_);
  nor (_26781_, _26779_, _26778_);
  not (_26782_, _26682_);
  nor (_26783_, _26716_, _26713_);
  nor (_26784_, _26783_, _26717_);
  nor (_26785_, _26784_, _22920_);
  nor (_26786_, _26785_, _23025_);
  nor (_26787_, _26786_, _26684_);
  nor (_26788_, _26787_, _26715_);
  nor (_26789_, _26788_, _26782_);
  not (_26790_, _26789_);
  not (_26791_, _26732_);
  nor (_26792_, _26088_, _26791_);
  not (_26793_, _26792_);
  and (_26794_, _24634_, _24577_);
  and (_26795_, _26681_, _24577_);
  nor (_26796_, _26795_, _26794_);
  nor (_26797_, _22768_, _23154_);
  and (_26798_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_26799_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_26800_, _26799_, _26798_);
  and (_26801_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_26802_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_26803_, _26802_, _26801_);
  and (_26804_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_26806_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_26807_, _26806_, _26804_);
  and (_26808_, _26807_, _26803_);
  and (_26809_, _26808_, _26800_);
  nor (_26810_, _26809_, _25729_);
  nor (_26811_, _26810_, _26797_);
  not (_26812_, _26811_);
  and (_26813_, _26812_, _26754_);
  not (_26814_, _26813_);
  and (_26815_, _26814_, _26796_);
  and (_26816_, _26815_, _26793_);
  and (_26817_, _26816_, _26790_);
  nor (_26818_, _26817_, _23034_);
  and (_26819_, _26817_, _23034_);
  nor (_26820_, _26819_, _26818_);
  nor (_26821_, _26712_, _26709_);
  nor (_26822_, _26821_, _26713_);
  nor (_26823_, _26822_, _22920_);
  nor (_26824_, _26823_, _23044_);
  nor (_26825_, _26824_, _26684_);
  nor (_26826_, _26825_, _26711_);
  nor (_26827_, _26826_, _26782_);
  not (_26829_, _26827_);
  nor (_26830_, _26065_, _26791_);
  not (_26831_, _26830_);
  and (_26832_, _26754_, _24576_);
  nor (_26833_, _22768_, _23191_);
  and (_26835_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_26836_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_26837_, _26836_, _26835_);
  and (_26838_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_26839_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_26840_, _26839_, _26838_);
  and (_26841_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00001_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_00002_, _00001_, _26841_);
  and (_00003_, _00002_, _26840_);
  and (_00004_, _00003_, _26837_);
  nor (_00005_, _00004_, _25729_);
  nor (_00006_, _00005_, _26833_);
  not (_00007_, _00006_);
  and (_00008_, _00007_, _26832_);
  not (_00009_, _00008_);
  and (_00010_, _26794_, _26680_);
  nor (_00011_, _26795_, _00010_);
  and (_00012_, _00011_, _00009_);
  and (_00013_, _00012_, _26831_);
  and (_00014_, _00013_, _26829_);
  nor (_00015_, _00014_, _23052_);
  and (_00016_, _00014_, _23052_);
  nor (_00017_, _00016_, _00015_);
  nor (_00018_, _26024_, _26791_);
  not (_00019_, _26145_);
  and (_00020_, _26832_, _00019_);
  nor (_00021_, _00020_, _00018_);
  not (_00022_, _26689_);
  or (_00023_, _26702_, _26693_);
  and (_00024_, _00023_, _00022_);
  nor (_00025_, _00024_, _26704_);
  nor (_00026_, _00025_, _22920_);
  nor (_00027_, _00026_, _22990_);
  nor (_00028_, _00027_, _26684_);
  nor (_00029_, _00028_, _26688_);
  not (_00030_, _00029_);
  and (_00031_, _00030_, _26682_);
  and (_00032_, _24634_, _24576_);
  and (_00033_, _00032_, _26680_);
  not (_00034_, _00033_);
  nor (_00035_, _00034_, _25780_);
  nor (_00036_, _00035_, _00031_);
  and (_00037_, _00036_, _00021_);
  nor (_00038_, _00037_, _23002_);
  and (_00039_, _00037_, _23002_);
  nor (_00040_, _00039_, _00038_);
  nor (_00041_, _26708_, _26704_);
  nor (_00042_, _00041_, _26709_);
  nor (_00043_, _00042_, _22920_);
  nor (_00044_, _00043_, _22954_);
  nor (_00045_, _00044_, _26684_);
  nor (_00046_, _00045_, _26707_);
  not (_00047_, _00046_);
  and (_00048_, _00047_, _26682_);
  not (_00049_, _00048_);
  nor (_00050_, _26043_, _26791_);
  not (_00051_, _25731_);
  and (_00052_, _26754_, _00051_);
  not (_00053_, _00052_);
  and (_00054_, _00033_, _25953_);
  nor (_00055_, _00054_, _26794_);
  nand (_00056_, _00055_, _00053_);
  nor (_00057_, _00056_, _00050_);
  and (_00058_, _00057_, _00049_);
  nor (_00059_, _00058_, _22970_);
  and (_00060_, _00058_, _22970_);
  nor (_00061_, _00060_, _00059_);
  or (_00062_, _00061_, _00040_);
  or (_00063_, _00062_, _00017_);
  or (_00064_, _00063_, _26820_);
  nor (_00065_, _00064_, _26781_);
  nor (_00066_, _25987_, _26791_);
  nor (_00067_, _24634_, _24576_);
  and (_00068_, _00032_, _24417_);
  or (_00069_, _00068_, _00067_);
  and (_00070_, _00069_, _26680_);
  nor (_00071_, _26700_, _26696_);
  nor (_00072_, _00071_, _26701_);
  nor (_00073_, _00072_, _22920_);
  nor (_00074_, _00073_, _22975_);
  nor (_00075_, _00074_, _26684_);
  not (_00076_, _00075_);
  and (_00077_, _00076_, _26695_);
  not (_00078_, _00077_);
  and (_00079_, _00078_, _26682_);
  nor (_00080_, _22768_, _23343_);
  and (_00081_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00082_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_00083_, _00082_, _00081_);
  and (_00084_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00085_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_00086_, _00085_, _00084_);
  and (_00087_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00088_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_00089_, _00088_, _00087_);
  and (_00091_, _00089_, _00086_);
  and (_00092_, _00091_, _00083_);
  nor (_00093_, _00092_, _25729_);
  nor (_00094_, _00093_, _00080_);
  not (_00095_, _00094_);
  and (_00096_, _00095_, _26832_);
  or (_00097_, _00096_, _00079_);
  or (_00098_, _00097_, _00070_);
  nor (_00099_, _00098_, _00066_);
  and (_00100_, _00099_, _24289_);
  nor (_00101_, _00099_, _24289_);
  or (_00102_, _00101_, _00100_);
  not (_00103_, _00102_);
  nor (_00104_, _25968_, _26791_);
  not (_00105_, _00104_);
  nor (_00106_, _26699_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_00107_, _00106_, _26700_);
  nor (_00108_, _00107_, _22920_);
  nor (_00109_, _00108_, _23014_);
  nor (_00110_, _00109_, _26684_);
  not (_00111_, _00110_);
  and (_00112_, _00111_, _26698_);
  not (_00113_, _00112_);
  and (_00114_, _00113_, _26682_);
  nand (_00115_, _00033_, _24408_);
  nor (_00116_, _22768_, _23375_);
  and (_00117_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00118_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_00119_, _00118_, _00117_);
  and (_00120_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00121_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_00122_, _00121_, _00120_);
  and (_00123_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00124_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_00125_, _00124_, _00123_);
  and (_00126_, _00125_, _00122_);
  and (_00127_, _00126_, _00119_);
  nor (_00128_, _00127_, _25729_);
  nor (_00129_, _00128_, _00116_);
  not (_00130_, _00129_);
  nand (_00131_, _00130_, _26832_);
  nand (_00132_, _00131_, _00115_);
  nor (_00133_, _00132_, _00114_);
  and (_00134_, _00133_, _00105_);
  nor (_00135_, _00134_, _23018_);
  and (_00136_, _00134_, _23018_);
  nor (_00137_, _00136_, _00135_);
  not (_00138_, _00137_);
  nor (_00139_, _26006_, _26791_);
  not (_00140_, _00139_);
  and (_00141_, _00033_, _24440_);
  and (_00142_, _26702_, _26693_);
  nor (_00143_, _00142_, _26703_);
  nor (_00144_, _00143_, _22920_);
  nor (_00145_, _00144_, _23057_);
  nor (_00146_, _00145_, _26684_);
  nor (_00147_, _00146_, _26692_);
  not (_00148_, _00147_);
  and (_00149_, _00148_, _26682_);
  nor (_00150_, _22768_, _23322_);
  and (_00151_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00152_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_00153_, _00152_, _00151_);
  and (_00154_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00155_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_00156_, _00155_, _00154_);
  and (_00157_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00158_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_00159_, _00158_, _00157_);
  and (_00160_, _00159_, _00156_);
  and (_00161_, _00160_, _00153_);
  nor (_00162_, _00161_, _25729_);
  nor (_00163_, _00162_, _00150_);
  not (_00164_, _00163_);
  and (_00165_, _00164_, _26832_);
  or (_00166_, _00165_, _00149_);
  nor (_00167_, _00166_, _00141_);
  and (_00168_, _00167_, _00140_);
  nor (_00169_, _00168_, _23065_);
  and (_00170_, _00168_, _23065_);
  nor (_00171_, _00170_, _00169_);
  nor (_00172_, _00171_, _25181_);
  and (_00173_, _00172_, _00138_);
  and (_00174_, _00173_, _00103_);
  and (_00175_, _00174_, _00065_);
  and (_00176_, _22943_, _22948_);
  and (_00177_, _00176_, _00175_);
  not (_00178_, _00177_);
  nor (_00179_, _26597_, _26579_);
  nor (_00180_, _26597_, _24382_);
  nor (_00181_, _00180_, _00179_);
  not (_00182_, _00181_);
  nor (_00183_, _24654_, _24070_);
  and (_00184_, _00183_, _00065_);
  and (_00185_, _00184_, _00182_);
  and (_00186_, _23471_, _23483_);
  nor (_00187_, _23471_, _23483_);
  nor (_00188_, _00187_, _00186_);
  not (_00189_, _00188_);
  nor (_00190_, _23469_, _23259_);
  nor (_00191_, _00190_, _23470_);
  nor (_00192_, _23468_, _23262_);
  nor (_00193_, _00192_, _23469_);
  nor (_00194_, _23467_, _23266_);
  and (_00195_, _23467_, _23266_);
  nor (_00196_, _00195_, _00194_);
  not (_00197_, _00196_);
  and (_00198_, _23460_, _23411_);
  nor (_00199_, _00198_, _23461_);
  nor (_00201_, _26544_, _23416_);
  nor (_00202_, _23458_, _23414_);
  nor (_00204_, _00202_, _23459_);
  and (_00205_, _00204_, _00201_);
  and (_00207_, _00205_, _00199_);
  not (_00208_, _24569_);
  and (_00209_, _00181_, _00208_);
  and (_00210_, _00209_, _00207_);
  and (_00211_, _00210_, _00197_);
  and (_00212_, _00211_, _00193_);
  and (_00213_, _00212_, _00191_);
  and (_00214_, _00213_, _00189_);
  nor (_00215_, _00181_, _23561_);
  not (_00216_, _00215_);
  and (_00217_, _00181_, _24534_);
  nor (_00218_, _00217_, _00208_);
  and (_00219_, _00218_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_00220_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_00221_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_00222_, _00221_, _00220_);
  nor (_00223_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_00224_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_00225_, _00224_, _00223_);
  and (_00226_, _00225_, _00222_);
  and (_00227_, _00226_, _24630_);
  nor (_00228_, _00227_, _00219_);
  and (_00229_, _00228_, _00216_);
  not (_00230_, _00229_);
  nor (_00231_, _00230_, _00214_);
  nor (_00232_, _26600_, _26584_);
  not (_00233_, _24567_);
  and (_00234_, _24593_, _24538_);
  or (_00235_, _24589_, _24541_);
  nor (_00236_, _00235_, _00234_);
  nor (_00237_, _00236_, _00233_);
  nor (_00238_, _00237_, _26591_);
  and (_00239_, _00238_, _00232_);
  not (_00240_, _00239_);
  and (_00241_, _00240_, _00231_);
  and (_00242_, _26603_, _24615_);
  not (_00243_, _00242_);
  nor (_00244_, _00243_, _00241_);
  nand (_00245_, _25629_, _24544_);
  and (_00246_, _24568_, _24471_);
  nor (_00247_, _00246_, _26596_);
  and (_00248_, _00247_, _00245_);
  or (_00249_, _00248_, _00231_);
  and (_00250_, _00249_, _00244_);
  nor (_00251_, _24628_, _24566_);
  nor (_00252_, _00251_, _00250_);
  nor (_00253_, _00252_, _26570_);
  not (_00254_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_00255_, _22766_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_00256_, _00255_, _00254_);
  not (_00257_, _00256_);
  not (_00258_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_00259_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _22766_);
  and (_00260_, _00259_, _00258_);
  and (_00261_, _24733_, _23662_);
  and (_00262_, _00261_, _25770_);
  nor (_00263_, _00262_, _00260_);
  and (_00264_, _00263_, _00257_);
  nor (_00265_, _23052_, _23034_);
  and (_00266_, _00265_, _24645_);
  and (_00267_, _00266_, _25259_);
  not (_00268_, _00267_);
  and (_00270_, _00268_, _00264_);
  not (_00271_, _00270_);
  and (_00272_, _00271_, _24630_);
  nor (_00273_, _23053_, _23034_);
  and (_00274_, _00273_, _24645_);
  and (_00276_, _00274_, _25163_);
  nor (_00277_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_00278_, _00277_);
  nor (_00280_, _00278_, _00276_);
  and (_00281_, _00280_, _25774_);
  not (_00282_, _00281_);
  and (_00283_, _00282_, _00218_);
  nor (_00284_, _00283_, _00272_);
  not (_00285_, _00284_);
  nor (_00286_, _00285_, _00253_);
  not (_00287_, _00286_);
  nor (_00288_, _00287_, _00185_);
  and (_00289_, _00288_, _00178_);
  and (_00290_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  not (_00291_, _25566_);
  and (_00292_, _26573_, _00291_);
  and (_00293_, _24567_, _26572_);
  and (_00294_, _00293_, _24593_);
  nor (_00295_, _26591_, _24568_);
  and (_00297_, _00295_, _26603_);
  and (_00298_, _00297_, _25630_);
  and (_00300_, _00298_, _00232_);
  nor (_00301_, _00300_, _26579_);
  nor (_00302_, _00301_, _00294_);
  not (_00303_, _26571_);
  and (_00304_, _26594_, _26578_);
  and (_00305_, _00304_, _00303_);
  and (_00306_, _00305_, _00302_);
  and (_00307_, _00306_, _00130_);
  or (_00308_, _00307_, _00292_);
  or (_00310_, _00308_, _00290_);
  and (_00311_, _26595_, _00291_);
  and (_00312_, _00304_, _00130_);
  or (_00313_, _00312_, _00311_);
  nor (_00314_, _00313_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_00315_, _00313_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_00316_, _00315_, _00314_);
  nor (_00317_, _00305_, _00302_);
  and (_00318_, _00317_, _00316_);
  nor (_00319_, _00318_, _00310_);
  nand (_00320_, _00319_, _00289_);
  or (_00321_, _00320_, _26613_);
  or (_00322_, _00289_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00323_, _00322_, _22762_);
  and (_26890_[0], _00323_, _00321_);
  not (_00324_, _26536_);
  nor (_00325_, _26539_, _00324_);
  and (_00326_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  and (_00327_, _26530_, _26464_);
  nand (_00328_, _00327_, _26533_);
  nand (_00329_, _00328_, _00326_);
  or (_00330_, _00328_, _00326_);
  nand (_00331_, _00330_, _00329_);
  or (_00332_, _00331_, _00325_);
  nand (_00333_, _00331_, _00325_);
  and (_00334_, _00333_, _00332_);
  nand (_00335_, _00334_, _23596_);
  nand (_00336_, _26365_, _26172_);
  or (_00337_, _26339_, _26337_);
  and (_00338_, _00337_, _26340_);
  or (_00339_, _00338_, _00336_);
  or (_00340_, _26366_, _26334_);
  and (_00341_, _00340_, _00339_);
  nand (_00342_, _00341_, _23599_);
  nor (_00343_, _23419_, _23367_);
  or (_00344_, _00343_, _23485_);
  and (_00345_, _00344_, _23492_);
  nor (_00346_, _00344_, _23492_);
  or (_00347_, _00346_, _00345_);
  and (_00348_, _00347_, _23480_);
  nor (_00349_, _23457_, _23417_);
  nor (_00350_, _00349_, _23458_);
  nor (_00351_, _00350_, _23088_);
  nor (_00352_, _00351_, _00348_);
  nor (_00353_, _23530_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_00354_, _00353_, _23359_);
  nor (_00355_, _00353_, _23359_);
  nor (_00356_, _00355_, _00354_);
  nor (_00357_, _00356_, _23539_);
  not (_00358_, _00357_);
  not (_00359_, _23604_);
  nor (_00360_, _00359_, _23392_);
  not (_00361_, _00360_);
  nand (_00362_, _23602_, _23326_);
  and (_00363_, _23579_, _23359_);
  not (_00364_, _00363_);
  and (_00365_, _00364_, _00362_);
  and (_00366_, _00365_, _00361_);
  and (_00367_, _00366_, _23889_);
  and (_00368_, _00367_, _00358_);
  and (_00369_, _00368_, _23878_);
  and (_00370_, _00369_, _00352_);
  and (_00371_, _00370_, _00342_);
  and (_00372_, _00371_, _00335_);
  not (_00373_, _00372_);
  and (_00374_, _00373_, _26612_);
  nor (_00375_, _22768_, _23341_);
  and (_00376_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_00377_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00378_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00379_, _00378_, _00377_);
  and (_00380_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00381_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_00382_, _00381_, _00380_);
  or (_00383_, _00382_, _00379_);
  and (_00384_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00386_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00387_, _00386_, _00384_);
  or (_00388_, _00387_, _00383_);
  and (_00389_, _00388_, _23839_);
  or (_00390_, _00389_, _00376_);
  and (_00391_, _00390_, _22768_);
  nor (_00392_, _00391_, _00375_);
  or (_00393_, _00392_, _00304_);
  or (_00394_, _26595_, _00094_);
  and (_00395_, _00394_, _00393_);
  or (_00396_, _00395_, _23336_);
  nand (_00397_, _00395_, _23336_);
  and (_00398_, _00397_, _00396_);
  and (_00399_, _00398_, _00315_);
  not (_00400_, _00305_);
  and (_00401_, _00400_, _26609_);
  or (_00402_, _00398_, _00315_);
  nand (_00403_, _00402_, _00401_);
  or (_00404_, _00403_, _00399_);
  and (_00405_, _26610_, _00303_);
  and (_00406_, _00405_, _00095_);
  nor (_00407_, _00392_, _26574_);
  and (_00408_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00409_, _00408_, _00407_);
  nor (_00410_, _00409_, _00406_);
  and (_00411_, _00410_, _00404_);
  nand (_00412_, _00411_, _00289_);
  or (_00413_, _00412_, _00374_);
  or (_00414_, _00289_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00415_, _00414_, _22762_);
  and (_26890_[1], _00415_, _00413_);
  not (_00416_, _00289_);
  not (_00417_, _26352_);
  and (_00418_, _26351_, _26341_);
  nor (_00419_, _00418_, _00417_);
  or (_00420_, _00419_, _00336_);
  or (_00421_, _26366_, _26347_);
  and (_00422_, _00421_, _00420_);
  nand (_00423_, _00422_, _23599_);
  and (_00424_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  nand (_00425_, _00332_, _00329_);
  nand (_00426_, _00425_, _00424_);
  or (_00427_, _00425_, _00424_);
  and (_00428_, _00427_, _00426_);
  nand (_00429_, _00428_, _23596_);
  nor (_00430_, _00204_, _23088_);
  or (_00431_, _23603_, _23291_);
  and (_00432_, _23579_, _23326_);
  not (_00433_, _00432_);
  nand (_00434_, _23604_, _23359_);
  and (_00435_, _00434_, _00433_);
  and (_00436_, _00435_, _00431_);
  and (_00437_, _00436_, _23811_);
  not (_00438_, _00437_);
  nor (_00439_, _00438_, _00430_);
  nor (_00440_, _23495_, _23493_);
  nor (_00441_, _00440_, _23481_);
  and (_00442_, _00441_, _23497_);
  and (_00443_, _23529_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_00444_, _00355_, _23610_);
  nor (_00445_, _00444_, _00443_);
  nor (_00446_, _00445_, _23539_);
  nor (_00447_, _00446_, _00442_);
  and (_00448_, _00447_, _00439_);
  and (_00449_, _00448_, _23803_);
  and (_00450_, _00449_, _00429_);
  nand (_00451_, _00450_, _00423_);
  and (_00452_, _00451_, _26612_);
  and (_00453_, _00405_, _00164_);
  nor (_00454_, _22768_, _23302_);
  and (_00455_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_00456_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00457_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00458_, _00457_, _00456_);
  and (_00459_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00460_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_00461_, _00460_, _00459_);
  or (_00462_, _00461_, _00458_);
  and (_00463_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00464_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00465_, _00464_, _00463_);
  or (_00466_, _00465_, _00462_);
  and (_00467_, _00466_, _23839_);
  or (_00468_, _00467_, _00455_);
  and (_00469_, _00468_, _22768_);
  nor (_00470_, _00469_, _00454_);
  not (_00471_, _00470_);
  and (_00472_, _00471_, _26573_);
  and (_00473_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_00474_, _00473_, _00472_);
  or (_00475_, _00474_, _00453_);
  not (_00476_, _00396_);
  or (_00477_, _00399_, _00476_);
  and (_00478_, _00471_, _26595_);
  and (_00479_, _00304_, _00164_);
  nor (_00480_, _00479_, _00478_);
  nor (_00481_, _00480_, _23307_);
  and (_00482_, _00480_, _23307_);
  nor (_00483_, _00482_, _00481_);
  or (_00484_, _00483_, _00477_);
  and (_00485_, _00483_, _00477_);
  not (_00486_, _00485_);
  and (_00487_, _00486_, _00317_);
  and (_00488_, _00487_, _00484_);
  or (_00489_, _00488_, _00475_);
  or (_00490_, _00489_, _00452_);
  or (_00491_, _00490_, _00416_);
  not (_00492_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00493_, _23953_, _00492_);
  and (_00494_, _23953_, _00492_);
  nor (_00495_, _00494_, _00493_);
  or (_00496_, _00495_, _00289_);
  and (_00497_, _00496_, _22762_);
  and (_26890_[2], _00497_, _00491_);
  or (_00498_, _00331_, _26536_);
  nand (_00499_, _00498_, _00329_);
  and (_00500_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_00501_, _00500_, _00424_);
  and (_00502_, _00501_, _00499_);
  and (_00503_, _00330_, _00329_);
  and (_00504_, _00503_, _26538_);
  and (_00505_, _00501_, _00504_);
  and (_00506_, _00505_, _26523_);
  or (_00507_, _00506_, _00502_);
  not (_00508_, _00507_);
  not (_00509_, _00500_);
  nand (_00510_, _00509_, _00426_);
  and (_00511_, _00510_, _00508_);
  nand (_00512_, _00511_, _23596_);
  or (_00513_, _26353_, _26328_);
  and (_00514_, _26352_, _26348_);
  or (_00515_, _00514_, _00513_);
  nand (_00516_, _00514_, _00513_);
  nand (_00517_, _00516_, _00515_);
  nand (_00518_, _00517_, _26366_);
  or (_00519_, _26366_, _26327_);
  and (_00520_, _00519_, _00518_);
  nand (_00521_, _00520_, _23599_);
  nor (_00522_, _00199_, _23088_);
  not (_00523_, _00522_);
  and (_00524_, _23497_, _23491_);
  or (_00525_, _00524_, _23481_);
  nor (_00526_, _00525_, _23498_);
  not (_00527_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_00528_, _23529_, _00527_);
  nor (_00529_, _00528_, _23616_);
  and (_00530_, _23579_, _23616_);
  nor (_00531_, _23530_, _23539_);
  nor (_00532_, _00531_, _00530_);
  nor (_00533_, _00532_, _00529_);
  not (_00534_, _00533_);
  or (_00535_, _23603_, _23244_);
  nand (_00536_, _23604_, _23326_);
  and (_00537_, _00536_, _00535_);
  and (_00538_, _00537_, _23736_);
  and (_00539_, _00538_, _00534_);
  and (_00540_, _00539_, _23725_);
  not (_00541_, _00540_);
  nor (_00542_, _00541_, _00526_);
  and (_00543_, _00542_, _00523_);
  and (_00544_, _00543_, _00521_);
  nand (_00545_, _00544_, _00512_);
  and (_00546_, _00545_, _26612_);
  and (_00547_, _00405_, _00019_);
  and (_00548_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00549_, _22768_, _23273_);
  and (_00550_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_00551_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00552_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_00553_, _00552_, _00551_);
  and (_00554_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00555_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_00556_, _00555_, _00554_);
  and (_00557_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00558_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_00559_, _00558_, _00557_);
  and (_00560_, _00559_, _00556_);
  and (_00561_, _00560_, _00553_);
  nor (_00563_, _00561_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_00564_, _00563_, _00550_);
  nor (_00565_, _00564_, _23950_);
  nor (_00566_, _00565_, _00549_);
  not (_00567_, _00566_);
  and (_00568_, _00567_, _26573_);
  or (_00569_, _00568_, _00548_);
  or (_00570_, _00569_, _00547_);
  or (_00571_, _00485_, _00481_);
  and (_00572_, _00567_, _26595_);
  and (_00573_, _00304_, _00019_);
  nor (_00574_, _00573_, _00572_);
  nor (_00575_, _00574_, _23268_);
  and (_00576_, _00574_, _23268_);
  nor (_00577_, _00576_, _00575_);
  nand (_00578_, _00577_, _00571_);
  or (_00579_, _00577_, _00571_);
  and (_00580_, _00579_, _00578_);
  and (_00581_, _00580_, _00317_);
  or (_00582_, _00581_, _00570_);
  or (_00583_, _00582_, _00546_);
  and (_00584_, _00583_, _00289_);
  and (_00585_, _00493_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00586_, _00493_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00587_, _00586_, _00585_);
  and (_00588_, _00587_, _00416_);
  or (_00589_, _00588_, _00584_);
  and (_26890_[3], _00589_, _22762_);
  nand (_00590_, _26359_, _26357_);
  or (_00591_, _26359_, _26357_);
  and (_00592_, _00591_, _00590_);
  or (_00593_, _00592_, _00336_);
  or (_00594_, _26366_, _26315_);
  and (_00595_, _00594_, _00593_);
  and (_00596_, _00595_, _23599_);
  and (_00597_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_00598_, _00597_, _00507_);
  nor (_00599_, _00597_, _00507_);
  nor (_00600_, _00599_, _00598_);
  and (_00601_, _00600_, _23596_);
  and (_00602_, _00196_, _23087_);
  or (_00603_, _23501_, _23266_);
  nor (_00604_, _23502_, _23481_);
  and (_00605_, _00604_, _00603_);
  or (_00606_, _23531_, _23525_);
  nor (_00607_, _23532_, _23539_);
  and (_00608_, _00607_, _00606_);
  and (_00609_, _23602_, _23208_);
  and (_00610_, _23579_, _23525_);
  nor (_00611_, _00359_, _23291_);
  or (_00612_, _00611_, _00610_);
  or (_00613_, _00612_, _00609_);
  or (_00614_, _00613_, _00608_);
  or (_00615_, _00614_, _23641_);
  or (_00616_, _00615_, _00605_);
  or (_00618_, _00616_, _00602_);
  or (_00619_, _00618_, _00601_);
  or (_00620_, _00619_, _00596_);
  and (_00621_, _00620_, _26612_);
  and (_00622_, _00405_, _00051_);
  nor (_00623_, _22768_, _23225_);
  and (_00624_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_00625_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00627_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_00628_, _00627_, _00625_);
  and (_00629_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00630_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_00631_, _00630_, _00629_);
  and (_00632_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00633_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_00634_, _00633_, _00632_);
  and (_00635_, _00634_, _00631_);
  and (_00636_, _00635_, _00628_);
  nor (_00637_, _00636_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_00638_, _00637_, _00624_);
  nor (_00639_, _00638_, _23950_);
  nor (_00640_, _00639_, _00623_);
  not (_00641_, _00640_);
  and (_00642_, _00641_, _26573_);
  and (_00643_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00644_, _00643_, _00642_);
  or (_00645_, _00644_, _00622_);
  and (_00646_, _00641_, _26595_);
  and (_00647_, _00304_, _00051_);
  nor (_00648_, _00647_, _00646_);
  or (_00649_, _00648_, _23220_);
  nand (_00650_, _00648_, _23220_);
  and (_00651_, _00650_, _00649_);
  nor (_00652_, _00575_, _00571_);
  nor (_00653_, _00652_, _00576_);
  or (_00654_, _00653_, _00651_);
  nand (_00655_, _00653_, _00651_);
  and (_00656_, _00655_, _00317_);
  and (_00657_, _00656_, _00654_);
  nor (_00658_, _00657_, _00645_);
  nand (_00659_, _00658_, _00289_);
  or (_00660_, _00659_, _00621_);
  and (_00661_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_00662_, _00661_, _00493_);
  nor (_00663_, _00585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00664_, _00663_, _00662_);
  or (_00665_, _00664_, _00289_);
  and (_00666_, _00665_, _22762_);
  and (_26890_[4], _00666_, _00660_);
  and (_00667_, _00590_, _26317_);
  nand (_00668_, _26319_, _00667_);
  or (_00669_, _26319_, _00667_);
  and (_00670_, _00669_, _00668_);
  or (_00671_, _00670_, _00336_);
  or (_00672_, _26366_, _26309_);
  and (_00673_, _00672_, _00671_);
  and (_00674_, _00673_, _23599_);
  and (_00675_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_00676_, _00675_, _00597_);
  nand (_00677_, _00676_, _00507_);
  or (_00678_, _00675_, _00598_);
  and (_00679_, _00678_, _00677_);
  and (_00680_, _00679_, _23596_);
  nor (_00681_, _23264_, _23219_);
  nor (_00682_, _00681_, _23506_);
  or (_00683_, _00682_, _23502_);
  nor (_00684_, _23503_, _23481_);
  and (_00685_, _00684_, _00683_);
  nor (_00686_, _00193_, _23088_);
  and (_00687_, _23532_, _23208_);
  nor (_00688_, _23532_, _23208_);
  nor (_00689_, _23523_, _23131_);
  nor (_00690_, _00689_, _23531_);
  and (_00691_, _00690_, _23521_);
  or (_00692_, _00691_, _00688_);
  or (_00693_, _00692_, _00687_);
  and (_00694_, _00691_, _23522_);
  nor (_00695_, _00694_, _23539_);
  and (_00696_, _00695_, _00693_);
  and (_00697_, _23579_, _23208_);
  nor (_00698_, _00359_, _23244_);
  nor (_00699_, _23603_, _23171_);
  or (_00700_, _00699_, _00698_);
  nor (_00701_, _00700_, _00697_);
  nand (_00702_, _00701_, _23935_);
  nor (_00703_, _00702_, _00696_);
  nand (_00704_, _00703_, _23926_);
  or (_00705_, _00704_, _00686_);
  or (_00706_, _00705_, _00685_);
  or (_00707_, _00706_, _00680_);
  or (_00708_, _00707_, _00674_);
  and (_00709_, _00708_, _26612_);
  nand (_00710_, _00655_, _00649_);
  nor (_00711_, _22768_, _23188_);
  and (_00712_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_00713_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00714_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_00715_, _00714_, _00713_);
  and (_00716_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00717_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_00718_, _00717_, _00716_);
  and (_00719_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_00720_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_00721_, _00720_, _00719_);
  and (_00722_, _00721_, _00718_);
  and (_00723_, _00722_, _00715_);
  nor (_00724_, _00723_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_00725_, _00724_, _00712_);
  nor (_00726_, _00725_, _23950_);
  nor (_00727_, _00726_, _00711_);
  nor (_00728_, _00727_, _00304_);
  and (_00729_, _00304_, _00007_);
  nor (_00730_, _00729_, _00728_);
  nor (_00731_, _00730_, _23183_);
  and (_00732_, _00730_, _23183_);
  nor (_00733_, _00732_, _00731_);
  or (_00734_, _00733_, _00710_);
  and (_00735_, _00733_, _00710_);
  not (_00736_, _00735_);
  and (_00737_, _00736_, _00401_);
  nand (_00738_, _00737_, _00734_);
  nand (_00739_, _00405_, _00007_);
  and (_00741_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_00742_, _00728_, _26570_);
  nor (_00743_, _00742_, _00741_);
  and (_00744_, _00743_, _00739_);
  and (_00745_, _00744_, _00738_);
  nand (_00746_, _00745_, _00289_);
  or (_00747_, _00746_, _00709_);
  nor (_00748_, _00662_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_00749_, _00662_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00750_, _00749_, _00748_);
  or (_00751_, _00750_, _00289_);
  and (_00752_, _00751_, _22762_);
  and (_26890_[5], _00752_, _00747_);
  not (_00753_, _23599_);
  and (_00754_, _26363_, _26300_);
  nor (_00755_, _26363_, _26300_);
  or (_00756_, _00755_, _00754_);
  and (_00757_, _00756_, _26366_);
  nor (_00758_, _26366_, _26294_);
  or (_00759_, _00758_, _00757_);
  or (_00760_, _00759_, _00753_);
  and (_00761_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  not (_00762_, _00761_);
  nor (_00763_, _00762_, _00677_);
  and (_00765_, _00762_, _00677_);
  or (_00766_, _00765_, _00763_);
  or (_00767_, _00766_, _23597_);
  nor (_00768_, _00191_, _23088_);
  not (_00769_, _00768_);
  nor (_00770_, _23511_, _23503_);
  nor (_00771_, _00770_, _23481_);
  and (_00772_, _00771_, _23514_);
  and (_00773_, _24041_, _24026_);
  not (_00774_, _00688_);
  nor (_00775_, _00694_, _00774_);
  nor (_00776_, _00775_, _24028_);
  not (_00777_, _00776_);
  and (_00778_, _00775_, _24028_);
  nor (_00779_, _00778_, _23539_);
  and (_00780_, _00779_, _00777_);
  nand (_00781_, _23604_, _23208_);
  or (_00782_, _23603_, _23131_);
  and (_00783_, _23579_, _24028_);
  not (_00784_, _00783_);
  and (_00785_, _00784_, _00782_);
  nand (_00786_, _00785_, _00781_);
  nor (_00787_, _00786_, _00780_);
  and (_00788_, _00787_, _00773_);
  not (_00789_, _00788_);
  nor (_00790_, _00789_, _00772_);
  and (_00791_, _00790_, _00769_);
  and (_00792_, _00791_, _00767_);
  and (_00793_, _00792_, _00760_);
  not (_00794_, _00793_);
  and (_00795_, _00794_, _26612_);
  and (_00796_, _00405_, _26812_);
  and (_00797_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00798_, _22768_, _23152_);
  and (_00799_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_00800_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00801_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00802_, _00801_, _00800_);
  and (_00803_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00804_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_00805_, _00804_, _00803_);
  or (_00806_, _00805_, _00802_);
  and (_00807_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00808_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00809_, _00808_, _00807_);
  or (_00810_, _00809_, _00806_);
  and (_00811_, _00810_, _23839_);
  or (_00812_, _00811_, _00799_);
  and (_00813_, _00812_, _22768_);
  nor (_00814_, _00813_, _00798_);
  not (_00815_, _00814_);
  and (_00816_, _00815_, _26573_);
  or (_00817_, _00816_, _00797_);
  or (_00818_, _00817_, _00796_);
  or (_00819_, _00735_, _00731_);
  and (_00820_, _00815_, _26595_);
  and (_00821_, _00304_, _26812_);
  nor (_00822_, _00821_, _00820_);
  or (_00823_, _00822_, _23147_);
  nand (_00824_, _00822_, _23147_);
  and (_00825_, _00824_, _00823_);
  or (_00826_, _00825_, _00819_);
  nand (_00827_, _00825_, _00819_);
  and (_00829_, _00827_, _00317_);
  and (_00830_, _00829_, _00826_);
  or (_00831_, _00830_, _00818_);
  or (_00833_, _00831_, _00795_);
  and (_00834_, _00833_, _00289_);
  and (_00835_, _00749_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00836_, _00749_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00837_, _00836_, _00835_);
  and (_00838_, _00837_, _00416_);
  or (_00839_, _00838_, _00834_);
  and (_26890_[6], _00839_, _22762_);
  or (_00840_, _26366_, _26286_);
  not (_00841_, _00754_);
  nand (_00842_, _00841_, _26295_);
  and (_00843_, _00842_, _26298_);
  or (_00844_, _00843_, _00336_);
  and (_00845_, _00844_, _00840_);
  and (_00846_, _00845_, _23599_);
  not (_00847_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  or (_00848_, _26372_, _00847_);
  nor (_00849_, _00848_, _00763_);
  and (_00850_, _00763_, _00847_);
  or (_00851_, _00850_, _00849_);
  and (_00852_, _00851_, _23596_);
  and (_00853_, _00188_, _23087_);
  nand (_00854_, _23516_, _23483_);
  and (_00855_, _23518_, _23480_);
  and (_00856_, _00855_, _00854_);
  nor (_00857_, _00691_, _23533_);
  and (_00858_, _00857_, _23131_);
  nor (_00859_, _00857_, _23131_);
  or (_00860_, _00859_, _00858_);
  and (_00861_, _00860_, _23528_);
  and (_00862_, _23568_, _23456_);
  and (_00863_, _23563_, _23567_);
  and (_00864_, _23579_, _23536_);
  nor (_00865_, _00359_, _23171_);
  or (_00866_, _00865_, _00864_);
  or (_00867_, _00866_, _00863_);
  or (_00868_, _00867_, _00862_);
  nor (_00869_, _00868_, _00861_);
  nand (_00870_, _00869_, _23701_);
  or (_00871_, _00870_, _00856_);
  or (_00872_, _00871_, _00853_);
  or (_00873_, _00872_, _00852_);
  or (_00875_, _00873_, _00846_);
  and (_00876_, _00875_, _26612_);
  and (_00877_, _00405_, _26772_);
  nor (_00878_, _26574_, _25713_);
  and (_00879_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_00880_, _00879_, _00878_);
  or (_00881_, _00880_, _00877_);
  or (_00882_, _00881_, _00876_);
  nand (_00883_, _00827_, _00823_);
  nor (_00884_, _00304_, _25713_);
  and (_00885_, _00304_, _26772_);
  nor (_00886_, _00885_, _00884_);
  nor (_00887_, _00886_, _23089_);
  and (_00888_, _00886_, _23089_);
  nor (_00889_, _00888_, _00887_);
  or (_00890_, _00889_, _00883_);
  nand (_00891_, _00889_, _00883_);
  and (_00892_, _00891_, _00890_);
  nand (_00893_, _00892_, _00317_);
  nand (_00894_, _00893_, _00289_);
  or (_00895_, _00894_, _00882_);
  nor (_00896_, _00835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_00897_, _00835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00898_, _00897_, _00896_);
  or (_00899_, _00898_, _00289_);
  and (_00900_, _00899_, _22762_);
  and (_26890_[7], _00900_, _00895_);
  and (_00901_, _26565_, _24628_);
  nor (_00902_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00903_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23370_);
  nor (_00904_, _00903_, _00902_);
  not (_00905_, _00904_);
  or (_00906_, _00905_, _23519_);
  and (_00907_, _00905_, _23519_);
  nor (_00908_, _00907_, _23481_);
  and (_00909_, _00908_, _00906_);
  nand (_00910_, _26366_, _23599_);
  nor (_00911_, _23540_, _23537_);
  and (_00912_, _00911_, _23680_);
  nor (_00913_, _00912_, _23397_);
  not (_00914_, _23609_);
  and (_00915_, _00912_, _23397_);
  or (_00916_, _00915_, _00914_);
  nor (_00917_, _00916_, _00913_);
  and (_00918_, _23579_, _23397_);
  and (_00919_, _26399_, _23567_);
  and (_00920_, _00919_, _23596_);
  and (_00922_, _23571_, _23525_);
  nor (_00923_, _23688_, _23392_);
  or (_00924_, _00923_, _00922_);
  or (_00925_, _00924_, _00920_);
  nor (_00926_, _00925_, _00918_);
  not (_00927_, _00926_);
  nor (_00928_, _00927_, _00917_);
  nand (_00929_, _00928_, _00910_);
  or (_00930_, _00929_, _00909_);
  and (_00931_, _00930_, _26566_);
  and (_00932_, _26573_, _00130_);
  not (_00933_, _24530_);
  and (_00934_, _00405_, _00933_);
  and (_00935_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_00936_, _00935_, _00934_);
  or (_00937_, _00936_, _00932_);
  or (_00938_, _00937_, _00931_);
  or (_00939_, _00938_, _00901_);
  not (_00940_, _00886_);
  not (_00941_, _00888_);
  and (_00942_, _00941_, _00883_);
  or (_00943_, _00942_, _00887_);
  nand (_00944_, _00943_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_00945_, _00943_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00946_, _00945_, _00944_);
  or (_00947_, _00946_, _00940_);
  nand (_00948_, _00946_, _00940_);
  and (_00949_, _00948_, _00947_);
  and (_00950_, _00949_, _00317_);
  or (_00951_, _00950_, _00416_);
  or (_00952_, _00951_, _00939_);
  nor (_00953_, _00897_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_00954_, _00897_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00955_, _00954_, _00953_);
  or (_00956_, _00955_, _00289_);
  and (_00957_, _00956_, _22762_);
  and (_26890_[8], _00957_, _00952_);
  not (_00958_, _26566_);
  nor (_00959_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00960_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23338_);
  nor (_00961_, _00960_, _00959_);
  not (_00962_, _00961_);
  and (_00963_, _00962_, _00906_);
  not (_00964_, _00963_);
  or (_00965_, _00962_, _00906_);
  and (_00966_, _00965_, _23480_);
  and (_00967_, _00966_, _00964_);
  not (_00968_, _00967_);
  and (_00969_, _26274_, _23599_);
  not (_00970_, _00969_);
  and (_00971_, _23579_, _23364_);
  or (_00972_, _23418_, _23131_);
  nor (_00973_, _00972_, _23678_);
  and (_00974_, _00973_, _23521_);
  and (_00975_, _23418_, _23131_);
  and (_00976_, _00975_, _23674_);
  and (_00977_, _00976_, _23456_);
  nor (_00978_, _00977_, _00974_);
  nor (_00979_, _00978_, _23400_);
  and (_00980_, _00978_, _23400_);
  or (_00981_, _00980_, _00914_);
  nor (_00982_, _00981_, _00979_);
  and (_00983_, _26437_, _26404_);
  nor (_00984_, _00983_, _26438_);
  and (_00985_, _00984_, _23596_);
  and (_00986_, _23571_, _23208_);
  and (_00987_, _23627_, _23359_);
  or (_00988_, _00987_, _00986_);
  or (_00989_, _00988_, _00985_);
  or (_00990_, _00989_, _00982_);
  nor (_00991_, _00990_, _00971_);
  and (_00992_, _00991_, _00970_);
  and (_00993_, _00992_, _00968_);
  nor (_00994_, _00993_, _00958_);
  and (_00996_, _26573_, _00095_);
  not (_00997_, _24486_);
  and (_00998_, _00405_, _00997_);
  or (_00999_, _00998_, _00996_);
  and (_01000_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_01001_, _01000_, _00999_);
  or (_01002_, _01001_, _00994_);
  nor (_01003_, _00945_, _00886_);
  nor (_01004_, _00944_, _00940_);
  nor (_01005_, _01004_, _01003_);
  nand (_01006_, _01005_, _23338_);
  or (_01007_, _01005_, _23338_);
  and (_01008_, _01007_, _00317_);
  and (_01009_, _01008_, _01006_);
  or (_01010_, _01009_, _01002_);
  not (_01011_, _24628_);
  or (_01012_, _00372_, _01011_);
  nand (_01013_, _01012_, _00289_);
  or (_01014_, _01013_, _01010_);
  and (_01015_, _00954_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_01016_, _00954_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_01017_, _01016_, _01015_);
  or (_01018_, _01017_, _00289_);
  and (_01019_, _01018_, _22762_);
  and (_26890_[9], _01019_, _01014_);
  and (_01021_, _01003_, _23338_);
  and (_01022_, _01004_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_01023_, _01022_, _01021_);
  nand (_01024_, _01023_, _23309_);
  or (_01025_, _01023_, _23309_);
  and (_01026_, _01025_, _00401_);
  and (_01027_, _01026_, _01024_);
  and (_01028_, _00451_, _24628_);
  nor (_01029_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01030_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23309_);
  nor (_01031_, _01030_, _01029_);
  not (_01032_, _01031_);
  and (_01033_, _01032_, _00965_);
  not (_01034_, _01033_);
  or (_01035_, _01032_, _00965_);
  and (_01036_, _01035_, _23480_);
  and (_01037_, _01036_, _01034_);
  not (_01038_, _01037_);
  and (_01039_, _00977_, _23400_);
  and (_01040_, _00973_, _23364_);
  and (_01041_, _01040_, _23521_);
  nor (_01042_, _01041_, _01039_);
  and (_01043_, _01042_, _23404_);
  nor (_01044_, _01042_, _23404_);
  or (_01045_, _01044_, _00914_);
  nor (_01046_, _01045_, _01043_);
  nor (_01047_, _26507_, _26504_);
  nor (_01048_, _01047_, _26508_);
  and (_01049_, _01048_, _23596_);
  nand (_01050_, _00865_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_01051_, _23627_, _23326_);
  and (_01052_, _23579_, _23332_);
  and (_01053_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or (_01054_, _01053_, _01052_);
  nor (_01055_, _01054_, _01051_);
  and (_01056_, _01055_, _01050_);
  not (_01057_, _01056_);
  nor (_01058_, _01057_, _01049_);
  not (_01059_, _01058_);
  nor (_01060_, _01059_, _01046_);
  and (_01061_, _01060_, _01038_);
  nor (_01062_, _01061_, _00958_);
  and (_01063_, _26573_, _00164_);
  not (_01064_, _24508_);
  and (_01065_, _00405_, _01064_);
  or (_01066_, _01065_, _01063_);
  and (_01067_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_01068_, _01067_, _01066_);
  nor (_01069_, _01068_, _01062_);
  nand (_01070_, _01069_, _00289_);
  or (_01071_, _01070_, _01028_);
  or (_01072_, _01071_, _01027_);
  nor (_01073_, _01015_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01074_, _01015_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01075_, _01074_, _01073_);
  or (_01076_, _01075_, _00289_);
  and (_01077_, _01076_, _22762_);
  and (_26890_[10], _01077_, _01072_);
  and (_01078_, _01074_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_01079_, _01074_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_01080_, _01079_, _01078_);
  or (_01081_, _00898_, _00837_);
  and (_01082_, _00495_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_01083_, _00955_, _00587_);
  or (_01084_, _01083_, _01082_);
  or (_01085_, _01017_, _00664_);
  or (_01086_, _01085_, _01084_);
  or (_01087_, _01075_, _00750_);
  or (_01088_, _01087_, _01086_);
  or (_01089_, _01088_, _01081_);
  and (_01090_, _01089_, _01080_);
  nor (_01091_, _01089_, _01080_);
  or (_01092_, _01091_, _01090_);
  nand (_01093_, _01092_, _00306_);
  and (_01094_, _00545_, _24628_);
  nor (_01095_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01096_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23270_);
  nor (_01097_, _01096_, _01095_);
  not (_01098_, _01097_);
  and (_01099_, _01098_, _01035_);
  nor (_01100_, _01098_, _01035_);
  nor (_01101_, _01100_, _01099_);
  and (_01102_, _01101_, _23480_);
  not (_01103_, _01102_);
  and (_01105_, _26511_, _26509_);
  not (_01106_, _01105_);
  and (_01107_, _01106_, _26512_);
  and (_01108_, _01107_, _23596_);
  not (_01109_, _01108_);
  and (_01110_, _01040_, _23332_);
  nor (_01111_, _01110_, _23456_);
  and (_01112_, _23400_, _23404_);
  and (_01113_, _01112_, _00976_);
  nor (_01114_, _01113_, _23521_);
  or (_01115_, _01114_, _01111_);
  and (_01116_, _01115_, _23296_);
  nor (_01117_, _01115_, _23296_);
  nor (_01118_, _01117_, _01116_);
  and (_01119_, _01118_, _23609_);
  and (_01120_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_01121_, _23688_, _23291_);
  and (_01122_, _23579_, _23462_);
  or (_01123_, _01122_, _01121_);
  or (_01124_, _01123_, _23572_);
  nor (_01125_, _01124_, _01120_);
  not (_01126_, _01125_);
  nor (_01127_, _01126_, _01119_);
  and (_01128_, _01127_, _01109_);
  and (_01129_, _01128_, _01103_);
  nor (_01131_, _01129_, _00958_);
  and (_01132_, _26573_, _00019_);
  and (_01133_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_01134_, _01133_, _01132_);
  or (_01135_, _01134_, _01131_);
  nor (_01136_, _01135_, _01094_);
  and (_01137_, _01136_, _01093_);
  nand (_01138_, _01137_, _00289_);
  nor (_01139_, \oc8051_top_1.oc8051_memory_interface1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_01140_, _01139_, _01003_);
  nand (_01141_, \oc8051_top_1.oc8051_memory_interface1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_01142_, _01141_, _00944_);
  nor (_01143_, _01142_, _00940_);
  nor (_01144_, _01143_, _01140_);
  nand (_01145_, _01144_, _23270_);
  or (_01146_, _01144_, _23270_);
  and (_01147_, _01146_, _01145_);
  and (_01148_, _01147_, _00317_);
  or (_01149_, _01148_, _01138_);
  or (_01150_, _01080_, _00289_);
  and (_01151_, _01150_, _22762_);
  and (_26890_[11], _01151_, _01149_);
  not (_01152_, _01091_);
  and (_01153_, _01078_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_01154_, _01078_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_01155_, _01154_, _01153_);
  and (_01156_, _01155_, _01152_);
  nor (_01157_, _01155_, _01152_);
  or (_01158_, _01157_, _01156_);
  and (_01159_, _01158_, _00306_);
  and (_01160_, _00620_, _24628_);
  nor (_01161_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01162_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23222_);
  nor (_01163_, _01162_, _01161_);
  or (_01164_, _01163_, _01100_);
  and (_01165_, _01163_, _01100_);
  nor (_01166_, _01165_, _23481_);
  and (_01167_, _01166_, _01164_);
  or (_01168_, _26515_, _26513_);
  and (_01169_, _01168_, _26516_);
  and (_01170_, _01169_, _23596_);
  and (_01171_, _01113_, _23296_);
  and (_01172_, _01171_, _23456_);
  and (_01173_, _01110_, _23462_);
  and (_01174_, _01173_, _23521_);
  nor (_01175_, _01174_, _01172_);
  nand (_01176_, _01175_, _23263_);
  or (_01177_, _01175_, _23263_);
  and (_01178_, _01177_, _23609_);
  and (_01179_, _01178_, _01176_);
  and (_01180_, _23456_, _23525_);
  and (_01181_, _23521_, _23250_);
  or (_01182_, _01181_, _01180_);
  and (_01183_, _01182_, _23627_);
  and (_01184_, _23571_, _23567_);
  and (_01185_, _23579_, _23250_);
  and (_01186_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or (_01187_, _01186_, _01185_);
  or (_01188_, _01187_, _01184_);
  or (_01189_, _01188_, _01183_);
  or (_01190_, _01189_, _01179_);
  or (_01191_, _01190_, _01170_);
  or (_01192_, _01191_, _01167_);
  and (_01193_, _01192_, _26566_);
  and (_01194_, _26573_, _00051_);
  and (_01195_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_01196_, _01195_, _01194_);
  or (_01197_, _01196_, _01193_);
  or (_01198_, _01197_, _01160_);
  nor (_01199_, _01198_, _01159_);
  nand (_01200_, _01199_, _00289_);
  and (_01201_, _01139_, _23270_);
  and (_01202_, _01201_, _01003_);
  or (_01203_, _01142_, _23270_);
  nor (_01204_, _01203_, _00940_);
  nor (_01205_, _01204_, _01202_);
  nand (_01206_, _01205_, _23222_);
  or (_01207_, _01205_, _23222_);
  and (_01208_, _01207_, _01206_);
  and (_01209_, _01208_, _00317_);
  or (_01210_, _01209_, _01200_);
  or (_01211_, _01155_, _00289_);
  and (_01212_, _01211_, _22762_);
  and (_26890_[12], _01212_, _01210_);
  or (_01213_, _01203_, _23222_);
  nor (_01214_, _01213_, _00940_);
  and (_01215_, _01201_, _23222_);
  and (_01216_, _01215_, _01003_);
  nor (_01217_, _01216_, _01214_);
  nand (_01218_, _01217_, _23185_);
  or (_01219_, _01217_, _23185_);
  and (_01220_, _01219_, _00401_);
  and (_01221_, _01220_, _01218_);
  and (_01222_, _00708_, _24628_);
  nor (_01223_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01224_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23185_);
  nor (_01225_, _01224_, _01223_);
  or (_01226_, _01225_, _01165_);
  nand (_01227_, _01225_, _01165_);
  and (_01228_, _01227_, _23480_);
  and (_01229_, _01228_, _01226_);
  or (_01230_, _26517_, _26493_);
  and (_01231_, _01230_, _26518_);
  and (_01232_, _01231_, _23596_);
  and (_01233_, _23296_, _23263_);
  and (_01234_, _01233_, _01113_);
  nor (_01235_, _01234_, _23521_);
  and (_01236_, _01173_, _23250_);
  nor (_01237_, _01236_, _23456_);
  nor (_01238_, _01237_, _01235_);
  nand (_01239_, _01238_, _23216_);
  or (_01240_, _01238_, _23216_);
  and (_01241_, _01240_, _23609_);
  and (_01242_, _01241_, _01239_);
  and (_01243_, _23521_, _23216_);
  and (_01244_, _23456_, _23208_);
  or (_01245_, _01244_, _01243_);
  and (_01246_, _01245_, _23627_);
  and (_01247_, _23571_, _23359_);
  and (_01248_, _23579_, _23216_);
  and (_01249_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_01250_, _01249_, _01248_);
  or (_01251_, _01250_, _01247_);
  or (_01252_, _01251_, _01246_);
  or (_01253_, _01252_, _01242_);
  or (_01254_, _01253_, _01232_);
  or (_01255_, _01254_, _01229_);
  and (_01256_, _01255_, _26566_);
  and (_01257_, _26573_, _00007_);
  not (_01258_, _01157_);
  or (_01259_, _01153_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_01260_, _01153_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_01261_, _01260_, _01259_);
  and (_01262_, _01261_, _01258_);
  nor (_01263_, _01261_, _01258_);
  or (_01264_, _01263_, _01262_);
  and (_01265_, _01264_, _00405_);
  or (_01266_, _01265_, _01257_);
  and (_01267_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_01268_, _01267_, _01266_);
  nor (_01269_, _01268_, _01256_);
  nand (_01270_, _01269_, _00289_);
  or (_01271_, _01270_, _01222_);
  or (_01272_, _01271_, _01221_);
  or (_01273_, _01261_, _00289_);
  and (_01274_, _01273_, _22762_);
  and (_26890_[13], _01274_, _01272_);
  nor (_01275_, _00793_, _01011_);
  nor (_01276_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01278_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23149_);
  nor (_01279_, _01278_, _01276_);
  not (_01280_, _01279_);
  and (_01281_, _01280_, _01227_);
  not (_01282_, _01281_);
  or (_01283_, _01280_, _01227_);
  and (_01284_, _01283_, _23480_);
  and (_01286_, _01284_, _01282_);
  not (_01287_, _01286_);
  and (_01288_, _26519_, _26487_);
  not (_01289_, _01288_);
  and (_01290_, _01289_, _26520_);
  and (_01291_, _01290_, _23596_);
  and (_01292_, _01236_, _23216_);
  and (_01293_, _01292_, _23521_);
  and (_01294_, _01234_, _23214_);
  and (_01295_, _01294_, _23456_);
  or (_01297_, _01295_, _01293_);
  and (_01298_, _01297_, _23177_);
  nor (_01299_, _01297_, _23177_);
  nor (_01300_, _01299_, _01298_);
  and (_01301_, _01300_, _23609_);
  and (_01302_, _23521_, _23179_);
  not (_01303_, _01302_);
  and (_01304_, _23456_, _23171_);
  nor (_01305_, _01304_, _23688_);
  and (_01306_, _01305_, _01303_);
  and (_01307_, _23579_, _23177_);
  and (_01308_, _23571_, _23326_);
  and (_01309_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or (_01310_, _01309_, _01308_);
  nor (_01311_, _01310_, _01307_);
  not (_01312_, _01311_);
  nor (_01313_, _01312_, _01306_);
  not (_01314_, _01313_);
  nor (_01315_, _01314_, _01301_);
  not (_01316_, _01315_);
  nor (_01317_, _01316_, _01291_);
  and (_01318_, _01317_, _01287_);
  nor (_01319_, _01318_, _00958_);
  and (_01320_, _26573_, _26812_);
  and (_01321_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01322_, _01321_, _01320_);
  or (_01323_, _01322_, _01319_);
  or (_01324_, _01323_, _01275_);
  or (_01325_, _00945_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_01326_, _01325_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_01327_, _01326_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_01328_, _01327_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_01329_, _01328_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_01330_, _01329_, _00886_);
  or (_01331_, _01213_, _23185_);
  or (_01332_, _01331_, _00940_);
  and (_01333_, _01332_, _01330_);
  nand (_01334_, _01333_, _23149_);
  or (_01335_, _01333_, _23149_);
  and (_01336_, _01335_, _00317_);
  and (_01337_, _01336_, _01334_);
  or (_01338_, _01337_, _01324_);
  not (_01339_, _01263_);
  and (_01340_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_01341_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01342_, _01341_, _01074_);
  and (_01343_, _01342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01345_, _01342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01346_, _01345_, _01343_);
  and (_01347_, _01346_, _01339_);
  nor (_01349_, _01346_, _01339_);
  or (_01350_, _01349_, _01347_);
  nand (_01351_, _01350_, _00306_);
  nand (_01352_, _01351_, _00289_);
  or (_01353_, _01352_, _01338_);
  or (_01354_, _01346_, _00289_);
  and (_01355_, _01354_, _22762_);
  and (_26890_[14], _01355_, _01353_);
  not (_01356_, _24402_);
  not (_01357_, _24352_);
  nor (_01358_, _01357_, _23866_);
  and (_01359_, _01358_, _24436_);
  and (_01360_, _01359_, _01356_);
  nor (_01361_, _24530_, _24486_);
  and (_01362_, _01361_, _01064_);
  and (_01363_, _01362_, _01360_);
  nor (_01364_, _01064_, _24486_);
  and (_01365_, _01364_, _00933_);
  not (_01366_, _01365_);
  nor (_01367_, _24436_, _01357_);
  and (_01368_, _01367_, _23866_);
  nor (_01369_, _01368_, _01359_);
  nor (_01370_, _01369_, _01366_);
  nor (_01371_, _01370_, _01363_);
  nor (_01373_, _01371_, _24464_);
  not (_01374_, _01373_);
  nor (_01375_, _00933_, _24464_);
  and (_01376_, _01375_, _01364_);
  and (_01377_, _01368_, _24402_);
  and (_01378_, _24508_, _24486_);
  and (_01379_, _01378_, _24530_);
  and (_01380_, _01379_, _01377_);
  nor (_01381_, _01380_, _01376_);
  and (_01383_, _01359_, _24402_);
  nor (_01385_, _01383_, _01377_);
  nor (_01387_, _01385_, _01381_);
  not (_01388_, _01387_);
  not (_01389_, _01360_);
  nor (_01390_, _24508_, _24486_);
  and (_01391_, _01390_, _01375_);
  not (_01392_, _01391_);
  and (_01394_, _01064_, _24486_);
  and (_01395_, _01394_, _24530_);
  and (_01397_, _01395_, _24464_);
  nor (_01398_, _01397_, _01378_);
  and (_01399_, _01398_, _01392_);
  nor (_01400_, _01399_, _01389_);
  and (_01401_, _01368_, _01356_);
  and (_01402_, _01401_, _01376_);
  and (_01403_, _24436_, _23866_);
  and (_01404_, _24464_, _24352_);
  and (_01405_, _01404_, _01403_);
  and (_01406_, _01394_, _00933_);
  nor (_01408_, _01406_, _01365_);
  not (_01409_, _01408_);
  and (_01410_, _01409_, _01405_);
  nor (_01411_, _01410_, _01402_);
  not (_01413_, _01411_);
  nor (_01414_, _01413_, _01400_);
  and (_01415_, _01414_, _01388_);
  and (_01416_, _01415_, _01374_);
  and (_01417_, _24530_, _24464_);
  and (_01418_, _01417_, _01364_);
  and (_01420_, _01418_, _01401_);
  not (_01421_, _01420_);
  and (_01422_, _01390_, _01417_);
  and (_01423_, _01422_, _01360_);
  not (_01424_, _23866_);
  and (_01425_, _01367_, _01424_);
  and (_01426_, _01425_, _24402_);
  and (_01427_, _00933_, _24464_);
  not (_01428_, _01427_);
  not (_01429_, _01378_);
  nor (_01430_, _01429_, _01375_);
  and (_01431_, _01430_, _01428_);
  and (_01432_, _01431_, _01426_);
  and (_01433_, _01406_, _24464_);
  and (_01434_, _01433_, _01359_);
  or (_01435_, _01434_, _01432_);
  nor (_01436_, _01435_, _01423_);
  and (_01437_, _01436_, _01421_);
  not (_01439_, _01418_);
  nor (_01440_, _01377_, _01359_);
  nor (_01441_, _01440_, _01439_);
  not (_01442_, _01426_);
  and (_01443_, _24530_, _00997_);
  and (_01444_, _01443_, _01064_);
  nor (_01445_, _01444_, _01376_);
  nor (_01446_, _01433_, _01395_);
  and (_01447_, _01446_, _01445_);
  not (_01448_, _24464_);
  and (_01449_, _01406_, _01448_);
  and (_01450_, _01427_, _01378_);
  nor (_01451_, _01450_, _01418_);
  not (_01453_, _01451_);
  nor (_01454_, _01453_, _01449_);
  and (_01456_, _01454_, _01447_);
  nor (_01458_, _01456_, _01442_);
  nor (_01459_, _01458_, _01441_);
  not (_01460_, _01406_);
  and (_01461_, _01365_, _24464_);
  nor (_01462_, _01461_, _01422_);
  and (_01463_, _01462_, _01460_);
  nor (_01464_, _01463_, _24352_);
  not (_01465_, _01377_);
  nor (_01467_, _01433_, _01391_);
  and (_01468_, _01467_, _01462_);
  nor (_01469_, _01468_, _01465_);
  nor (_01470_, _01469_, _01464_);
  and (_01471_, _01470_, _01459_);
  and (_01472_, _01394_, _01375_);
  and (_01473_, _01472_, _01377_);
  and (_01474_, _01426_, _01365_);
  nor (_01475_, _01474_, _01473_);
  or (_01476_, _01449_, _01397_);
  and (_01477_, _01476_, _01377_);
  and (_01478_, _01378_, _00933_);
  not (_01479_, _01478_);
  nor (_01480_, _01461_, _01397_);
  and (_01481_, _01480_, _01479_);
  not (_01482_, _01481_);
  and (_01483_, _01482_, _01383_);
  nor (_01484_, _01483_, _01477_);
  and (_01485_, _01484_, _01475_);
  and (_01486_, _01403_, _24352_);
  and (_01487_, _01394_, _01448_);
  and (_01488_, _01487_, _01486_);
  not (_01489_, _01488_);
  and (_01490_, _01472_, _01357_);
  and (_01491_, _01425_, _01356_);
  nor (_01492_, _01491_, _01490_);
  and (_01493_, _01492_, _01489_);
  nor (_01494_, _01472_, _01461_);
  nor (_01496_, _01494_, _01389_);
  and (_01497_, _01362_, _24464_);
  nor (_01498_, _01497_, _01376_);
  nor (_01499_, _01498_, _01389_);
  nor (_01500_, _01499_, _01496_);
  and (_01501_, _01500_, _01493_);
  and (_01502_, _01501_, _01485_);
  and (_01503_, _01502_, _01471_);
  and (_01504_, _01503_, _01437_);
  and (_01505_, _01504_, _01416_);
  and (_01506_, _01365_, _01448_);
  and (_01507_, _01506_, _01401_);
  or (_01508_, _01403_, _01357_);
  and (_01509_, _01508_, _01433_);
  or (_01510_, _01509_, _01507_);
  nor (_01511_, _01510_, _01496_);
  or (_01512_, _01450_, _01397_);
  and (_01513_, _01512_, _01426_);
  or (_01514_, _01402_, _01380_);
  nor (_01515_, _01514_, _01513_);
  and (_01516_, _01515_, _01511_);
  nand (_01517_, _01516_, _01437_);
  nor (_01518_, _01517_, _01505_);
  and (_01519_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_01520_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_01522_, _01520_, _01519_);
  not (_01523_, _01522_);
  nand (_01525_, _01523_, _01518_);
  nor (_01526_, _01523_, _01518_);
  nor (_01527_, _01526_, _25729_);
  and (_01528_, _01527_, _01525_);
  nor (_01529_, _25728_, _23368_);
  or (_01530_, _01529_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01531_, _01530_, _01528_);
  not (_01532_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01533_, _01532_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_01534_, _01533_, _22762_);
  and (_26891_[0], _01534_, _01531_);
  and (_01535_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_01536_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_01537_, _01536_, _01535_);
  and (_01539_, _01537_, _01519_);
  nor (_01540_, _01537_, _01519_);
  nor (_01541_, _01540_, _01539_);
  not (_01543_, _01541_);
  nor (_01544_, _01543_, _01505_);
  and (_01545_, _01543_, _01505_);
  nor (_01546_, _01545_, _01544_);
  nand (_01547_, _01546_, _01526_);
  or (_01548_, _01546_, _01526_);
  and (_01549_, _01548_, _01547_);
  or (_01550_, _01549_, _25729_);
  or (_01551_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01552_, _01551_, _01532_);
  and (_01553_, _01552_, _01550_);
  and (_01554_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_01555_, _01554_, _01553_);
  and (_26891_[1], _01555_, _22762_);
  not (_01556_, _01544_);
  and (_01557_, _01547_, _01556_);
  not (_01558_, _01557_);
  nor (_01559_, _01539_, _01535_);
  and (_01560_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_01561_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_01562_, _01561_, _01560_);
  not (_01563_, _01562_);
  nor (_01564_, _01563_, _01559_);
  and (_01565_, _01563_, _01559_);
  nor (_01567_, _01565_, _01564_);
  and (_01568_, _01567_, _01558_);
  nor (_01569_, _01567_, _01558_);
  nor (_01570_, _01569_, _01568_);
  or (_01571_, _01570_, _25729_);
  or (_01572_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01573_, _01572_, _01532_);
  and (_01574_, _01573_, _01571_);
  and (_01575_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01576_, _01575_, _01574_);
  and (_26891_[2], _01576_, _22762_);
  nor (_01577_, _01564_, _01560_);
  nor (_01578_, _01577_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01579_, _01577_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_01580_, _01579_, _01578_);
  and (_01581_, _01580_, _01568_);
  nor (_01582_, _01580_, _01568_);
  nor (_01583_, _01582_, _01581_);
  or (_01584_, _01583_, _25729_);
  or (_01585_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01586_, _01585_, _01532_);
  and (_01587_, _01586_, _01584_);
  and (_01588_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01589_, _01588_, _01587_);
  and (_26891_[3], _01589_, _22762_);
  nor (_01590_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_01591_, _01590_, _00661_);
  nand (_01592_, _01591_, _01578_);
  or (_01593_, _01591_, _01578_);
  and (_01594_, _01593_, _01592_);
  and (_01595_, _01594_, _01581_);
  nor (_01596_, _01594_, _01581_);
  nor (_01597_, _01596_, _01595_);
  or (_01598_, _01597_, _25729_);
  or (_01599_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01600_, _01599_, _01532_);
  and (_01601_, _01600_, _01598_);
  and (_01602_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01603_, _01602_, _01601_);
  and (_26891_[4], _01603_, _22762_);
  or (_01604_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _01532_);
  and (_01605_, _01604_, _22762_);
  nand (_01606_, _01590_, _01577_);
  and (_01607_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not (_01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_01609_, _01590_, _01608_);
  and (_01610_, _01609_, _01577_);
  or (_01611_, _01610_, _01607_);
  or (_01612_, _01611_, _01595_);
  and (_01613_, _01611_, _01594_);
  and (_01614_, _01613_, _01581_);
  nor (_01615_, _01614_, _25729_);
  and (_01616_, _01615_, _01612_);
  nor (_01617_, _25728_, _23183_);
  or (_01618_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01619_, _01618_, _01616_);
  and (_26891_[5], _01619_, _01605_);
  not (_01620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_01621_, _01610_, _01620_);
  and (_01622_, _01609_, _01620_);
  and (_01623_, _01622_, _01577_);
  nor (_01624_, _01623_, _01621_);
  not (_01625_, _01624_);
  and (_01626_, _01625_, _01614_);
  or (_01627_, _01625_, _01614_);
  nand (_01628_, _01627_, _25728_);
  nor (_01629_, _01628_, _01626_);
  nor (_01630_, _25728_, _23147_);
  or (_01631_, _01630_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01632_, _01631_, _01629_);
  or (_01633_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _01532_);
  and (_01634_, _01633_, _22762_);
  and (_26891_[6], _01634_, _01632_);
  not (_01635_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_01636_, _01623_, _01635_);
  and (_01637_, _01622_, _01635_);
  and (_01638_, _01637_, _01577_);
  nor (_01639_, _01638_, _01636_);
  not (_01640_, _01639_);
  and (_01641_, _01640_, _01626_);
  nor (_01642_, _01640_, _01626_);
  nor (_01643_, _01642_, _01641_);
  or (_01644_, _01643_, _25729_);
  or (_01645_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01646_, _01645_, _01532_);
  and (_01647_, _01646_, _01644_);
  and (_01648_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_01649_, _01648_, _01647_);
  and (_26891_[7], _01649_, _22762_);
  not (_01650_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_01651_, _01638_, _01650_);
  and (_01652_, _01637_, _01650_);
  and (_01653_, _01652_, _01577_);
  or (_01654_, _01653_, _01651_);
  and (_01655_, _01654_, _01641_);
  nor (_01656_, _01654_, _01641_);
  nor (_01657_, _01656_, _01655_);
  or (_01658_, _01657_, _25729_);
  or (_01659_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01660_, _01659_, _01532_);
  and (_01661_, _01660_, _01658_);
  and (_01662_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01663_, _01662_, _01661_);
  and (_26891_[8], _01663_, _22762_);
  or (_01664_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _01532_);
  and (_01665_, _01664_, _22762_);
  not (_01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01667_, _01652_, _01666_);
  and (_01668_, _01667_, _01577_);
  nor (_01669_, _01653_, _01666_);
  nor (_01670_, _01669_, _01668_);
  not (_01671_, _01670_);
  and (_01672_, _01671_, _01655_);
  or (_01673_, _01671_, _01655_);
  nand (_01674_, _01673_, _25728_);
  nor (_01675_, _01674_, _01672_);
  nor (_01676_, _25728_, _23338_);
  or (_01677_, _01676_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01678_, _01677_, _01675_);
  and (_26891_[9], _01678_, _01665_);
  not (_01679_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01680_, _01668_, _01679_);
  and (_01681_, _01667_, _01679_);
  and (_01682_, _01681_, _01577_);
  nor (_01683_, _01682_, _01680_);
  not (_01684_, _01683_);
  and (_01685_, _01684_, _01672_);
  nor (_01686_, _01684_, _01672_);
  nor (_01687_, _01686_, _01685_);
  or (_01688_, _01687_, _25729_);
  or (_01689_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01691_, _01689_, _01532_);
  and (_01692_, _01691_, _01688_);
  and (_01693_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01695_, _01693_, _01692_);
  and (_26891_[10], _01695_, _22762_);
  not (_01697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01698_, _01681_, _01697_);
  and (_01699_, _01698_, _01577_);
  nor (_01700_, _01682_, _01697_);
  nor (_01701_, _01700_, _01699_);
  not (_01702_, _01701_);
  and (_01703_, _01702_, _01685_);
  or (_01704_, _01702_, _01685_);
  nand (_01705_, _01704_, _25728_);
  nor (_01706_, _01705_, _01703_);
  nor (_01707_, _25728_, _23270_);
  or (_01708_, _01707_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01709_, _01708_, _01706_);
  or (_01710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _01532_);
  and (_01711_, _01710_, _22762_);
  and (_26891_[11], _01711_, _01709_);
  not (_01712_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_01713_, _01699_, _01712_);
  and (_01714_, _01698_, _01712_);
  and (_01715_, _01714_, _01577_);
  nor (_01717_, _01715_, _01713_);
  not (_01718_, _01717_);
  or (_01719_, _01718_, _01703_);
  and (_01720_, _01718_, _01703_);
  nor (_01721_, _01720_, _25729_);
  and (_01722_, _01721_, _01719_);
  nor (_01723_, _25728_, _23222_);
  or (_01724_, _01723_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01725_, _01724_, _01722_);
  or (_01726_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _01532_);
  and (_01727_, _01726_, _22762_);
  and (_26891_[12], _01727_, _01725_);
  not (_01728_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01729_, _01715_, _01728_);
  and (_01730_, _01715_, _01728_);
  nor (_01731_, _01730_, _01729_);
  not (_01732_, _01731_);
  and (_01733_, _01732_, _01720_);
  nor (_01734_, _01732_, _01720_);
  nor (_01735_, _01734_, _01733_);
  or (_01736_, _01735_, _25729_);
  or (_01737_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01738_, _01737_, _01532_);
  and (_01739_, _01738_, _01736_);
  and (_01740_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_01741_, _01740_, _01739_);
  and (_26891_[13], _01741_, _22762_);
  not (_01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01743_, _01730_, _01742_);
  and (_01744_, _01730_, _01742_);
  nor (_01745_, _01744_, _01743_);
  not (_01746_, _01745_);
  and (_01747_, _01746_, _01733_);
  nor (_01748_, _01746_, _01733_);
  nor (_01749_, _01748_, _01747_);
  or (_01751_, _01749_, _25729_);
  or (_01752_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01753_, _01752_, _01532_);
  and (_01754_, _01753_, _01751_);
  and (_01755_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01756_, _01755_, _01754_);
  and (_26891_[14], _01756_, _22762_);
  nand (_01757_, _23074_, _22946_);
  and (_01758_, _23661_, _01757_);
  and (_01759_, _01758_, _24275_);
  and (_01760_, _01759_, _23946_);
  not (_01762_, _01759_);
  and (_01763_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_22631_, _01763_, _01760_);
  and (_01764_, _01759_, _23649_);
  and (_01765_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_22632_, _01765_, _01764_);
  nor (_01766_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_01767_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_01768_, _01767_, _01766_);
  nor (_01769_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor (_01770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_01771_, _01770_, _01769_);
  and (_01772_, _01771_, _01768_);
  and (_01773_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_01774_, _01773_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_26895_[0], _01774_, _22762_);
  and (_01775_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_01776_, _01775_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_26895_[1], _01776_, _22762_);
  and (_01777_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_01778_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_26895_[2], _01778_, _22762_);
  and (_01779_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_01781_, _01779_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_26895_[3], _01781_, _22762_);
  and (_01782_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_01783_, _01782_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_26895_[4], _01783_, _22762_);
  and (_01785_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_01786_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_26895_[5], _01786_, _22762_);
  and (_01787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22762_);
  and (_01788_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _22762_);
  and (_01790_, _01788_, _01772_);
  or (_26895_[6], _01790_, _01787_);
  nor (_01791_, _01518_, _23950_);
  nand (_01792_, _01791_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01793_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  or (_01794_, _01791_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_01795_, _01794_, _01793_);
  and (_26896_[0], _01795_, _01792_);
  not (_01796_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01797_, _01518_, _01796_);
  or (_01798_, _01505_, _23855_);
  nand (_01799_, _01505_, _23855_);
  and (_01800_, _01799_, _01798_);
  nand (_01801_, _01800_, _01797_);
  or (_01802_, _01800_, _01797_);
  and (_01803_, _01802_, _01801_);
  or (_01804_, _01803_, _23950_);
  or (_01805_, _22768_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01807_, _01805_, _01793_);
  and (_26896_[1], _01807_, _01804_);
  and (_01808_, _23901_, _23068_);
  and (_01809_, _23905_, _23662_);
  and (_01810_, _01809_, _01808_);
  and (_01811_, _01810_, _23747_);
  not (_01812_, _01810_);
  and (_01813_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_22633_, _01813_, _01811_);
  and (_22634_, t0_i, _22762_);
  and (_01814_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _23978_);
  and (_01815_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01816_, _01815_, _01814_);
  and (_26899_[0], _01816_, _22762_);
  and (_01817_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _23978_);
  and (_01818_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01819_, _01818_, _01817_);
  and (_26899_[1], _01819_, _22762_);
  and (_01821_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _23978_);
  and (_01822_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01823_, _01822_, _01821_);
  and (_26899_[2], _01823_, _22762_);
  and (_01824_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _23978_);
  and (_01825_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01826_, _01825_, _01824_);
  and (_26899_[3], _01826_, _22762_);
  and (_01827_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _23978_);
  and (_01828_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01829_, _01828_, _01827_);
  and (_26899_[4], _01829_, _22762_);
  and (_01830_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _23978_);
  and (_01831_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01832_, _01831_, _01830_);
  and (_26899_[5], _01832_, _22762_);
  and (_01834_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _23978_);
  and (_01835_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01836_, _01835_, _01834_);
  and (_26899_[6], _01836_, _22762_);
  and (_26902_[0], _23968_, _22762_);
  nor (_26902_[1], _23973_, rst);
  and (_26902_[2], _23976_, _22762_);
  and (_01838_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_01839_, _23953_, _25783_);
  or (_01840_, _01839_, _01838_);
  and (_26904_[0], _01840_, _22762_);
  and (_01841_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_01842_, _23953_, _25788_);
  or (_01843_, _01842_, _01841_);
  and (_26904_[1], _01843_, _22762_);
  and (_01844_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_01845_, _23953_, _25793_);
  or (_01846_, _01845_, _01844_);
  and (_26904_[2], _01846_, _22762_);
  and (_01847_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_01848_, _23953_, _25798_);
  or (_01849_, _01848_, _01847_);
  and (_26904_[3], _01849_, _22762_);
  and (_01850_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_01851_, _23953_, _25803_);
  or (_01852_, _01851_, _01850_);
  and (_26904_[4], _01852_, _22762_);
  and (_01853_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_01854_, _23953_, _25807_);
  or (_01855_, _01854_, _01853_);
  and (_26904_[5], _01855_, _22762_);
  and (_01856_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_01857_, _23953_, _25811_);
  or (_01858_, _01857_, _01856_);
  and (_26904_[6], _01858_, _22762_);
  and (_01859_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_01861_, _23953_, _25817_);
  or (_01862_, _01861_, _01859_);
  and (_26904_[7], _01862_, _22762_);
  and (_01863_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_01864_, _23953_, _25822_);
  or (_01865_, _01864_, _01863_);
  and (_26904_[8], _01865_, _22762_);
  and (_01867_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_01868_, _23953_, _25826_);
  or (_01869_, _01868_, _01867_);
  and (_26904_[9], _01869_, _22762_);
  and (_01870_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_01871_, _23953_, _25830_);
  or (_01872_, _01871_, _01870_);
  and (_26904_[10], _01872_, _22762_);
  and (_01873_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_01874_, _23953_, _25834_);
  or (_01875_, _01874_, _01873_);
  and (_26904_[11], _01875_, _22762_);
  and (_01876_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_01877_, _23953_, _25838_);
  or (_01879_, _01877_, _01876_);
  and (_26904_[12], _01879_, _22762_);
  and (_01880_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_01882_, _23953_, _25842_);
  or (_01883_, _01882_, _01880_);
  and (_26904_[13], _01883_, _22762_);
  and (_01884_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_01886_, _23953_, _25846_);
  or (_01887_, _01886_, _01884_);
  and (_26904_[14], _01887_, _22762_);
  and (_01888_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_01889_, _23953_, _25850_);
  or (_01890_, _01889_, _01888_);
  and (_26904_[15], _01890_, _22762_);
  and (_01891_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_01892_, _23953_, _25854_);
  or (_01893_, _01892_, _01891_);
  and (_26904_[16], _01893_, _22762_);
  and (_01894_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_01895_, _23953_, _25858_);
  or (_01896_, _01895_, _01894_);
  and (_26904_[17], _01896_, _22762_);
  and (_01897_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01898_, _23953_, _25862_);
  or (_01899_, _01898_, _01897_);
  and (_26904_[18], _01899_, _22762_);
  and (_01900_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_01902_, _23953_, _25866_);
  or (_01903_, _01902_, _01900_);
  and (_26904_[19], _01903_, _22762_);
  and (_01904_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_01905_, _23953_, _25870_);
  or (_01906_, _01905_, _01904_);
  and (_26904_[20], _01906_, _22762_);
  and (_01907_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_01908_, _23953_, _25876_);
  or (_01909_, _01908_, _01907_);
  and (_26904_[21], _01909_, _22762_);
  and (_01910_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_01911_, _23953_, _25880_);
  or (_01912_, _01911_, _01910_);
  and (_26904_[22], _01912_, _22762_);
  and (_01913_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_01914_, _23953_, _25884_);
  or (_01915_, _01914_, _01913_);
  and (_26904_[23], _01915_, _22762_);
  and (_01916_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_01917_, _25888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_01918_, _01917_, _01916_);
  and (_26904_[24], _01918_, _22762_);
  and (_01919_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_01920_, _23953_, _25892_);
  or (_01921_, _01920_, _01919_);
  and (_26904_[25], _01921_, _22762_);
  and (_01922_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_01923_, _23953_, _25896_);
  or (_01924_, _01923_, _01922_);
  and (_26904_[26], _01924_, _22762_);
  and (_01925_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_01926_, _23953_, _25900_);
  or (_01927_, _01926_, _01925_);
  and (_26904_[27], _01927_, _22762_);
  and (_01929_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_01930_, _23953_, _25904_);
  or (_01931_, _01930_, _01929_);
  and (_26904_[28], _01931_, _22762_);
  and (_01932_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_01934_, _23953_, _25908_);
  or (_01935_, _01934_, _01932_);
  and (_26904_[29], _01935_, _22762_);
  and (_01936_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_01937_, _23953_, _25912_);
  or (_01938_, _01937_, _01936_);
  and (_26904_[30], _01938_, _22762_);
  and (_01939_, _01759_, _23707_);
  and (_01940_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_22635_, _01940_, _01939_);
  and (_01941_, _25733_, _23946_);
  and (_01942_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_22636_, _01942_, _01941_);
  and (_01944_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_01945_, _25763_, _23898_);
  or (_22637_, _01945_, _01944_);
  and (_01947_, _25733_, _24050_);
  and (_01948_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_22638_, _01948_, _01947_);
  and (_01949_, _25733_, _23747_);
  and (_01950_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_22639_, _01950_, _01949_);
  and (_01951_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_01952_, _25763_, _23778_);
  or (_22640_, _01952_, _01951_);
  not (_01954_, _24096_);
  or (_01955_, _26565_, _01954_);
  or (_01956_, _24096_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_01957_, _01956_, _22762_);
  and (_26908_[0], _01957_, _01955_);
  nand (_01958_, _00372_, _24096_);
  or (_01959_, _24096_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_01960_, _01959_, _22762_);
  and (_26908_[1], _01960_, _01958_);
  or (_01961_, _00451_, _01954_);
  or (_01962_, _24096_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_01963_, _01962_, _22762_);
  and (_26908_[2], _01963_, _01961_);
  or (_01964_, _00545_, _01954_);
  or (_01965_, _24096_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_01966_, _01965_, _22762_);
  and (_26908_[3], _01966_, _01964_);
  and (_01967_, _25078_, _24201_);
  not (_01968_, _01967_);
  and (_01969_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and (_01970_, _01967_, _24050_);
  or (_22641_, _01970_, _01969_);
  and (_01971_, _24329_, _23664_);
  and (_01972_, _01971_, _23778_);
  not (_01973_, _01971_);
  and (_01974_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or (_22642_, _01974_, _01972_);
  and (_01975_, _24063_, _23662_);
  and (_01977_, _01975_, _24297_);
  and (_01978_, _01975_, _24126_);
  nor (_01979_, _01978_, _01977_);
  or (_01980_, _01979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_01981_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_01982_, _01981_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_01983_, _01982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_01984_, _01983_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_01985_, _01984_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_01986_, _01985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_01987_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_01988_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_01989_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_01990_, _01989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_01992_, _01990_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_01993_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_01994_, _01993_, _01992_);
  and (_01995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_01996_, _01995_, _01994_);
  not (_01997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nor (_01998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_01999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_02000_, _01999_, _01998_);
  and (_02001_, _02000_, _01997_);
  not (_02002_, _02001_);
  or (_02004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_02005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_02006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _02005_);
  and (_02007_, _02006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_02009_, _02007_, _02004_);
  and (_02010_, _02009_, _01998_);
  and (_02011_, _02010_, _02002_);
  nand (_02012_, _02011_, _01996_);
  nand (_02014_, _02012_, _01979_);
  and (_02015_, _02014_, _22762_);
  and (_22644_, _02015_, _01980_);
  nand (_02016_, _01978_, _23702_);
  not (_02017_, _01977_);
  and (_02018_, _02009_, _01994_);
  and (_02019_, _02018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_02020_, _02019_, _02001_);
  and (_02021_, _02020_, _02017_);
  or (_02022_, _02021_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_02023_, _02019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_02024_, _02023_, _02002_);
  and (_02025_, _01998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not (_02026_, _02025_);
  and (_02027_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_02028_, _02027_, _01977_);
  or (_02029_, _02028_, _02024_);
  and (_02030_, _02029_, _02022_);
  or (_02031_, _02030_, _01978_);
  and (_02032_, _02031_, _22762_);
  and (_22645_, _02032_, _02016_);
  and (_02034_, _24655_, _24064_);
  or (_02035_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_02036_, _02035_, _22762_);
  not (_02037_, _02034_);
  or (_02038_, _02037_, _23816_);
  and (_22646_, _02038_, _02036_);
  nor (_02039_, _02017_, _23702_);
  and (_02040_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_02041_, _02009_, _01996_);
  and (_02042_, _02041_, _02040_);
  and (_02043_, _02009_, _01986_);
  or (_02044_, _02043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_02045_, _02043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_02046_, _02045_, _02044_);
  or (_02047_, _02046_, _02001_);
  or (_02048_, _02047_, _02042_);
  or (_02049_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_02050_, _02049_, _01979_);
  and (_02051_, _02050_, _02048_);
  and (_02052_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_02053_, _02052_, _02051_);
  or (_02054_, _02053_, _02039_);
  and (_22647_, _02054_, _22762_);
  not (_02055_, _01998_);
  and (_02056_, _02009_, _02055_);
  and (_02057_, _02056_, _01979_);
  or (_02058_, _02057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_02059_, _01996_);
  nand (_02061_, _02057_, _02059_);
  and (_02063_, _02061_, _22762_);
  and (_22648_, _02063_, _02058_);
  nor (_02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_02065_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _22762_);
  and (_02067_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_22649_, _02067_, _02065_);
  and (_02069_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_02070_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_22650_, _02070_, _02069_);
  and (_02071_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_02072_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_22651_, _02072_, _02071_);
  and (_02073_, _01975_, _24119_);
  nand (_02074_, _02073_, _23702_);
  and (_02075_, _02025_, _01999_);
  not (_02076_, _02075_);
  and (_02077_, _01975_, _24292_);
  nor (_02078_, _02077_, _02076_);
  not (_02079_, _02078_);
  and (_02080_, _02079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_02081_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_02082_, _02081_, _02080_);
  or (_02083_, _02082_, _02073_);
  and (_02084_, _02083_, _22762_);
  and (_22652_, _02084_, _02074_);
  and (_22653_, t2ex_i, _22762_);
  nand (_02086_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _22762_);
  nor (_22654_, _02086_, t2_i);
  and (_22655_, t2_i, _22762_);
  and (_02087_, _01758_, _23991_);
  and (_02088_, _02087_, _23707_);
  not (_02089_, _02087_);
  and (_02090_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_22656_, _02090_, _02088_);
  and (_02091_, _24173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_02092_, _24177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or (_02093_, _02092_, _24257_);
  and (_02094_, _02093_, _24255_);
  or (_02095_, _02092_, _24243_);
  and (_02096_, _02095_, _24132_);
  and (_02097_, _25584_, _24145_);
  or (_02099_, _02097_, _02092_);
  and (_02100_, _02099_, _24184_);
  or (_02101_, _02100_, _02096_);
  or (_02102_, _02101_, _02094_);
  or (_02103_, _02102_, _02091_);
  and (_02104_, _02103_, _24128_);
  and (_22657_, _02104_, _24166_);
  and (_02105_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_02106_, _25763_, _23824_);
  or (_22658_, _02106_, _02105_);
  and (_02107_, _24356_, _23069_);
  and (_02108_, _02107_, _23649_);
  not (_02109_, _02107_);
  and (_02110_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or (_22659_, _02110_, _02108_);
  and (_02111_, _23790_, _23707_);
  and (_02112_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or (_22660_, _02112_, _02111_);
  and (_02113_, _01759_, _23778_);
  and (_02114_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_22661_, _02114_, _02113_);
  and (_02115_, _01759_, _23824_);
  and (_02116_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_22662_, _02116_, _02115_);
  and (_22663_, _01787_, _24862_);
  and (_02117_, _24862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_02118_, _02117_, _24951_);
  and (_22664_, _02118_, _22762_);
  or (_02119_, _25057_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_02120_, _02119_, _25056_);
  and (_02121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _24865_);
  nand (_02122_, _02121_, _24904_);
  nand (_02123_, _02122_, _24913_);
  or (_02124_, _02123_, _02120_);
  or (_02125_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_02126_, _02125_, _24913_);
  and (_02127_, _02126_, _24908_);
  and (_02128_, _02127_, _02124_);
  and (_02129_, _02121_, _24907_);
  or (_02130_, _02129_, _02128_);
  and (_02131_, _02130_, _24949_);
  nand (_02132_, _24917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nand (_02133_, _02132_, _25004_);
  or (_02134_, _02133_, _02131_);
  or (_02135_, _24954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_02136_, _02135_, _22762_);
  not (_02137_, _24895_);
  nor (_02138_, _02121_, _02137_);
  nor (_02139_, _02138_, _25136_);
  or (_02140_, _25041_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_02141_, _02140_, _25044_);
  nand (_02142_, _02121_, _24891_);
  nand (_02143_, _02142_, _24888_);
  or (_02144_, _02143_, _02141_);
  or (_02145_, _02125_, _24888_);
  and (_02146_, _02145_, _24883_);
  and (_02147_, _02146_, _02144_);
  or (_02148_, _02147_, _24862_);
  or (_02149_, _02148_, _02139_);
  and (_02150_, _02149_, _02136_);
  and (_22665_, _02150_, _02134_);
  or (_02151_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _24865_);
  or (_02152_, _02151_, _24913_);
  and (_02153_, _02152_, _24908_);
  or (_02154_, _24980_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_02155_, _02154_, _24979_);
  and (_02156_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_02157_, _02156_, _24904_);
  nand (_02158_, _02157_, _24913_);
  or (_02159_, _02158_, _02155_);
  and (_02160_, _02159_, _02153_);
  and (_02161_, _02156_, _24907_);
  or (_02162_, _02161_, _02160_);
  and (_02163_, _02162_, _24949_);
  nand (_02164_, _24917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nand (_02165_, _02164_, _25004_);
  or (_02166_, _02165_, _02163_);
  or (_02167_, _24954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_02168_, _02167_, _22762_);
  nor (_02169_, _02156_, _02137_);
  nor (_02170_, _02169_, _25136_);
  or (_02171_, _24958_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_02172_, _02171_, _24956_);
  nand (_02173_, _02156_, _24891_);
  nand (_02174_, _02173_, _24888_);
  or (_02175_, _02174_, _02172_);
  or (_02176_, _02151_, _24888_);
  and (_02177_, _02176_, _24883_);
  and (_02178_, _02177_, _02175_);
  or (_02179_, _02178_, _24862_);
  or (_02180_, _02179_, _02170_);
  and (_02181_, _02180_, _02168_);
  and (_22666_, _02181_, _02166_);
  and (_02182_, _24730_, _24125_);
  nand (_02183_, _02182_, _23594_);
  or (_02184_, _02182_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_02185_, _02184_, _24737_);
  and (_02186_, _02185_, _02183_);
  and (_02187_, _24736_, _23939_);
  or (_02188_, _02187_, _02186_);
  and (_22667_, _02188_, _22762_);
  and (_02189_, _24648_, _24296_);
  nand (_02190_, _02189_, _23594_);
  or (_02191_, _02189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_02192_, _02191_, _24659_);
  and (_02193_, _02192_, _02190_);
  and (_02194_, _24658_, _23642_);
  or (_02195_, _02194_, _02193_);
  and (_22668_, _02195_, _22762_);
  and (_02196_, _01759_, _23898_);
  and (_02197_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_22669_, _02197_, _02196_);
  and (_02198_, _23707_, _23077_);
  and (_02199_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or (_22670_, _02199_, _02198_);
  and (_02200_, _24356_, _23986_);
  and (_02201_, _02200_, _23898_);
  not (_02202_, _02200_);
  and (_02203_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_22671_, _02203_, _02201_);
  and (_02204_, _24766_, _23986_);
  not (_02205_, _02204_);
  and (_02206_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_02207_, _02204_, _23747_);
  or (_22672_, _02207_, _02206_);
  and (_02208_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_02209_, _02204_, _23649_);
  or (_27039_, _02209_, _02208_);
  and (_02211_, _02087_, _23778_);
  and (_02212_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_27008_, _02212_, _02211_);
  and (_02213_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_02214_, _02204_, _23824_);
  or (_27038_, _02214_, _02213_);
  and (_02215_, _01758_, _23903_);
  and (_02216_, _02215_, _23707_);
  not (_02217_, _02215_);
  and (_02218_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_22673_, _02218_, _02216_);
  nor (_26897_[2], _00470_, rst);
  nor (_26887_[5], _00006_, rst);
  and (_02219_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_02220_, _02204_, _24050_);
  or (_22674_, _02220_, _02219_);
  and (_02221_, _02087_, _23898_);
  and (_02222_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_22675_, _02222_, _02221_);
  and (_02223_, _02087_, _23747_);
  and (_02224_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_22676_, _02224_, _02223_);
  and (_02225_, _02087_, _23824_);
  and (_02226_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_22677_, _02226_, _02225_);
  and (_02227_, _24331_, _23707_);
  and (_02228_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_22678_, _02228_, _02227_);
  and (_02229_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_02230_, _02204_, _23946_);
  or (_27040_, _02230_, _02229_);
  nor (_26860_[0], _24402_, rst);
  nor (_26860_[6], _24486_, rst);
  and (_02231_, _24852_, _23707_);
  and (_02232_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or (_22679_, _02232_, _02231_);
  and (_02233_, _24006_, _23946_);
  and (_02234_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or (_22680_, _02234_, _02233_);
  and (_02235_, _02215_, _23778_);
  and (_02236_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_22681_, _02236_, _02235_);
  and (_02237_, _02215_, _23824_);
  and (_02238_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_22682_, _02238_, _02237_);
  and (_02239_, _02215_, _23898_);
  and (_02240_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_22683_, _02240_, _02239_);
  and (_02241_, _24275_, _23789_);
  and (_02242_, _02241_, _23747_);
  not (_02243_, _02241_);
  and (_02244_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_27293_, _02244_, _02242_);
  and (_02245_, _24766_, _23069_);
  not (_02246_, _02245_);
  and (_02247_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  and (_02248_, _02245_, _23707_);
  or (_27037_, _02248_, _02247_);
  and (_02249_, _24050_, _23077_);
  and (_02250_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or (_22684_, _02250_, _02249_);
  and (_02251_, _23946_, _23077_);
  and (_02252_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or (_22685_, _02252_, _02251_);
  and (_02253_, _25618_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_02254_, _24596_, _24539_);
  or (_02255_, _02254_, _24585_);
  and (_02256_, _24556_, _24546_);
  or (_02257_, _02256_, _25640_);
  and (_02258_, _24613_, _26650_);
  or (_02259_, _02258_, _26666_);
  and (_02260_, _24613_, _24604_);
  and (_02261_, _26625_, _24582_);
  and (_02262_, _26625_, _24540_);
  or (_02263_, _02262_, _02261_);
  or (_02264_, _02263_, _02260_);
  or (_02265_, _02264_, _26591_);
  or (_02266_, _02265_, _02259_);
  and (_02267_, _26650_, _26582_);
  and (_02268_, _24567_, _24546_);
  or (_02269_, _02268_, _02267_);
  and (_02270_, _24604_, _24556_);
  and (_02271_, _24593_, _24556_);
  or (_02272_, _02271_, _02270_);
  and (_02273_, _24606_, _24556_);
  and (_02274_, _24589_, _24556_);
  or (_02275_, _02274_, _02273_);
  or (_02276_, _02275_, _02272_);
  or (_02277_, _02276_, _02269_);
  or (_02278_, _02277_, _02266_);
  or (_02279_, _02278_, _02257_);
  or (_02280_, _02279_, _02255_);
  and (_02281_, _02280_, _25644_);
  or (_26867_[0], _02281_, _02253_);
  and (_02282_, _24283_, _23898_);
  and (_02283_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or (_22686_, _02283_, _02282_);
  and (_02284_, _01809_, _24329_);
  and (_02285_, _02284_, _24050_);
  not (_02286_, _02284_);
  and (_02287_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  or (_22687_, _02287_, _02285_);
  and (_02288_, _02284_, _23649_);
  and (_02289_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  or (_22688_, _02289_, _02288_);
  and (_02290_, _02284_, _23747_);
  and (_02291_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or (_22689_, _02291_, _02290_);
  and (_02292_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and (_02293_, _24692_, _24050_);
  or (_22690_, _02293_, _02292_);
  and (_02294_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and (_02295_, _24692_, _23707_);
  or (_27236_, _02295_, _02294_);
  and (_02296_, _02284_, _23778_);
  and (_02297_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  or (_27115_, _02297_, _02296_);
  and (_02298_, _24201_, _23752_);
  not (_02299_, _02298_);
  and (_02300_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  and (_02301_, _02298_, _23778_);
  or (_22691_, _02301_, _02300_);
  and (_02302_, _01809_, _23752_);
  and (_02303_, _02302_, _23707_);
  not (_02304_, _02302_);
  and (_02305_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_22692_, _02305_, _02303_);
  and (_02306_, _24201_, _23069_);
  not (_02307_, _02306_);
  and (_02308_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  and (_02309_, _02306_, _23824_);
  or (_22693_, _02309_, _02308_);
  and (_02310_, _24678_, _23003_);
  and (_02311_, _25769_, _23073_);
  and (_02312_, _02311_, _02310_);
  and (_02313_, _02312_, _25926_);
  and (_02314_, _02313_, _24043_);
  not (_02315_, _02313_);
  and (_02316_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_22694_, _02316_, _02314_);
  and (_02317_, _02302_, _23946_);
  and (_02318_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_22695_, _02318_, _02317_);
  and (_02319_, _02302_, _23747_);
  and (_02320_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_22696_, _02320_, _02319_);
  and (_02321_, _24356_, _23752_);
  and (_02322_, _02321_, _23649_);
  not (_02323_, _02321_);
  and (_02324_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  or (_22697_, _02324_, _02322_);
  and (_02325_, _23662_, _23072_);
  and (_02326_, _02325_, _24329_);
  and (_02327_, _02326_, _23778_);
  not (_02328_, _02326_);
  and (_02329_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_22698_, _02329_, _02327_);
  and (_02330_, _02302_, _23898_);
  and (_02331_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_22699_, _02331_, _02330_);
  and (_02332_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and (_02333_, _24692_, _23649_);
  or (_27235_, _02333_, _02332_);
  and (_02334_, _02215_, _23946_);
  and (_02335_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_26992_, _02335_, _02334_);
  and (_02336_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_02337_, _02204_, _23778_);
  or (_22700_, _02337_, _02336_);
  and (_02339_, _02215_, _23649_);
  and (_02340_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_22701_, _02340_, _02339_);
  nor (_26887_[0], _00129_, rst);
  and (_02341_, _25748_, _23824_);
  and (_02342_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_22702_, _02342_, _02341_);
  and (_02343_, _02215_, _23747_);
  and (_02344_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_22703_, _02344_, _02343_);
  and (_02345_, _01808_, _24370_);
  and (_02346_, _02345_, _23778_);
  not (_02347_, _02345_);
  and (_02349_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_22704_, _02349_, _02346_);
  and (_02350_, _01758_, _24005_);
  and (_02351_, _02350_, _23649_);
  not (_02352_, _02350_);
  and (_02353_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_22705_, _02353_, _02351_);
  nor (_02354_, _23596_, _26379_);
  and (_02355_, _26385_, _23596_);
  or (_02356_, _02355_, _02354_);
  and (_22706_, _02356_, _22762_);
  and (_02357_, _02200_, _23649_);
  and (_02358_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_27166_, _02358_, _02357_);
  and (_02359_, _02325_, _01808_);
  and (_02360_, _02359_, _24050_);
  not (_02361_, _02359_);
  and (_02363_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  or (_27155_, _02363_, _02360_);
  and (_02364_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and (_02365_, _24692_, _23946_);
  or (_22707_, _02365_, _02364_);
  and (_02366_, _01971_, _23898_);
  and (_02367_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  or (_22708_, _02367_, _02366_);
  and (_02368_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and (_02369_, _24692_, _23747_);
  or (_22709_, _02369_, _02368_);
  and (_02370_, _24005_, _23754_);
  and (_02371_, _02370_, _23898_);
  not (_02372_, _02370_);
  and (_02373_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_22710_, _02373_, _02371_);
  and (_02374_, _01809_, _23656_);
  and (_02375_, _02374_, _24050_);
  not (_02376_, _02374_);
  and (_02377_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  or (_22711_, _02377_, _02375_);
  nor (_02378_, _26656_, _26668_);
  nand (_02379_, _02378_, _26597_);
  or (_02380_, _26644_, _26652_);
  or (_02381_, _26660_, _26641_);
  or (_02382_, _02381_, _26637_);
  or (_02383_, _02382_, _02380_);
  or (_02384_, _02383_, _02379_);
  and (_02385_, _02384_, _26572_);
  and (_02386_, _25629_, _24566_);
  nor (_02387_, _02386_, _02385_);
  not (_02388_, _02387_);
  nor (_02389_, _02388_, _00099_);
  not (_02390_, _02389_);
  or (_02391_, _02387_, _26777_);
  or (_02392_, _02391_, _00058_);
  and (_02393_, _02392_, _02390_);
  and (_02394_, _02393_, _22985_);
  nor (_02395_, _02393_, _22985_);
  or (_02396_, _02395_, _02394_);
  not (_02397_, _00058_);
  and (_02398_, _02391_, _02397_);
  nor (_02399_, _02398_, _23904_);
  and (_02400_, _02391_, _00014_);
  nor (_02401_, _02400_, _23658_);
  nor (_02402_, _02401_, _02399_);
  not (_02403_, _23786_);
  not (_02404_, _26817_);
  and (_02405_, _02391_, _02404_);
  nor (_02406_, _02405_, _02403_);
  and (_02407_, _02405_, _02403_);
  nor (_02408_, _02407_, _02406_);
  and (_02409_, _02408_, _02402_);
  and (_02410_, _02409_, _02396_);
  not (_02411_, _02391_);
  and (_02412_, _02411_, _26817_);
  and (_02413_, _02391_, _00037_);
  nor (_02414_, _02413_, _02412_);
  and (_02415_, _02414_, _23039_);
  nor (_02416_, _02414_, _23039_);
  or (_02417_, _02416_, _02415_);
  not (_02418_, _23067_);
  nor (_02419_, _02388_, _00168_);
  nor (_02420_, _02391_, _00014_);
  nor (_02421_, _02420_, _02419_);
  nor (_02422_, _02421_, _02418_);
  and (_02423_, _02421_, _02418_);
  nor (_02424_, _02423_, _02422_);
  not (_02425_, _02424_);
  nor (_02426_, _02425_, _02417_);
  or (_02427_, _02388_, _00134_);
  or (_02428_, _02391_, _00037_);
  nand (_02429_, _02428_, _02427_);
  and (_02430_, _02429_, _23020_);
  nor (_02431_, _02429_, _23020_);
  nor (_02432_, _02431_, _02430_);
  and (_02433_, _02400_, _23658_);
  not (_02434_, _02433_);
  and (_02435_, _02398_, _23904_);
  not (_02436_, _02435_);
  nor (_02438_, _26781_, _22947_);
  and (_02439_, _02438_, _02436_);
  and (_02440_, _02439_, _02434_);
  and (_02441_, _02440_, _02432_);
  and (_02442_, _02441_, _02426_);
  and (_02443_, _02442_, _02410_);
  not (_02444_, _26777_);
  not (_02445_, _02393_);
  and (_02447_, _02428_, _02427_);
  and (_02448_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_02449_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_02450_, _02449_, _02448_);
  and (_02451_, _02450_, _02445_);
  and (_02452_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_02453_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_02454_, _02453_, _02452_);
  and (_02455_, _02454_, _02393_);
  or (_02456_, _02455_, _02451_);
  or (_02457_, _02456_, _02421_);
  not (_02458_, _02414_);
  not (_02459_, _02421_);
  and (_02460_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_02461_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_02462_, _02461_, _02460_);
  and (_02463_, _02462_, _02445_);
  and (_02464_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_02465_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_02466_, _02465_, _02464_);
  and (_02467_, _02466_, _02393_);
  or (_02468_, _02467_, _02463_);
  or (_02469_, _02468_, _02459_);
  and (_02470_, _02469_, _02458_);
  and (_02471_, _02470_, _02457_);
  or (_02472_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_02473_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_02474_, _02473_, _02393_);
  and (_02475_, _02474_, _02472_);
  or (_02476_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_02477_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_02478_, _02477_, _02445_);
  and (_02479_, _02478_, _02476_);
  or (_02480_, _02479_, _02475_);
  or (_02481_, _02480_, _02459_);
  or (_02482_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_02483_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_02484_, _02483_, _02393_);
  and (_02485_, _02484_, _02482_);
  or (_02486_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_02487_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_02488_, _02487_, _02445_);
  and (_02489_, _02488_, _02486_);
  or (_02490_, _02489_, _02485_);
  or (_02491_, _02490_, _02421_);
  and (_02492_, _02491_, _02414_);
  and (_02493_, _02492_, _02481_);
  or (_02494_, _02493_, _02471_);
  or (_02495_, _02494_, _02398_);
  not (_02496_, _02398_);
  and (_02497_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and (_02498_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_02499_, _02498_, _02393_);
  or (_02500_, _02499_, _02497_);
  and (_02501_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and (_02502_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_02503_, _02502_, _02445_);
  or (_02504_, _02503_, _02501_);
  and (_02505_, _02504_, _02500_);
  or (_02506_, _02505_, _02459_);
  and (_02507_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and (_02508_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_02509_, _02508_, _02393_);
  or (_02510_, _02509_, _02507_);
  and (_02511_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and (_02512_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_02513_, _02512_, _02445_);
  or (_02514_, _02513_, _02511_);
  and (_02515_, _02514_, _02510_);
  or (_02516_, _02515_, _02421_);
  and (_02517_, _02516_, _02458_);
  and (_02518_, _02517_, _02506_);
  or (_02519_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_02520_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and (_02521_, _02520_, _02519_);
  or (_02522_, _02521_, _02445_);
  or (_02523_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_02524_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and (_02525_, _02524_, _02523_);
  or (_02526_, _02525_, _02393_);
  and (_02527_, _02526_, _02522_);
  or (_02528_, _02527_, _02459_);
  or (_02529_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_02530_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and (_02531_, _02530_, _02529_);
  or (_02532_, _02531_, _02445_);
  or (_02533_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_02534_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and (_02535_, _02534_, _02533_);
  or (_02536_, _02535_, _02393_);
  and (_02537_, _02536_, _02532_);
  or (_02538_, _02537_, _02421_);
  and (_02540_, _02538_, _02414_);
  and (_02541_, _02540_, _02528_);
  or (_02542_, _02541_, _02518_);
  or (_02543_, _02542_, _02496_);
  and (_02544_, _02543_, _02400_);
  and (_02545_, _02544_, _02495_);
  not (_02546_, _02400_);
  and (_02547_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and (_02548_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_02549_, _02548_, _02547_);
  and (_02550_, _02549_, _02393_);
  and (_02551_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and (_02552_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_02553_, _02552_, _02551_);
  and (_02554_, _02553_, _02445_);
  or (_02556_, _02554_, _02550_);
  or (_02557_, _02556_, _02459_);
  and (_02558_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and (_02559_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_02560_, _02559_, _02558_);
  and (_02561_, _02560_, _02393_);
  and (_02562_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and (_02563_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_02564_, _02563_, _02562_);
  and (_02565_, _02564_, _02445_);
  or (_02566_, _02565_, _02561_);
  or (_02567_, _02566_, _02421_);
  and (_02568_, _02567_, _02458_);
  and (_02569_, _02568_, _02557_);
  or (_02570_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_02572_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and (_02573_, _02572_, _02445_);
  and (_02574_, _02573_, _02570_);
  or (_02575_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_02576_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and (_02577_, _02576_, _02393_);
  and (_02578_, _02577_, _02575_);
  or (_02579_, _02578_, _02574_);
  or (_02580_, _02579_, _02459_);
  or (_02581_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_02583_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and (_02584_, _02583_, _02445_);
  and (_02585_, _02584_, _02581_);
  or (_02586_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_02587_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and (_02588_, _02587_, _02393_);
  and (_02589_, _02588_, _02586_);
  or (_02590_, _02589_, _02585_);
  or (_02591_, _02590_, _02421_);
  and (_02592_, _02591_, _02414_);
  and (_02593_, _02592_, _02580_);
  or (_02594_, _02593_, _02569_);
  and (_02595_, _02594_, _02496_);
  and (_02596_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_02597_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_02598_, _02597_, _02596_);
  and (_02599_, _02598_, _02393_);
  and (_02600_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and (_02601_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_02602_, _02601_, _02600_);
  and (_02603_, _02602_, _02445_);
  or (_02604_, _02603_, _02599_);
  or (_02605_, _02604_, _02459_);
  and (_02606_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and (_02607_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_02608_, _02607_, _02606_);
  and (_02609_, _02608_, _02393_);
  and (_02610_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and (_02611_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_02612_, _02611_, _02610_);
  and (_02613_, _02612_, _02445_);
  or (_02614_, _02613_, _02609_);
  or (_02615_, _02614_, _02421_);
  and (_02616_, _02615_, _02458_);
  and (_02617_, _02616_, _02605_);
  or (_02618_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_02619_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and (_02620_, _02619_, _02618_);
  and (_02621_, _02620_, _02393_);
  or (_02622_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_02623_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and (_02624_, _02623_, _02622_);
  and (_02625_, _02624_, _02445_);
  or (_02626_, _02625_, _02621_);
  or (_02627_, _02626_, _02459_);
  or (_02628_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_02629_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and (_02630_, _02629_, _02628_);
  and (_02631_, _02630_, _02393_);
  or (_02632_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_02633_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and (_02634_, _02633_, _02632_);
  and (_02635_, _02634_, _02445_);
  or (_02636_, _02635_, _02631_);
  or (_02637_, _02636_, _02421_);
  and (_02638_, _02637_, _02414_);
  and (_02639_, _02638_, _02627_);
  or (_02640_, _02639_, _02617_);
  and (_02641_, _02640_, _02398_);
  or (_02642_, _02641_, _02595_);
  and (_02643_, _02642_, _02546_);
  or (_02644_, _02643_, _02545_);
  or (_02645_, _02644_, _02405_);
  not (_02646_, _02405_);
  and (_02647_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  and (_02648_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or (_02649_, _02648_, _02647_);
  and (_02650_, _02649_, _02393_);
  and (_02651_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and (_02652_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or (_02653_, _02652_, _02651_);
  and (_02654_, _02653_, _02445_);
  or (_02655_, _02654_, _02650_);
  and (_02656_, _02655_, _02421_);
  and (_02657_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  and (_02658_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or (_02659_, _02658_, _02657_);
  and (_02660_, _02659_, _02393_);
  and (_02661_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and (_02662_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or (_02664_, _02662_, _02661_);
  and (_02665_, _02664_, _02445_);
  or (_02666_, _02665_, _02660_);
  and (_02667_, _02666_, _02459_);
  or (_02668_, _02667_, _02414_);
  or (_02669_, _02668_, _02656_);
  or (_02670_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or (_02671_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and (_02672_, _02671_, _02670_);
  and (_02673_, _02672_, _02393_);
  or (_02674_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or (_02675_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  and (_02676_, _02675_, _02674_);
  and (_02677_, _02676_, _02445_);
  or (_02678_, _02677_, _02673_);
  and (_02679_, _02678_, _02421_);
  or (_02680_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or (_02681_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  and (_02682_, _02681_, _02680_);
  and (_02683_, _02682_, _02393_);
  or (_02684_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or (_02685_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and (_02686_, _02685_, _02684_);
  and (_02687_, _02686_, _02445_);
  or (_02688_, _02687_, _02683_);
  and (_02689_, _02688_, _02459_);
  or (_02690_, _02689_, _02458_);
  or (_02691_, _02690_, _02679_);
  and (_02692_, _02691_, _02669_);
  or (_02693_, _02692_, _02398_);
  and (_02694_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and (_02695_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_02696_, _02695_, _02694_);
  and (_02697_, _02696_, _02393_);
  and (_02698_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and (_02699_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_02700_, _02699_, _02698_);
  and (_02701_, _02700_, _02445_);
  or (_02702_, _02701_, _02697_);
  and (_02703_, _02702_, _02421_);
  and (_02704_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and (_02705_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_02706_, _02705_, _02704_);
  and (_02707_, _02706_, _02393_);
  and (_02708_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and (_02709_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_02710_, _02709_, _02708_);
  and (_02711_, _02710_, _02445_);
  or (_02712_, _02711_, _02707_);
  and (_02713_, _02712_, _02459_);
  or (_02715_, _02713_, _02414_);
  or (_02716_, _02715_, _02703_);
  or (_02717_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_02718_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and (_02719_, _02718_, _02717_);
  and (_02720_, _02719_, _02393_);
  or (_02721_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_02722_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and (_02723_, _02722_, _02721_);
  and (_02724_, _02723_, _02445_);
  or (_02725_, _02724_, _02720_);
  and (_02726_, _02725_, _02421_);
  or (_02727_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_02728_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and (_02729_, _02728_, _02727_);
  and (_02730_, _02729_, _02393_);
  or (_02731_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_02732_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and (_02733_, _02732_, _02731_);
  and (_02734_, _02733_, _02445_);
  or (_02735_, _02734_, _02730_);
  and (_02736_, _02735_, _02459_);
  or (_02737_, _02736_, _02458_);
  or (_02738_, _02737_, _02726_);
  and (_02739_, _02738_, _02716_);
  or (_02740_, _02739_, _02496_);
  and (_02741_, _02740_, _02400_);
  and (_02742_, _02741_, _02693_);
  and (_02743_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and (_02744_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_02745_, _02744_, _02743_);
  and (_02746_, _02745_, _02445_);
  and (_02747_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and (_02748_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_02749_, _02748_, _02747_);
  and (_02750_, _02749_, _02393_);
  or (_02751_, _02750_, _02746_);
  or (_02752_, _02751_, _02459_);
  and (_02753_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and (_02754_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_02755_, _02754_, _02753_);
  and (_02756_, _02755_, _02445_);
  and (_02757_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and (_02758_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_02759_, _02758_, _02757_);
  and (_02760_, _02759_, _02393_);
  or (_02761_, _02760_, _02756_);
  or (_02762_, _02761_, _02421_);
  and (_02763_, _02762_, _02458_);
  and (_02764_, _02763_, _02752_);
  or (_02765_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_02766_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and (_02767_, _02766_, _02393_);
  and (_02768_, _02767_, _02765_);
  or (_02769_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_02770_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and (_02771_, _02770_, _02445_);
  and (_02772_, _02771_, _02769_);
  or (_02773_, _02772_, _02768_);
  or (_02774_, _02773_, _02459_);
  or (_02775_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_02776_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and (_02777_, _02776_, _02393_);
  and (_02778_, _02777_, _02775_);
  or (_02779_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_02780_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and (_02781_, _02780_, _02445_);
  and (_02782_, _02781_, _02779_);
  or (_02783_, _02782_, _02778_);
  or (_02784_, _02783_, _02421_);
  and (_02785_, _02784_, _02414_);
  and (_02786_, _02785_, _02774_);
  or (_02787_, _02786_, _02764_);
  and (_02788_, _02787_, _02496_);
  and (_02789_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and (_02790_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_02791_, _02790_, _02393_);
  or (_02792_, _02791_, _02789_);
  and (_02793_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and (_02794_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_02795_, _02794_, _02445_);
  or (_02796_, _02795_, _02793_);
  and (_02797_, _02796_, _02792_);
  or (_02798_, _02797_, _02459_);
  and (_02799_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and (_02800_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_02801_, _02800_, _02393_);
  or (_02802_, _02801_, _02799_);
  and (_02803_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and (_02804_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_02805_, _02804_, _02445_);
  or (_02806_, _02805_, _02803_);
  and (_02807_, _02806_, _02802_);
  or (_02808_, _02807_, _02421_);
  and (_02809_, _02808_, _02458_);
  and (_02810_, _02809_, _02798_);
  or (_02811_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_02812_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and (_02813_, _02812_, _02811_);
  or (_02814_, _02813_, _02445_);
  or (_02815_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_02816_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and (_02817_, _02816_, _02815_);
  or (_02818_, _02817_, _02393_);
  and (_02819_, _02818_, _02814_);
  or (_02820_, _02819_, _02459_);
  or (_02821_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_02822_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and (_02823_, _02822_, _02821_);
  or (_02824_, _02823_, _02445_);
  or (_02825_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_02827_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and (_02828_, _02827_, _02825_);
  or (_02829_, _02828_, _02393_);
  and (_02830_, _02829_, _02824_);
  or (_02831_, _02830_, _02421_);
  and (_02832_, _02831_, _02414_);
  and (_02833_, _02832_, _02820_);
  or (_02834_, _02833_, _02810_);
  and (_02835_, _02834_, _02398_);
  or (_02836_, _02835_, _02788_);
  and (_02837_, _02836_, _02546_);
  or (_02838_, _02837_, _02742_);
  or (_02839_, _02838_, _02646_);
  and (_02840_, _02839_, _02645_);
  and (_02841_, _02840_, _02444_);
  and (_02842_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and (_02843_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_02845_, _02843_, _02842_);
  and (_02846_, _02845_, _02393_);
  and (_02847_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and (_02848_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_02849_, _02848_, _02847_);
  and (_02850_, _02849_, _02445_);
  or (_02851_, _02850_, _02846_);
  or (_02852_, _02851_, _02459_);
  and (_02853_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and (_02854_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_02855_, _02854_, _02853_);
  and (_02856_, _02855_, _02393_);
  and (_02857_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and (_02858_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_02859_, _02858_, _02857_);
  and (_02860_, _02859_, _02445_);
  or (_02861_, _02860_, _02856_);
  or (_02862_, _02861_, _02421_);
  and (_02863_, _02862_, _02458_);
  and (_02864_, _02863_, _02852_);
  or (_02865_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_02866_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and (_02868_, _02866_, _02865_);
  and (_02869_, _02868_, _02393_);
  or (_02870_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_02871_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and (_02872_, _02871_, _02870_);
  and (_02873_, _02872_, _02445_);
  or (_02875_, _02873_, _02869_);
  or (_02877_, _02875_, _02459_);
  or (_02878_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_02879_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and (_02881_, _02879_, _02878_);
  and (_02883_, _02881_, _02393_);
  or (_02884_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_02885_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and (_02886_, _02885_, _02884_);
  and (_02887_, _02886_, _02445_);
  or (_02888_, _02887_, _02883_);
  or (_02889_, _02888_, _02421_);
  and (_02890_, _02889_, _02414_);
  and (_02891_, _02890_, _02877_);
  or (_02892_, _02891_, _02864_);
  and (_02894_, _02892_, _02398_);
  and (_02895_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_02896_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or (_02897_, _02896_, _02895_);
  and (_02898_, _02897_, _02393_);
  and (_02899_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_02900_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or (_02901_, _02900_, _02899_);
  and (_02902_, _02901_, _02445_);
  or (_02904_, _02902_, _02898_);
  or (_02905_, _02904_, _02459_);
  and (_02907_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_02909_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or (_02910_, _02909_, _02907_);
  and (_02912_, _02910_, _02393_);
  and (_02913_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_02914_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or (_02915_, _02914_, _02913_);
  and (_02916_, _02915_, _02445_);
  or (_02917_, _02916_, _02912_);
  or (_02918_, _02917_, _02421_);
  and (_02919_, _02918_, _02458_);
  and (_02920_, _02919_, _02905_);
  or (_02921_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or (_02922_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_02924_, _02922_, _02445_);
  and (_02925_, _02924_, _02921_);
  or (_02926_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or (_02927_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_02928_, _02927_, _02393_);
  and (_02929_, _02928_, _02926_);
  or (_02930_, _02929_, _02925_);
  or (_02931_, _02930_, _02459_);
  or (_02932_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or (_02933_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_02934_, _02933_, _02445_);
  and (_02935_, _02934_, _02932_);
  or (_02936_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or (_02937_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_02938_, _02937_, _02393_);
  and (_02939_, _02938_, _02936_);
  or (_02940_, _02939_, _02935_);
  or (_02941_, _02940_, _02421_);
  and (_02942_, _02941_, _02414_);
  and (_02943_, _02942_, _02931_);
  or (_02944_, _02943_, _02920_);
  and (_02945_, _02944_, _02496_);
  or (_02946_, _02945_, _02894_);
  and (_02947_, _02946_, _02546_);
  and (_02948_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and (_02949_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or (_02950_, _02949_, _02948_);
  and (_02951_, _02950_, _02393_);
  and (_02952_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and (_02953_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or (_02954_, _02953_, _02952_);
  and (_02955_, _02954_, _02445_);
  or (_02956_, _02955_, _02951_);
  and (_02957_, _02956_, _02421_);
  and (_02958_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and (_02959_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or (_02960_, _02959_, _02958_);
  and (_02961_, _02960_, _02393_);
  and (_02962_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and (_02963_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or (_02964_, _02963_, _02962_);
  and (_02965_, _02964_, _02445_);
  or (_02966_, _02965_, _02961_);
  and (_02967_, _02966_, _02459_);
  or (_02968_, _02967_, _02957_);
  and (_02969_, _02968_, _02458_);
  or (_02970_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or (_02971_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and (_02973_, _02971_, _02445_);
  and (_02974_, _02973_, _02970_);
  or (_02975_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or (_02976_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and (_02977_, _02976_, _02393_);
  and (_02978_, _02977_, _02975_);
  or (_02979_, _02978_, _02974_);
  and (_02980_, _02979_, _02421_);
  or (_02981_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or (_02982_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and (_02983_, _02982_, _02445_);
  and (_02984_, _02983_, _02981_);
  or (_02985_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or (_02986_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and (_02987_, _02986_, _02393_);
  and (_02988_, _02987_, _02985_);
  or (_02989_, _02988_, _02984_);
  and (_02990_, _02989_, _02459_);
  or (_02991_, _02990_, _02980_);
  and (_02992_, _02991_, _02414_);
  or (_02993_, _02992_, _02969_);
  and (_02994_, _02993_, _02496_);
  and (_02995_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_02997_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_02998_, _02997_, _02995_);
  and (_02999_, _02998_, _02393_);
  and (_03000_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_03001_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or (_03002_, _03001_, _03000_);
  and (_03003_, _03002_, _02445_);
  or (_03004_, _03003_, _02999_);
  and (_03005_, _03004_, _02421_);
  and (_03006_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_03007_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_03008_, _03007_, _03006_);
  and (_03009_, _03008_, _02393_);
  and (_03010_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and (_03011_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or (_03012_, _03011_, _03010_);
  and (_03013_, _03012_, _02445_);
  or (_03014_, _03013_, _03009_);
  and (_03015_, _03014_, _02459_);
  or (_03016_, _03015_, _03005_);
  and (_03017_, _03016_, _02458_);
  or (_03018_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or (_03019_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_03020_, _03019_, _03018_);
  and (_03021_, _03020_, _02393_);
  or (_03022_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_03023_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_03024_, _03023_, _03022_);
  and (_03025_, _03024_, _02445_);
  or (_03026_, _03025_, _03021_);
  and (_03027_, _03026_, _02421_);
  or (_03028_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or (_03029_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_03030_, _03029_, _03028_);
  and (_03031_, _03030_, _02393_);
  or (_03032_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_03033_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and (_03034_, _03033_, _03032_);
  and (_03035_, _03034_, _02445_);
  or (_03036_, _03035_, _03031_);
  and (_03037_, _03036_, _02459_);
  or (_03038_, _03037_, _03027_);
  and (_03039_, _03038_, _02414_);
  or (_03040_, _03039_, _03017_);
  and (_03041_, _03040_, _02398_);
  or (_03042_, _03041_, _02994_);
  and (_03043_, _03042_, _02400_);
  or (_03044_, _03043_, _02947_);
  or (_03045_, _03044_, _02405_);
  and (_03047_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and (_03048_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_03049_, _03048_, _03047_);
  and (_03050_, _03049_, _02393_);
  and (_03051_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and (_03053_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_03054_, _03053_, _03051_);
  and (_03055_, _03054_, _02445_);
  or (_03056_, _03055_, _03050_);
  or (_03057_, _03056_, _02459_);
  and (_03058_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and (_03059_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_03060_, _03059_, _03058_);
  and (_03061_, _03060_, _02393_);
  and (_03062_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and (_03063_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_03064_, _03063_, _03062_);
  and (_03065_, _03064_, _02445_);
  or (_03066_, _03065_, _03061_);
  or (_03067_, _03066_, _02421_);
  and (_03068_, _03067_, _02458_);
  and (_03070_, _03068_, _03057_);
  or (_03071_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_03072_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and (_03073_, _03072_, _02445_);
  and (_03074_, _03073_, _03071_);
  or (_03075_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_03076_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and (_03077_, _03076_, _02393_);
  and (_03078_, _03077_, _03075_);
  or (_03079_, _03078_, _03074_);
  or (_03080_, _03079_, _02459_);
  or (_03081_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_03082_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and (_03084_, _03082_, _02445_);
  and (_03085_, _03084_, _03081_);
  or (_03086_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_03087_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and (_03088_, _03087_, _02393_);
  and (_03089_, _03088_, _03086_);
  or (_03090_, _03089_, _03085_);
  or (_03091_, _03090_, _02421_);
  and (_03092_, _03091_, _02414_);
  and (_03093_, _03092_, _03080_);
  or (_03094_, _03093_, _03070_);
  and (_03095_, _03094_, _02496_);
  and (_03096_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and (_03097_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_03098_, _03097_, _03096_);
  and (_03099_, _03098_, _02393_);
  and (_03100_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and (_03101_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_03102_, _03101_, _03100_);
  and (_03103_, _03102_, _02445_);
  or (_03104_, _03103_, _03099_);
  or (_03105_, _03104_, _02459_);
  and (_03106_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and (_03107_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_03109_, _03107_, _03106_);
  and (_03110_, _03109_, _02393_);
  and (_03111_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and (_03112_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_03113_, _03112_, _03111_);
  and (_03115_, _03113_, _02445_);
  or (_03116_, _03115_, _03110_);
  or (_03118_, _03116_, _02421_);
  and (_03119_, _03118_, _02458_);
  and (_03120_, _03119_, _03105_);
  or (_03121_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_03122_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_03124_, _03122_, _03121_);
  and (_03126_, _03124_, _02393_);
  or (_03127_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_03128_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and (_03130_, _03128_, _03127_);
  and (_03131_, _03130_, _02445_);
  or (_03132_, _03131_, _03126_);
  or (_03133_, _03132_, _02459_);
  or (_03134_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_03135_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and (_03136_, _03135_, _03134_);
  and (_03137_, _03136_, _02393_);
  or (_03138_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_03140_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and (_03141_, _03140_, _03138_);
  and (_03142_, _03141_, _02445_);
  or (_03143_, _03142_, _03137_);
  or (_03145_, _03143_, _02421_);
  and (_03146_, _03145_, _02414_);
  and (_03147_, _03146_, _03133_);
  or (_03148_, _03147_, _03120_);
  and (_03149_, _03148_, _02398_);
  or (_03150_, _03149_, _03095_);
  and (_03151_, _03150_, _02546_);
  or (_03152_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_03153_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and (_03154_, _03153_, _03152_);
  and (_03155_, _03154_, _02393_);
  or (_03156_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_03157_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_03158_, _03157_, _03156_);
  and (_03159_, _03158_, _02445_);
  or (_03161_, _03159_, _03155_);
  and (_03162_, _03161_, _02459_);
  or (_03163_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_03165_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_03166_, _03165_, _03163_);
  and (_03167_, _03166_, _02393_);
  or (_03169_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or (_03170_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_03171_, _03170_, _03169_);
  and (_03172_, _03171_, _02445_);
  or (_03173_, _03172_, _03167_);
  and (_03174_, _03173_, _02421_);
  or (_03176_, _03174_, _03162_);
  and (_03178_, _03176_, _02414_);
  and (_03179_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_03180_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or (_03181_, _03180_, _03179_);
  and (_03182_, _03181_, _02393_);
  and (_03183_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_03184_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_03185_, _03184_, _03183_);
  and (_03186_, _03185_, _02445_);
  or (_03187_, _03186_, _03182_);
  and (_03188_, _03187_, _02459_);
  and (_03189_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_03190_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_03191_, _03190_, _03189_);
  and (_03192_, _03191_, _02393_);
  and (_03193_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_03195_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or (_03196_, _03195_, _03193_);
  and (_03197_, _03196_, _02445_);
  or (_03198_, _03197_, _03192_);
  and (_03200_, _03198_, _02421_);
  or (_03201_, _03200_, _03188_);
  and (_03202_, _03201_, _02458_);
  or (_03203_, _03202_, _03178_);
  and (_03204_, _03203_, _02398_);
  or (_03205_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_03206_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and (_03207_, _03206_, _02445_);
  and (_03208_, _03207_, _03205_);
  or (_03210_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_03212_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and (_03213_, _03212_, _02393_);
  and (_03214_, _03213_, _03210_);
  or (_03215_, _03214_, _03208_);
  and (_03216_, _03215_, _02459_);
  or (_03217_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_03218_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and (_03219_, _03218_, _02445_);
  and (_03220_, _03219_, _03217_);
  or (_03221_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_03223_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and (_03224_, _03223_, _02393_);
  and (_03226_, _03224_, _03221_);
  or (_03228_, _03226_, _03220_);
  and (_03229_, _03228_, _02421_);
  or (_03230_, _03229_, _03216_);
  and (_03232_, _03230_, _02414_);
  and (_03234_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and (_03235_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_03236_, _03235_, _03234_);
  and (_03237_, _03236_, _02393_);
  and (_03238_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and (_03239_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_03240_, _03239_, _03238_);
  and (_03241_, _03240_, _02445_);
  or (_03242_, _03241_, _03237_);
  and (_03243_, _03242_, _02459_);
  and (_03245_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and (_03246_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_03247_, _03246_, _03245_);
  and (_03248_, _03247_, _02393_);
  and (_03249_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and (_03250_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_03251_, _03250_, _03249_);
  and (_03252_, _03251_, _02445_);
  or (_03253_, _03252_, _03248_);
  and (_03254_, _03253_, _02421_);
  or (_03255_, _03254_, _03243_);
  and (_03256_, _03255_, _02458_);
  or (_03257_, _03256_, _03232_);
  and (_03258_, _03257_, _02496_);
  or (_03259_, _03258_, _03204_);
  and (_03260_, _03259_, _02400_);
  or (_03261_, _03260_, _03151_);
  or (_03262_, _03261_, _02646_);
  and (_03263_, _03262_, _03045_);
  and (_03264_, _03263_, _26777_);
  or (_03265_, _03264_, _02841_);
  or (_03266_, _03265_, _02443_);
  not (_03267_, _02443_);
  or (_03268_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_03269_, _03268_, _22762_);
  and (_22712_, _03269_, _03266_);
  and (_03271_, _02374_, _23649_);
  and (_03272_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or (_22713_, _03272_, _03271_);
  or (_03273_, _02268_, _24537_);
  and (_03274_, _26625_, _24584_);
  and (_03275_, _25621_, _26582_);
  or (_03276_, _03275_, _24585_);
  or (_03277_, _03276_, _03274_);
  or (_03278_, _03277_, _03273_);
  and (_03279_, _03278_, _22768_);
  and (_03280_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  or (_03281_, _03280_, _25664_);
  or (_03283_, _03281_, _03279_);
  and (_26866_[1], _03283_, _22762_);
  and (_03284_, _25656_, _23898_);
  and (_03285_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_22714_, _03285_, _03284_);
  and (_03286_, _25142_, _23946_);
  and (_03288_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or (_22715_, _03288_, _03286_);
  and (_03290_, _02350_, _23747_);
  and (_03292_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_26978_, _03292_, _03290_);
  and (_03293_, _25649_, _23747_);
  and (_03295_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_22716_, _03295_, _03293_);
  and (_03296_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  and (_03297_, _02245_, _23747_);
  or (_22717_, _03297_, _03296_);
  and (_03298_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and (_03299_, _02245_, _23824_);
  or (_22718_, _03299_, _03298_);
  and (_03300_, _23752_, _23664_);
  and (_03301_, _03300_, _23747_);
  not (_03302_, _03300_);
  and (_03303_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_22719_, _03303_, _03301_);
  and (_03305_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _22762_);
  and (_03306_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _22762_);
  and (_03307_, _03306_, _01772_);
  or (_26895_[7], _03307_, _03305_);
  or (_03308_, _26622_, _26646_);
  and (_03309_, _26645_, _24613_);
  and (_03311_, _24597_, _24538_);
  and (_03312_, _03311_, _25667_);
  or (_03313_, _03312_, _03309_);
  or (_03314_, _03313_, _03308_);
  or (_03315_, _26669_, _26657_);
  or (_03316_, _26581_, _26615_);
  or (_03317_, _26636_, _26665_);
  or (_03318_, _03317_, _03316_);
  or (_03319_, _03318_, _03315_);
  or (_03320_, _03319_, _03314_);
  and (_03321_, _26568_, _24538_);
  and (_03322_, _24552_, _24445_);
  or (_03323_, _03322_, _03321_);
  or (_03324_, _26661_, _24608_);
  or (_03325_, _03324_, _03323_);
  or (_03327_, _03325_, _03320_);
  and (_03328_, _03327_, _22768_);
  and (_03329_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_03330_, _03321_, _03309_);
  and (_03331_, _03330_, _24566_);
  or (_03332_, _03331_, _25664_);
  and (_03334_, _26645_, _24567_);
  and (_03335_, _03334_, _24566_);
  or (_03336_, _03335_, _03332_);
  or (_03337_, _03336_, _03329_);
  or (_03338_, _03337_, _03328_);
  and (_26868_[0], _03338_, _22762_);
  and (_03339_, _01809_, _24282_);
  and (_03340_, _03339_, _23649_);
  not (_03342_, _03339_);
  and (_03343_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_22720_, _03343_, _03340_);
  and (_03344_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_03345_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_03347_, _03345_, _03344_);
  and (_03348_, _03347_, _02393_);
  and (_03349_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and (_03350_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or (_03351_, _03350_, _03349_);
  and (_03352_, _03351_, _02445_);
  or (_03353_, _03352_, _03348_);
  and (_03354_, _03353_, _02421_);
  and (_03355_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_03356_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_03358_, _03356_, _03355_);
  and (_03359_, _03358_, _02393_);
  and (_03360_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and (_03361_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or (_03363_, _03361_, _03360_);
  and (_03364_, _03363_, _02445_);
  or (_03366_, _03364_, _03359_);
  and (_03367_, _03366_, _02459_);
  or (_03368_, _03367_, _03354_);
  and (_03369_, _03368_, _02458_);
  or (_03370_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or (_03372_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_03373_, _03372_, _03370_);
  and (_03374_, _03373_, _02393_);
  or (_03375_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_03376_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_03377_, _03376_, _03375_);
  and (_03378_, _03377_, _02445_);
  or (_03379_, _03378_, _03374_);
  and (_03380_, _03379_, _02421_);
  or (_03381_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or (_03382_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_03383_, _03382_, _03381_);
  and (_03384_, _03383_, _02393_);
  or (_03385_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or (_03386_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_03387_, _03386_, _03385_);
  and (_03388_, _03387_, _02445_);
  or (_03389_, _03388_, _03384_);
  and (_03390_, _03389_, _02459_);
  or (_03392_, _03390_, _03380_);
  and (_03393_, _03392_, _02414_);
  or (_03394_, _03393_, _03369_);
  and (_03395_, _03394_, _02398_);
  and (_03396_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and (_03397_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or (_03399_, _03397_, _03396_);
  and (_03401_, _03399_, _02393_);
  and (_03402_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and (_03403_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_03404_, _03403_, _03402_);
  and (_03405_, _03404_, _02445_);
  or (_03407_, _03405_, _03401_);
  and (_03408_, _03407_, _02421_);
  and (_03410_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and (_03411_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or (_03412_, _03411_, _03410_);
  and (_03413_, _03412_, _02393_);
  and (_03414_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and (_03415_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or (_03416_, _03415_, _03414_);
  and (_03417_, _03416_, _02445_);
  or (_03419_, _03417_, _03413_);
  and (_03420_, _03419_, _02459_);
  or (_03421_, _03420_, _03408_);
  and (_03422_, _03421_, _02458_);
  or (_03423_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or (_03424_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and (_03425_, _03424_, _02445_);
  and (_03426_, _03425_, _03423_);
  or (_03427_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_03428_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and (_03429_, _03428_, _02393_);
  and (_03430_, _03429_, _03427_);
  or (_03431_, _03430_, _03426_);
  and (_03432_, _03431_, _02421_);
  or (_03434_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_03435_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and (_03437_, _03435_, _02445_);
  and (_03438_, _03437_, _03434_);
  or (_03440_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or (_03442_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and (_03443_, _03442_, _02393_);
  and (_03445_, _03443_, _03440_);
  or (_03446_, _03445_, _03438_);
  and (_03447_, _03446_, _02459_);
  or (_03449_, _03447_, _03432_);
  and (_03450_, _03449_, _02414_);
  or (_03451_, _03450_, _03422_);
  and (_03452_, _03451_, _02496_);
  or (_03454_, _03452_, _03395_);
  and (_03455_, _03454_, _02400_);
  and (_03456_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_03457_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or (_03458_, _03457_, _03456_);
  and (_03459_, _03458_, _02393_);
  and (_03460_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_03461_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or (_03462_, _03461_, _03460_);
  and (_03464_, _03462_, _02445_);
  or (_03465_, _03464_, _03459_);
  or (_03466_, _03465_, _02459_);
  and (_03467_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_03468_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or (_03469_, _03468_, _03467_);
  and (_03470_, _03469_, _02393_);
  and (_03471_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_03472_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or (_03473_, _03472_, _03471_);
  and (_03474_, _03473_, _02445_);
  or (_03475_, _03474_, _03470_);
  or (_03476_, _03475_, _02421_);
  and (_03478_, _03476_, _02458_);
  and (_03479_, _03478_, _03466_);
  or (_03480_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or (_03481_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_03482_, _03481_, _02445_);
  and (_03483_, _03482_, _03480_);
  or (_03484_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or (_03485_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_03487_, _03485_, _02393_);
  and (_03488_, _03487_, _03484_);
  or (_03489_, _03488_, _03483_);
  or (_03490_, _03489_, _02459_);
  or (_03491_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or (_03492_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_03493_, _03492_, _02445_);
  and (_03494_, _03493_, _03491_);
  or (_03495_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or (_03496_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_03497_, _03496_, _02393_);
  and (_03498_, _03497_, _03495_);
  or (_03499_, _03498_, _03494_);
  or (_03501_, _03499_, _02421_);
  and (_03502_, _03501_, _02414_);
  and (_03503_, _03502_, _03490_);
  or (_03504_, _03503_, _03479_);
  and (_03506_, _03504_, _02496_);
  and (_03507_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and (_03508_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_03510_, _03508_, _03507_);
  and (_03511_, _03510_, _02393_);
  and (_03512_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and (_03513_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_03514_, _03513_, _03512_);
  and (_03515_, _03514_, _02445_);
  or (_03516_, _03515_, _03511_);
  or (_03517_, _03516_, _02459_);
  and (_03519_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and (_03520_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_03521_, _03520_, _03519_);
  and (_03522_, _03521_, _02393_);
  and (_03523_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and (_03525_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_03526_, _03525_, _03523_);
  and (_03527_, _03526_, _02445_);
  or (_03528_, _03527_, _03522_);
  or (_03529_, _03528_, _02421_);
  and (_03530_, _03529_, _02458_);
  and (_03531_, _03530_, _03517_);
  or (_03532_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_03533_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and (_03534_, _03533_, _03532_);
  and (_03535_, _03534_, _02393_);
  or (_03536_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_03537_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and (_03538_, _03537_, _03536_);
  and (_03540_, _03538_, _02445_);
  or (_03541_, _03540_, _03535_);
  or (_03543_, _03541_, _02459_);
  or (_03544_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_03545_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and (_03546_, _03545_, _03544_);
  and (_03547_, _03546_, _02393_);
  or (_03548_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_03549_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and (_03550_, _03549_, _03548_);
  and (_03551_, _03550_, _02445_);
  or (_03552_, _03551_, _03547_);
  or (_03553_, _03552_, _02421_);
  and (_03554_, _03553_, _02414_);
  and (_03555_, _03554_, _03543_);
  or (_03556_, _03555_, _03531_);
  and (_03558_, _03556_, _02398_);
  or (_03559_, _03558_, _03506_);
  and (_03560_, _03559_, _02546_);
  or (_03561_, _03560_, _03455_);
  and (_03562_, _03561_, _02646_);
  or (_03563_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_03564_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and (_03565_, _03564_, _02445_);
  and (_03566_, _03565_, _03563_);
  or (_03567_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_03568_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and (_03569_, _03568_, _02393_);
  and (_03570_, _03569_, _03567_);
  or (_03571_, _03570_, _03566_);
  and (_03572_, _03571_, _02459_);
  or (_03573_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_03575_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and (_03576_, _03575_, _02445_);
  and (_03578_, _03576_, _03573_);
  or (_03579_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_03580_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and (_03581_, _03580_, _02393_);
  and (_03582_, _03581_, _03579_);
  or (_03583_, _03582_, _03578_);
  and (_03584_, _03583_, _02421_);
  or (_03585_, _03584_, _03572_);
  and (_03586_, _03585_, _02414_);
  and (_03587_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and (_03588_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_03589_, _03588_, _03587_);
  and (_03590_, _03589_, _02393_);
  and (_03591_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and (_03592_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_03593_, _03592_, _03591_);
  and (_03594_, _03593_, _02445_);
  or (_03595_, _03594_, _03590_);
  and (_03596_, _03595_, _02459_);
  and (_03597_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and (_03598_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_03599_, _03598_, _03597_);
  and (_03600_, _03599_, _02393_);
  and (_03601_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and (_03602_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_03603_, _03602_, _03601_);
  and (_03604_, _03603_, _02445_);
  or (_03606_, _03604_, _03600_);
  and (_03607_, _03606_, _02421_);
  or (_03609_, _03607_, _03596_);
  and (_03610_, _03609_, _02458_);
  or (_03611_, _03610_, _03586_);
  and (_03612_, _03611_, _02496_);
  or (_03614_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_03615_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and (_03616_, _03615_, _03614_);
  and (_03617_, _03616_, _02393_);
  or (_03618_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or (_03619_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_03620_, _03619_, _03618_);
  and (_03621_, _03620_, _02445_);
  or (_03622_, _03621_, _03617_);
  and (_03623_, _03622_, _02459_);
  or (_03624_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or (_03625_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and (_03626_, _03625_, _03624_);
  and (_03627_, _03626_, _02393_);
  or (_03629_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or (_03630_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_03631_, _03630_, _03629_);
  and (_03632_, _03631_, _02445_);
  or (_03633_, _03632_, _03627_);
  and (_03634_, _03633_, _02421_);
  or (_03635_, _03634_, _03623_);
  and (_03636_, _03635_, _02414_);
  and (_03637_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_03639_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_03640_, _03639_, _03637_);
  and (_03641_, _03640_, _02393_);
  and (_03642_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and (_03643_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or (_03644_, _03643_, _03642_);
  and (_03645_, _03644_, _02445_);
  or (_03646_, _03645_, _03641_);
  and (_03647_, _03646_, _02459_);
  and (_03648_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and (_03649_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or (_03650_, _03649_, _03648_);
  and (_03651_, _03650_, _02393_);
  and (_03652_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_03653_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_03654_, _03653_, _03652_);
  and (_03655_, _03654_, _02445_);
  or (_03657_, _03655_, _03651_);
  and (_03658_, _03657_, _02421_);
  or (_03659_, _03658_, _03647_);
  and (_03660_, _03659_, _02458_);
  or (_03661_, _03660_, _03636_);
  and (_03662_, _03661_, _02398_);
  or (_03663_, _03662_, _03612_);
  and (_03665_, _03663_, _02400_);
  and (_03666_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and (_03667_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_03668_, _03667_, _03666_);
  and (_03669_, _03668_, _02393_);
  and (_03670_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and (_03671_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_03672_, _03671_, _03670_);
  and (_03673_, _03672_, _02445_);
  or (_03674_, _03673_, _03669_);
  or (_03675_, _03674_, _02459_);
  and (_03677_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_03678_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_03679_, _03678_, _03677_);
  and (_03681_, _03679_, _02393_);
  and (_03682_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and (_03684_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_03685_, _03684_, _03682_);
  and (_03686_, _03685_, _02445_);
  or (_03687_, _03686_, _03681_);
  or (_03688_, _03687_, _02421_);
  and (_03689_, _03688_, _02458_);
  and (_03690_, _03689_, _03675_);
  or (_03691_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_03692_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and (_03693_, _03692_, _03691_);
  and (_03694_, _03693_, _02393_);
  or (_03695_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_03696_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_03697_, _03696_, _03695_);
  and (_03698_, _03697_, _02445_);
  or (_03699_, _03698_, _03694_);
  or (_03700_, _03699_, _02459_);
  or (_03702_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_03704_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and (_03705_, _03704_, _03702_);
  and (_03706_, _03705_, _02393_);
  or (_03707_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_03708_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and (_03709_, _03708_, _03707_);
  and (_03711_, _03709_, _02445_);
  or (_03712_, _03711_, _03706_);
  or (_03714_, _03712_, _02421_);
  and (_03715_, _03714_, _02414_);
  and (_03716_, _03715_, _03700_);
  or (_03717_, _03716_, _03690_);
  and (_03718_, _03717_, _02398_);
  and (_03719_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and (_03720_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_03721_, _03720_, _03719_);
  and (_03722_, _03721_, _02393_);
  and (_03723_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and (_03725_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_03726_, _03725_, _03723_);
  and (_03727_, _03726_, _02445_);
  or (_03728_, _03727_, _03722_);
  or (_03729_, _03728_, _02459_);
  and (_03730_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and (_03731_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_03732_, _03731_, _03730_);
  and (_03733_, _03732_, _02393_);
  and (_03734_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and (_03735_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_03736_, _03735_, _03734_);
  and (_03737_, _03736_, _02445_);
  or (_03738_, _03737_, _03733_);
  or (_03739_, _03738_, _02421_);
  and (_03740_, _03739_, _02458_);
  and (_03741_, _03740_, _03729_);
  or (_03743_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_03744_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and (_03745_, _03744_, _02445_);
  and (_03746_, _03745_, _03743_);
  or (_03747_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_03749_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and (_03750_, _03749_, _02393_);
  and (_03752_, _03750_, _03747_);
  or (_03753_, _03752_, _03746_);
  or (_03754_, _03753_, _02459_);
  or (_03755_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_03756_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and (_03757_, _03756_, _02445_);
  and (_03758_, _03757_, _03755_);
  or (_03759_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_03760_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and (_03761_, _03760_, _02393_);
  and (_03762_, _03761_, _03759_);
  or (_03764_, _03762_, _03758_);
  or (_03766_, _03764_, _02421_);
  and (_03767_, _03766_, _02414_);
  and (_03769_, _03767_, _03754_);
  or (_03770_, _03769_, _03741_);
  and (_03771_, _03770_, _02496_);
  or (_03772_, _03771_, _03718_);
  and (_03773_, _03772_, _02546_);
  or (_03774_, _03773_, _03665_);
  and (_03776_, _03774_, _02405_);
  or (_03777_, _03776_, _03562_);
  and (_03778_, _03777_, _26777_);
  and (_03779_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and (_03780_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_03781_, _03780_, _03779_);
  and (_03782_, _03781_, _02393_);
  and (_03783_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and (_03784_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_03785_, _03784_, _03783_);
  and (_03786_, _03785_, _02445_);
  or (_03787_, _03786_, _03782_);
  and (_03789_, _03787_, _02421_);
  and (_03790_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and (_03791_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_03793_, _03791_, _03790_);
  and (_03794_, _03793_, _02393_);
  and (_03795_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and (_03796_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_03797_, _03796_, _03795_);
  and (_03798_, _03797_, _02445_);
  or (_03799_, _03798_, _03794_);
  and (_03800_, _03799_, _02459_);
  or (_03801_, _03800_, _03789_);
  and (_03803_, _03801_, _02458_);
  or (_03804_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_03805_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and (_03806_, _03805_, _03804_);
  and (_03807_, _03806_, _02393_);
  or (_03808_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_03810_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and (_03811_, _03810_, _03808_);
  and (_03812_, _03811_, _02445_);
  or (_03813_, _03812_, _03807_);
  and (_03814_, _03813_, _02421_);
  or (_03815_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_03816_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and (_03817_, _03816_, _03815_);
  and (_03818_, _03817_, _02393_);
  or (_03819_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_03820_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and (_03821_, _03820_, _03819_);
  and (_03823_, _03821_, _02445_);
  or (_03824_, _03823_, _03818_);
  and (_03825_, _03824_, _02459_);
  or (_03826_, _03825_, _03814_);
  and (_03827_, _03826_, _02414_);
  or (_03828_, _03827_, _03803_);
  and (_03829_, _03828_, _02398_);
  and (_03830_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_03831_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_03832_, _03831_, _03830_);
  and (_03833_, _03832_, _02393_);
  and (_03834_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_03835_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_03836_, _03835_, _03834_);
  and (_03837_, _03836_, _02445_);
  or (_03838_, _03837_, _03833_);
  and (_03839_, _03838_, _02421_);
  and (_03840_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_03841_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_03842_, _03841_, _03840_);
  and (_03843_, _03842_, _02393_);
  and (_03844_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_03845_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_03847_, _03845_, _03844_);
  and (_03848_, _03847_, _02445_);
  or (_03850_, _03848_, _03843_);
  and (_03851_, _03850_, _02459_);
  or (_03852_, _03851_, _03839_);
  and (_03853_, _03852_, _02458_);
  or (_03854_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_03856_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_03857_, _03856_, _02445_);
  and (_03858_, _03857_, _03854_);
  or (_03859_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_03860_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_03861_, _03860_, _02393_);
  and (_03862_, _03861_, _03859_);
  or (_03863_, _03862_, _03858_);
  and (_03864_, _03863_, _02421_);
  or (_03866_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_03867_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_03868_, _03867_, _02445_);
  and (_03869_, _03868_, _03866_);
  or (_03870_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_03872_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_03873_, _03872_, _02393_);
  and (_03874_, _03873_, _03870_);
  or (_03875_, _03874_, _03869_);
  and (_03876_, _03875_, _02459_);
  or (_03877_, _03876_, _03864_);
  and (_03879_, _03877_, _02414_);
  or (_03881_, _03879_, _03853_);
  and (_03882_, _03881_, _02496_);
  or (_03884_, _03882_, _03829_);
  and (_03885_, _03884_, _02400_);
  and (_03886_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and (_03887_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_03888_, _03887_, _03886_);
  and (_03889_, _03888_, _02393_);
  and (_03890_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and (_03891_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_03892_, _03891_, _03890_);
  and (_03893_, _03892_, _02445_);
  or (_03895_, _03893_, _03889_);
  or (_03896_, _03895_, _02459_);
  and (_03897_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and (_03898_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_03899_, _03898_, _03897_);
  and (_03900_, _03899_, _02393_);
  and (_03901_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and (_03902_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_03903_, _03902_, _03901_);
  and (_03904_, _03903_, _02445_);
  or (_03905_, _03904_, _03900_);
  or (_03906_, _03905_, _02421_);
  and (_03907_, _03906_, _02458_);
  and (_03908_, _03907_, _03896_);
  or (_03909_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_03910_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and (_03911_, _03910_, _02445_);
  and (_03912_, _03911_, _03909_);
  or (_03913_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_03914_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and (_03915_, _03914_, _02393_);
  and (_03916_, _03915_, _03913_);
  or (_03917_, _03916_, _03912_);
  or (_03918_, _03917_, _02459_);
  or (_03919_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_03920_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and (_03921_, _03920_, _02445_);
  and (_03922_, _03921_, _03919_);
  or (_03923_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_03924_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and (_03925_, _03924_, _02393_);
  and (_03926_, _03925_, _03923_);
  or (_03927_, _03926_, _03922_);
  or (_03928_, _03927_, _02421_);
  and (_03929_, _03928_, _02414_);
  and (_03930_, _03929_, _03918_);
  or (_03931_, _03930_, _03908_);
  and (_03932_, _03931_, _02496_);
  and (_03933_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and (_03934_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_03935_, _03934_, _03933_);
  and (_03937_, _03935_, _02393_);
  and (_03938_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and (_03939_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_03940_, _03939_, _03938_);
  and (_03941_, _03940_, _02445_);
  or (_03942_, _03941_, _03937_);
  or (_03943_, _03942_, _02459_);
  and (_03944_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and (_03945_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_03946_, _03945_, _03944_);
  and (_03947_, _03946_, _02393_);
  and (_03948_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and (_03949_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_03950_, _03949_, _03948_);
  and (_03951_, _03950_, _02445_);
  or (_03952_, _03951_, _03947_);
  or (_03953_, _03952_, _02421_);
  and (_03954_, _03953_, _02458_);
  and (_03955_, _03954_, _03943_);
  or (_03956_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_03957_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and (_03958_, _03957_, _03956_);
  and (_03959_, _03958_, _02393_);
  or (_03960_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_03961_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and (_03962_, _03961_, _03960_);
  and (_03963_, _03962_, _02445_);
  or (_03964_, _03963_, _03959_);
  or (_03965_, _03964_, _02459_);
  or (_03966_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_03967_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and (_03968_, _03967_, _03966_);
  and (_03970_, _03968_, _02393_);
  or (_03971_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_03972_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and (_03973_, _03972_, _03971_);
  and (_03974_, _03973_, _02445_);
  or (_03975_, _03974_, _03970_);
  or (_03976_, _03975_, _02421_);
  and (_03977_, _03976_, _02414_);
  and (_03978_, _03977_, _03965_);
  or (_03979_, _03978_, _03955_);
  and (_03981_, _03979_, _02398_);
  or (_03982_, _03981_, _03932_);
  and (_03983_, _03982_, _02546_);
  or (_03985_, _03983_, _03885_);
  and (_03986_, _03985_, _02646_);
  or (_03988_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_03989_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and (_03990_, _03989_, _02445_);
  and (_03991_, _03990_, _03988_);
  or (_03992_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_03993_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and (_03994_, _03993_, _02393_);
  and (_03996_, _03994_, _03992_);
  or (_03998_, _03996_, _03991_);
  and (_03999_, _03998_, _02459_);
  or (_04000_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_04001_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and (_04002_, _04001_, _02445_);
  and (_04004_, _04002_, _04000_);
  or (_04005_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_04006_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and (_04008_, _04006_, _02393_);
  and (_04009_, _04008_, _04005_);
  or (_04010_, _04009_, _04004_);
  and (_04011_, _04010_, _02421_);
  or (_04012_, _04011_, _03999_);
  and (_04013_, _04012_, _02414_);
  and (_04014_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and (_04015_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_04016_, _04015_, _04014_);
  and (_04017_, _04016_, _02393_);
  and (_04018_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and (_04019_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_04020_, _04019_, _04018_);
  and (_04021_, _04020_, _02445_);
  or (_04022_, _04021_, _04017_);
  and (_04023_, _04022_, _02459_);
  and (_04024_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and (_04026_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_04027_, _04026_, _04024_);
  and (_04028_, _04027_, _02393_);
  and (_04029_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and (_04030_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_04032_, _04030_, _04029_);
  and (_04034_, _04032_, _02445_);
  or (_04035_, _04034_, _04028_);
  and (_04036_, _04035_, _02421_);
  or (_04037_, _04036_, _04023_);
  and (_04038_, _04037_, _02458_);
  or (_04039_, _04038_, _04013_);
  and (_04040_, _04039_, _02496_);
  or (_04041_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_04042_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and (_04043_, _04042_, _04041_);
  and (_04044_, _04043_, _02393_);
  or (_04046_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_04047_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and (_04048_, _04047_, _04046_);
  and (_04050_, _04048_, _02445_);
  or (_04051_, _04050_, _04044_);
  and (_04052_, _04051_, _02459_);
  or (_04053_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_04054_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and (_04055_, _04054_, _04053_);
  and (_04056_, _04055_, _02393_);
  or (_04057_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_04058_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and (_04059_, _04058_, _04057_);
  and (_04060_, _04059_, _02445_);
  or (_04061_, _04060_, _04056_);
  and (_04062_, _04061_, _02421_);
  or (_04063_, _04062_, _04052_);
  and (_04064_, _04063_, _02414_);
  and (_04065_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and (_04066_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_04067_, _04066_, _04065_);
  and (_04068_, _04067_, _02393_);
  and (_04069_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and (_04070_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_04071_, _04070_, _04069_);
  and (_04072_, _04071_, _02445_);
  or (_04073_, _04072_, _04068_);
  and (_04074_, _04073_, _02459_);
  and (_04075_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and (_04076_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_04077_, _04076_, _04075_);
  and (_04078_, _04077_, _02393_);
  and (_04079_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and (_04081_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_04082_, _04081_, _04079_);
  and (_04083_, _04082_, _02445_);
  or (_04084_, _04083_, _04078_);
  and (_04085_, _04084_, _02421_);
  or (_04086_, _04085_, _04074_);
  and (_04087_, _04086_, _02458_);
  or (_04088_, _04087_, _04064_);
  and (_04089_, _04088_, _02398_);
  or (_04091_, _04089_, _04040_);
  and (_04092_, _04091_, _02400_);
  and (_04093_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and (_04094_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_04095_, _04094_, _04093_);
  and (_04096_, _04095_, _02393_);
  and (_04097_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and (_04099_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_04100_, _04099_, _04097_);
  and (_04101_, _04100_, _02445_);
  or (_04102_, _04101_, _04096_);
  or (_04103_, _04102_, _02459_);
  and (_04104_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and (_04105_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_04106_, _04105_, _04104_);
  and (_04107_, _04106_, _02393_);
  and (_04108_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and (_04109_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_04110_, _04109_, _04108_);
  and (_04112_, _04110_, _02445_);
  or (_04113_, _04112_, _04107_);
  or (_04115_, _04113_, _02421_);
  and (_04116_, _04115_, _02458_);
  and (_04118_, _04116_, _04103_);
  or (_04119_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_04121_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and (_04122_, _04121_, _04119_);
  and (_04123_, _04122_, _02393_);
  or (_04124_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_04126_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and (_04127_, _04126_, _04124_);
  and (_04128_, _04127_, _02445_);
  or (_04129_, _04128_, _04123_);
  or (_04130_, _04129_, _02459_);
  or (_04131_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_04132_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and (_04134_, _04132_, _04131_);
  and (_04135_, _04134_, _02393_);
  or (_04136_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_04137_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and (_04138_, _04137_, _04136_);
  and (_04139_, _04138_, _02445_);
  or (_04141_, _04139_, _04135_);
  or (_04142_, _04141_, _02421_);
  and (_04143_, _04142_, _02414_);
  and (_04144_, _04143_, _04130_);
  or (_04145_, _04144_, _04118_);
  and (_04146_, _04145_, _02398_);
  and (_04147_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and (_04148_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_04149_, _04148_, _04147_);
  and (_04150_, _04149_, _02393_);
  and (_04151_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and (_04152_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_04153_, _04152_, _04151_);
  and (_04154_, _04153_, _02445_);
  or (_04155_, _04154_, _04150_);
  or (_04156_, _04155_, _02459_);
  and (_04157_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and (_04158_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_04159_, _04158_, _04157_);
  and (_04160_, _04159_, _02393_);
  and (_04161_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and (_04162_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_04163_, _04162_, _04161_);
  and (_04164_, _04163_, _02445_);
  or (_04165_, _04164_, _04160_);
  or (_04166_, _04165_, _02421_);
  and (_04167_, _04166_, _02458_);
  and (_04168_, _04167_, _04156_);
  or (_04169_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_04170_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and (_04172_, _04170_, _02445_);
  and (_04173_, _04172_, _04169_);
  or (_04175_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_04176_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and (_04177_, _04176_, _02393_);
  and (_04178_, _04177_, _04175_);
  or (_04179_, _04178_, _04173_);
  or (_04180_, _04179_, _02459_);
  or (_04181_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_04182_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and (_04183_, _04182_, _02445_);
  and (_04184_, _04183_, _04181_);
  or (_04185_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_04186_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and (_04187_, _04186_, _02393_);
  and (_04188_, _04187_, _04185_);
  or (_04189_, _04188_, _04184_);
  or (_04190_, _04189_, _02421_);
  and (_04191_, _04190_, _02414_);
  and (_04192_, _04191_, _04180_);
  or (_04194_, _04192_, _04168_);
  and (_04196_, _04194_, _02496_);
  or (_04197_, _04196_, _04146_);
  and (_04198_, _04197_, _02546_);
  or (_04200_, _04198_, _04092_);
  and (_04201_, _04200_, _02405_);
  or (_04202_, _04201_, _03986_);
  and (_04204_, _04202_, _02444_);
  or (_04205_, _04204_, _03778_);
  or (_04206_, _04205_, _02443_);
  or (_04207_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_04208_, _04207_, _22762_);
  and (_22721_, _04208_, _04206_);
  nor (_04210_, _01772_, rst);
  nand (_04211_, _22768_, _01532_);
  and (_26893_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _22762_);
  and (_04213_, _26893_, _04211_);
  or (_26894_, _04213_, _04210_);
  and (_04215_, _03339_, _23824_);
  and (_04216_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_27112_, _04216_, _04215_);
  and (_04218_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  and (_04219_, _02298_, _24050_);
  or (_27237_, _04219_, _04218_);
  and (_04220_, _25656_, _23824_);
  and (_04221_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_22723_, _04221_, _04220_);
  and (_04222_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _22762_);
  and (_04223_, _04222_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_04224_, _01744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_04226_, _01744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_04227_, _04226_, _04224_);
  not (_04228_, _04227_);
  nor (_04229_, _04228_, _01747_);
  and (_04230_, _04228_, _01747_);
  or (_04231_, _04230_, _04229_);
  or (_04232_, _04231_, _25729_);
  or (_04233_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_04234_, _04233_, _01793_);
  and (_04235_, _04234_, _04232_);
  or (_26891_[15], _04235_, _04223_);
  and (_04236_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  and (_04237_, _02306_, _23898_);
  or (_22724_, _04237_, _04236_);
  and (_04239_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_04240_, _04239_, _03332_);
  and (_04241_, _04240_, _22762_);
  and (_04242_, _03311_, _24581_);
  or (_04243_, _04242_, _24617_);
  or (_04244_, _04243_, _26616_);
  and (_04245_, _26621_, _24471_);
  or (_04247_, _04245_, _24585_);
  or (_04248_, _04247_, _03330_);
  or (_04249_, _04248_, _04244_);
  and (_04250_, _04249_, _25644_);
  or (_26868_[1], _04250_, _04241_);
  and (_26889_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _22762_);
  and (_04251_, _03339_, _23778_);
  and (_04252_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_22725_, _04252_, _04251_);
  and (_04253_, _02350_, _23707_);
  and (_04254_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_22726_, _04254_, _04253_);
  and (_04255_, _02350_, _24050_);
  and (_04256_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_22727_, _04256_, _04255_);
  nand (_04257_, _00886_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_04259_, _04257_, _01213_);
  and (_04260_, _04259_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_04261_, _01216_, _23185_);
  and (_04262_, _04261_, _23149_);
  or (_04263_, _04262_, _04260_);
  nand (_04264_, _04263_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_04265_, _04263_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_04266_, _04265_, _00401_);
  and (_04267_, _04266_, _04264_);
  and (_04268_, _00875_, _24628_);
  nor (_04269_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_04271_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23095_);
  nor (_04272_, _04271_, _04269_);
  nor (_04273_, _04272_, _01283_);
  and (_04274_, _04272_, _01283_);
  or (_04276_, _04274_, _04273_);
  and (_04277_, _04276_, _23480_);
  or (_04278_, _26521_, _26481_);
  and (_04279_, _04278_, _26522_);
  and (_04280_, _04279_, _23596_);
  and (_04281_, _01294_, _23179_);
  nor (_04282_, _04281_, _01293_);
  nor (_04283_, _04282_, _01302_);
  nand (_04284_, _04283_, _23142_);
  or (_04285_, _04283_, _23142_);
  and (_04286_, _04285_, _23609_);
  and (_04287_, _04286_, _04284_);
  and (_04288_, _23521_, _23142_);
  or (_04289_, _04288_, _23537_);
  and (_04290_, _04289_, _23627_);
  and (_04291_, _00611_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_04292_, _23579_, _23142_);
  and (_04293_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  or (_04294_, _04293_, _04292_);
  or (_04295_, _04294_, _04291_);
  or (_04296_, _04295_, _04290_);
  or (_04297_, _04296_, _04287_);
  or (_04298_, _04297_, _04280_);
  or (_04299_, _04298_, _04277_);
  and (_04300_, _04299_, _26566_);
  nor (_04301_, _01343_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_04302_, _01343_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_04303_, _04302_, _04301_);
  nand (_04304_, _04303_, _01349_);
  or (_04305_, _04303_, _01349_);
  and (_04306_, _04305_, _04304_);
  and (_04307_, _04306_, _00405_);
  and (_04308_, _26573_, _26772_);
  or (_04309_, _04308_, _04307_);
  and (_04310_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_04311_, _04310_, _04309_);
  nor (_04312_, _04311_, _04300_);
  nand (_04313_, _04312_, _00289_);
  or (_04314_, _04313_, _04268_);
  or (_04315_, _04314_, _04267_);
  or (_04316_, _04303_, _00289_);
  and (_04317_, _04316_, _22762_);
  and (_26890_[15], _04317_, _04315_);
  nor (_04318_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_26892_, _04318_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  nor (_04319_, _23953_, _23950_);
  and (_04320_, _01801_, _01798_);
  nor (_04321_, _04320_, _23950_);
  and (_04322_, _04321_, _23840_);
  nor (_04323_, _04321_, _23840_);
  nor (_04324_, _04323_, _04322_);
  nor (_04325_, _04324_, _04319_);
  and (_04326_, _23856_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_04327_, _04326_, _04319_);
  and (_04328_, _04327_, _01517_);
  or (_04329_, _04328_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_04331_, _04329_, _04325_);
  and (_26896_[2], _04331_, _22762_);
  and (_04333_, _24812_, _24647_);
  and (_04334_, _04333_, _24705_);
  nand (_04335_, _04334_, _23594_);
  and (_04336_, _25769_, _23753_);
  and (_04337_, _04336_, _24735_);
  not (_04339_, _04337_);
  or (_04340_, _04334_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_04341_, _04340_, _04339_);
  and (_04342_, _04341_, _04335_);
  and (_04343_, _04337_, _24043_);
  or (_04344_, _04343_, _04342_);
  and (_22728_, _04344_, _22762_);
  and (_04346_, _04333_, _24125_);
  nand (_04347_, _04346_, _23594_);
  or (_04348_, _04346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_04349_, _04348_, _04339_);
  and (_04350_, _04349_, _04347_);
  and (_04351_, _04337_, _23939_);
  or (_04353_, _04351_, _04350_);
  and (_22729_, _04353_, _22762_);
  and (_04354_, _24746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_04356_, _04354_, _24745_);
  and (_04357_, _04356_, _04333_);
  not (_04358_, _04333_);
  or (_04360_, _04358_, _24752_);
  and (_04362_, _04360_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_04363_, _04362_, _04337_);
  or (_04365_, _04363_, _04357_);
  or (_04366_, _04339_, _23642_);
  and (_04367_, _04366_, _22762_);
  and (_22730_, _04367_, _04365_);
  and (_04368_, _04333_, _24118_);
  nand (_04369_, _04368_, _23594_);
  or (_04370_, _04368_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_04372_, _04370_, _04339_);
  and (_04373_, _04372_, _04369_);
  and (_04374_, _04337_, _23738_);
  or (_04375_, _04374_, _04373_);
  and (_22731_, _04375_, _22762_);
  nor (_04376_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_04377_, _04376_);
  nor (_04378_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_04380_, _04378_, _04377_);
  and (_04381_, _04380_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_04383_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_04384_, _04380_, _04383_);
  or (_04386_, _04384_, _04381_);
  or (_04387_, _04386_, _04333_);
  not (_04388_, _24291_);
  nor (_04389_, _04388_, _23594_);
  or (_04390_, _24291_, _04383_);
  nand (_04391_, _04390_, _04333_);
  or (_04392_, _04391_, _04389_);
  and (_04393_, _04392_, _04387_);
  or (_04394_, _04393_, _04337_);
  or (_04395_, _04339_, _23816_);
  and (_04396_, _04395_, _22762_);
  and (_22732_, _04396_, _04394_);
  not (_04397_, _24067_);
  nor (_04398_, _04397_, _23594_);
  nand (_04399_, _04397_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_04401_, _04399_, _04333_);
  or (_04402_, _04401_, _04398_);
  or (_04403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_04404_, _04403_, _04333_);
  and (_04405_, _04404_, _04402_);
  or (_04406_, _04405_, _04337_);
  or (_04407_, _04339_, _23892_);
  and (_04408_, _04407_, _22762_);
  and (_22733_, _04408_, _04406_);
  not (_04410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_04411_, _04410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_04413_, _04411_, _04376_);
  and (_04414_, _04413_, _04378_);
  or (_04415_, _04414_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_04417_, _04415_, _04333_);
  and (_04418_, _24678_, _23711_);
  not (_04420_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_04421_, _24678_, _04420_);
  nand (_04423_, _04421_, _04333_);
  or (_04424_, _04423_, _04418_);
  and (_04425_, _04424_, _04417_);
  or (_04426_, _04425_, _04337_);
  nand (_04427_, _04337_, _23772_);
  and (_04428_, _04427_, _22762_);
  and (_22734_, _04428_, _04426_);
  or (_04429_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_04430_, _04429_, _22762_);
  or (_04431_, _02037_, _24043_);
  and (_22735_, _04431_, _04430_);
  or (_04432_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_04433_, _04432_, _22762_);
  or (_04434_, _02037_, _23939_);
  and (_22736_, _04434_, _04433_);
  or (_04435_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_04436_, _04435_, _22762_);
  or (_04437_, _02037_, _23738_);
  and (_22737_, _04437_, _04436_);
  or (_04438_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_04439_, _04438_, _22762_);
  or (_04440_, _02037_, _23892_);
  and (_22738_, _04440_, _04439_);
  nand (_04441_, _02034_, _23772_);
  or (_04442_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_04443_, _04442_, _22762_);
  and (_22739_, _04443_, _04441_);
  and (_04444_, _02350_, _23946_);
  and (_04445_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_22740_, _04445_, _04444_);
  and (_04447_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_04448_, _04447_, _04376_);
  and (_04449_, _04377_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_04451_, _04449_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_04452_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_04453_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_04454_, _04453_, _04452_);
  and (_04455_, _04454_, _04451_);
  nor (_04457_, _04455_, _04448_);
  not (_04458_, _04457_);
  and (_04459_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_04460_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_04461_, _04460_, _04459_);
  and (_04462_, _04336_, _24072_);
  nor (_04463_, _04462_, _04461_);
  not (_04464_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_04465_, _04464_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_04466_, _04465_, _04377_);
  and (_04467_, _04466_, _04462_);
  or (_04469_, _04467_, _04463_);
  and (_22741_, _04469_, _22762_);
  and (_04470_, _04462_, _04377_);
  nand (_04471_, _04470_, _23702_);
  and (_04473_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_04474_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_04475_, _04474_, _04473_);
  or (_04476_, _04475_, _04462_);
  and (_04477_, _04476_, _22762_);
  and (_22742_, _04477_, _04471_);
  and (_04478_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_04479_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_04480_, _04479_, _04478_);
  nor (_04481_, _04480_, _04462_);
  and (_04483_, _04470_, _24043_);
  or (_04484_, _04483_, _04481_);
  and (_04485_, _04462_, _04376_);
  and (_04486_, _04485_, _26750_);
  or (_04487_, _04486_, _04484_);
  and (_22743_, _04487_, _22762_);
  not (_04488_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_04490_, _04462_, _04464_);
  and (_04491_, _04490_, _04488_);
  and (_04493_, _04491_, _24043_);
  and (_04494_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_04495_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_04496_, _04495_, _04494_);
  nor (_04497_, _04496_, _04462_);
  and (_04498_, _04470_, _23939_);
  or (_04500_, _04498_, _04497_);
  or (_04501_, _04500_, _04493_);
  and (_22744_, _04501_, _22762_);
  and (_04504_, _04491_, _23939_);
  and (_04505_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_04506_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_04507_, _04506_, _04505_);
  nor (_04508_, _04507_, _04462_);
  and (_04509_, _04470_, _23642_);
  or (_04510_, _04509_, _04508_);
  or (_04511_, _04510_, _04504_);
  and (_22745_, _04511_, _22762_);
  and (_04513_, _04491_, _23642_);
  and (_04514_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_04515_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_04516_, _04515_, _04514_);
  nor (_04517_, _04516_, _04462_);
  and (_04518_, _04470_, _23738_);
  or (_04520_, _04518_, _04517_);
  or (_04521_, _04520_, _04513_);
  and (_22747_, _04521_, _22762_);
  and (_04522_, _04470_, _23816_);
  and (_04523_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_04524_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_04525_, _04524_, _04523_);
  nor (_04526_, _04525_, _04462_);
  and (_04527_, _04491_, _23738_);
  or (_04528_, _04527_, _04526_);
  or (_04529_, _04528_, _04522_);
  and (_22748_, _04529_, _22762_);
  and (_04531_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_04532_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_04533_, _04532_, _04531_);
  nor (_04535_, _04533_, _04462_);
  and (_04536_, _04470_, _23892_);
  or (_04537_, _04536_, _04535_);
  and (_04538_, _04485_, _23816_);
  or (_04540_, _04538_, _04537_);
  and (_22749_, _04540_, _22762_);
  and (_04541_, _04491_, _23892_);
  and (_04543_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_04544_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_04545_, _04544_, _04543_);
  nor (_04547_, _04545_, _04462_);
  and (_04549_, _04470_, _24685_);
  or (_04551_, _04549_, _04547_);
  or (_04552_, _04551_, _04541_);
  and (_22750_, _04552_, _22762_);
  or (_04554_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_04555_, _04448_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_04556_, _04555_, _04455_);
  and (_04557_, _04556_, _04554_);
  nor (_04558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor (_04559_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_04560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_04561_, _04560_, _04559_);
  and (_04563_, _04561_, _04558_);
  nor (_04564_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_04565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_04567_, _04565_, _04564_);
  and (_04568_, _04567_, _04448_);
  and (_04569_, _04568_, _04563_);
  and (_04570_, _04569_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_04571_, _04570_, _04557_);
  nor (_04572_, _04571_, _04462_);
  and (_04574_, _04485_, _24685_);
  or (_04575_, _04574_, _04572_);
  and (_22751_, _04575_, _22762_);
  not (_04576_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_04578_, _04376_, _04576_);
  and (_04579_, _04578_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_04581_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_04582_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _04581_);
  not (_04584_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_04586_, _04584_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_04588_, _04586_, _04582_);
  and (_04589_, _04588_, _04579_);
  and (_04591_, _04576_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_04593_, _04376_, _04420_);
  and (_04594_, _04593_, _04591_);
  and (_04595_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_04596_, _04595_, _04377_);
  nor (_04598_, _04596_, _04594_);
  nor (_04599_, _04598_, _04579_);
  or (_04600_, _04599_, _04589_);
  and (_04601_, _04376_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_04602_, _04601_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_04603_, _04602_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_04604_, _04603_, _04600_);
  nor (_04605_, _04602_, _04589_);
  or (_04606_, _04605_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_04607_, _04606_, _02066_);
  and (_04608_, _04607_, _04604_);
  or (_22752_, _04608_, _02065_);
  not (_04609_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not (_04611_, _04605_);
  nor (_04612_, _04611_, _04599_);
  nor (_04613_, _04612_, _04609_);
  or (_04615_, _04613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_04616_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _04609_);
  or (_04618_, _04616_, _04605_);
  and (_04619_, _04618_, _22762_);
  and (_22753_, _04619_, _04615_);
  and (_04621_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  and (_04623_, _02245_, _23946_);
  or (_22754_, _04623_, _04621_);
  and (_04625_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_04627_, _04611_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  not (_04628_, _04579_);
  nor (_04629_, _04588_, _04628_);
  and (_04630_, _04629_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_04631_, _04596_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nand (_04632_, _04631_, _04628_);
  nor (_04633_, _04632_, _04594_);
  nor (_04634_, _04633_, _04630_);
  nor (_04636_, _04634_, _04602_);
  or (_04637_, _04636_, _04627_);
  and (_04639_, _04637_, _02066_);
  or (_22755_, _04639_, _04625_);
  and (_04641_, _01810_, _23946_);
  and (_04643_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_22756_, _04643_, _04641_);
  and (_04644_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and (_04646_, _02245_, _23649_);
  or (_27036_, _04646_, _04644_);
  and (_04648_, _25656_, _23649_);
  and (_04650_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_27192_, _04650_, _04648_);
  and (_04652_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  and (_04654_, _02298_, _23707_);
  or (_27238_, _04654_, _04652_);
  and (_04656_, _01758_, _23986_);
  and (_04658_, _04656_, _23707_);
  not (_04660_, _04656_);
  and (_04661_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_22758_, _04661_, _04658_);
  and (_04663_, _01478_, _01377_);
  or (_04665_, _04663_, _01474_);
  and (_04666_, _01487_, _01383_);
  and (_04667_, _01426_, _01362_);
  or (_04668_, _04667_, _04666_);
  or (_04669_, _04668_, _04665_);
  and (_04671_, _01422_, _01357_);
  and (_04673_, _01472_, _01425_);
  and (_04674_, _01368_, _01362_);
  or (_04675_, _04674_, _04673_);
  or (_04676_, _04675_, _04671_);
  or (_04677_, _01509_, _01491_);
  or (_04678_, _04677_, _01380_);
  or (_04679_, _04678_, _04676_);
  or (_04680_, _04679_, _04669_);
  and (_04681_, _01461_, _01401_);
  and (_04682_, _01401_, _01395_);
  or (_04683_, _01453_, _01376_);
  and (_04684_, _04683_, _01426_);
  or (_04685_, _04684_, _04682_);
  nor (_04686_, _04685_, _04681_);
  nand (_04688_, _04686_, _01436_);
  or (_04690_, _04688_, _04680_);
  and (_04691_, _04690_, _22769_);
  and (_04693_, _22765_, _22766_);
  and (_04694_, _04693_, _24564_);
  nor (_04695_, _04694_, _25661_);
  or (_04696_, _04695_, rst);
  or (_26863_[1], _04696_, _04691_);
  and (_04698_, _04656_, _24050_);
  and (_04700_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_22759_, _04700_, _04698_);
  not (_04701_, _04612_);
  or (_04702_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_04703_, _04605_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_04704_, _04703_, _02066_);
  and (_04705_, _04704_, _04702_);
  or (_22760_, _04705_, _02071_);
  and (_04706_, _02370_, _23824_);
  and (_04707_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_22761_, _04707_, _04706_);
  and (_04708_, _02200_, _23778_);
  and (_04709_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_22774_, _04709_, _04708_);
  and (_04711_, _04588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_04712_, _04711_, _04598_);
  or (_04714_, _04712_, _04612_);
  and (_04715_, _04714_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_04717_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _04609_);
  nand (_04718_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_04720_, _04718_, _04605_);
  or (_04721_, _04720_, _04717_);
  or (_04723_, _04721_, _04715_);
  and (_22776_, _04723_, _22762_);
  nor (_04724_, _04596_, _04579_);
  or (_04725_, _04724_, _04609_);
  or (_04726_, _04725_, _04584_);
  and (_04727_, _04579_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_04728_, _04727_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_04729_, _04728_, _22762_);
  and (_22779_, _04729_, _04726_);
  and (_04730_, _24331_, _24050_);
  and (_04732_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_22787_, _04732_, _04730_);
  nand (_04734_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22762_);
  nor (_04735_, _04734_, _04613_);
  or (_04736_, _04712_, _04611_);
  and (_04737_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_04738_, _04737_, _04736_);
  or (_22790_, _04738_, _04735_);
  and (_04740_, _04725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_04741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_04743_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_04744_, _04743_, _04741_);
  and (_04745_, _04744_, _04727_);
  or (_04746_, _04745_, _04740_);
  and (_22792_, _04746_, _22762_);
  and (_04748_, _01808_, _24766_);
  not (_04749_, _04748_);
  and (_04751_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and (_04752_, _04748_, _23707_);
  or (_22818_, _04752_, _04751_);
  or (_04754_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_04756_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_04757_, _04756_, rst);
  nand (_04758_, _04757_, _04754_);
  nor (_22831_, _04758_, _04462_);
  and (_04760_, _23788_, _23072_);
  and (_04761_, _04760_, _01808_);
  not (_04762_, _04761_);
  and (_04763_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and (_04764_, _04761_, _23649_);
  or (_22835_, _04764_, _04763_);
  and (_04766_, _04741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_04767_, _04766_, _04581_);
  and (_04768_, _04727_, _04767_);
  or (_04769_, _04768_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not (_04770_, rxd_i);
  nand (_04771_, _04768_, _04770_);
  and (_04772_, _04771_, _22762_);
  and (_22851_, _04772_, _04769_);
  or (_04773_, _04756_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_04774_, _04756_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_04775_, _04774_, rst);
  nand (_04776_, _04775_, _04773_);
  nor (_22856_, _04776_, _04462_);
  nor (_04778_, _04774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_04780_, _04774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_04781_, _04780_, _04778_);
  nand (_04782_, _04781_, _22762_);
  nor (_22858_, _04782_, _04462_);
  and (_04783_, _02350_, _23898_);
  and (_04785_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_22863_, _04785_, _04783_);
  and (_04786_, _24006_, _23747_);
  and (_04787_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  or (_22866_, _04787_, _04786_);
  or (_04788_, _04613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_04789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _04609_);
  or (_04790_, _04789_, _04605_);
  and (_04791_, _04790_, _22762_);
  and (_22873_, _04791_, _04788_);
  and (_04792_, _02350_, _23778_);
  and (_04793_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_22880_, _04793_, _04792_);
  and (_04794_, _01971_, _23824_);
  and (_04795_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  or (_22898_, _04795_, _04794_);
  and (_04797_, _01809_, _23069_);
  and (_04799_, _04797_, _23824_);
  not (_04800_, _04797_);
  and (_04801_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_22902_, _04801_, _04799_);
  and (_04804_, _04725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor (_04805_, _04766_, _04628_);
  or (_04806_, _04805_, _04804_);
  and (_04807_, _04741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_04809_, _04807_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_04810_, _04809_, _22762_);
  and (_22911_, _04810_, _04806_);
  and (_04811_, _23754_, _23069_);
  and (_04812_, _04811_, _23946_);
  not (_04813_, _04811_);
  and (_04814_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  or (_22916_, _04814_, _04812_);
  and (_04816_, _24699_, _23649_);
  and (_04817_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  or (_22925_, _04817_, _04816_);
  and (_04819_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_22933_, _04819_, _04625_);
  and (_04820_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and (_04821_, _02245_, _23778_);
  or (_22936_, _04821_, _04820_);
  and (_04822_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_04823_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_22955_, _04823_, _04822_);
  and (_04825_, _04656_, _23778_);
  and (_04826_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_22959_, _04826_, _04825_);
  and (_04828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_04829_, _04828_, _04717_);
  and (_22965_, _04829_, _22762_);
  and (_04830_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_04831_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_22988_, _04831_, _04830_);
  and (_04832_, _01758_, _23069_);
  and (_04833_, _04832_, _23707_);
  not (_04834_, _04832_);
  and (_04835_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_22993_, _04835_, _04833_);
  and (_04836_, _03300_, _23824_);
  and (_04838_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_22998_, _04838_, _04836_);
  or (_04839_, _04613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_04840_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _04609_);
  or (_04842_, _04840_, _04605_);
  and (_04843_, _04842_, _22762_);
  and (_23001_, _04843_, _04839_);
  or (_04845_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_04846_, _04605_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_04848_, _04846_, _02066_);
  and (_04850_, _04848_, _04845_);
  or (_23007_, _04850_, _02069_);
  or (_04852_, _04613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_04853_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _04609_);
  or (_04854_, _04853_, _04605_);
  and (_04855_, _04854_, _22762_);
  and (_23010_, _04855_, _04852_);
  or (_04856_, _04613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_04857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _04609_);
  or (_04858_, _04857_, _04605_);
  and (_04859_, _04858_, _22762_);
  and (_23013_, _04859_, _04856_);
  and (_04860_, _26099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_04861_, _04860_, _26100_);
  not (_04862_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_04863_, _26117_, _26114_);
  and (_04864_, _04863_, _26110_);
  and (_04866_, _04864_, _24308_);
  and (_04867_, _04866_, _26099_);
  nor (_04869_, _04867_, _04862_);
  and (_04871_, _04867_, _04862_);
  or (_04872_, _04871_, _04869_);
  and (_04873_, _04872_, _04861_);
  and (_04874_, _24308_, _24300_);
  and (_04876_, _04874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_04877_, _04874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_04878_, _04877_, _24302_);
  nor (_04879_, _04878_, _04876_);
  and (_04880_, _26115_, _24307_);
  and (_04881_, _04880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_04882_, _04881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_04883_, _04881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_04885_, _04883_, _26097_);
  nor (_04886_, _04885_, _04882_);
  or (_04887_, _04886_, _04879_);
  or (_04888_, _04887_, _04873_);
  or (_04890_, _04888_, _24299_);
  not (_04891_, _24299_);
  or (_04892_, _04891_, _23738_);
  and (_04894_, _04892_, _04890_);
  or (_04895_, _04894_, _24293_);
  nand (_04896_, _24293_, _04862_);
  and (_04897_, _04896_, _22762_);
  and (_23032_, _04897_, _04895_);
  and (_04898_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  and (_04900_, _04748_, _23747_);
  or (_23037_, _04900_, _04898_);
  and (_04901_, _04656_, _23747_);
  and (_04903_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_23119_, _04903_, _04901_);
  and (_04905_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and (_04907_, _04748_, _23946_);
  or (_27031_, _04907_, _04905_);
  and (_04908_, _04656_, _23824_);
  and (_04909_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_23125_, _04909_, _04908_);
  and (_04911_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  and (_04913_, _04748_, _23649_);
  or (_23136_, _04913_, _04911_);
  and (_04914_, _25142_, _24050_);
  and (_04915_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or (_23162_, _04915_, _04914_);
  and (_04917_, _01809_, _23911_);
  and (_04918_, _04917_, _23707_);
  not (_04919_, _04917_);
  and (_04920_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_23176_, _04920_, _04918_);
  and (_04922_, _23991_, _23754_);
  and (_04924_, _04922_, _23898_);
  not (_04925_, _04922_);
  and (_04926_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or (_23189_, _04926_, _04924_);
  and (_04927_, _03300_, _23898_);
  and (_04928_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_23207_, _04928_, _04927_);
  and (_04929_, _04832_, _23747_);
  and (_04931_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_23210_, _04931_, _04929_);
  and (_04934_, _04832_, _23824_);
  and (_04935_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_26942_, _04935_, _04934_);
  and (_04936_, _04797_, _23946_);
  and (_04937_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_23234_, _04937_, _04936_);
  and (_04938_, _26589_, _24597_);
  or (_04939_, _04938_, _24586_);
  or (_04940_, _04939_, _04242_);
  or (_04941_, _04940_, _03330_);
  and (_04942_, _24546_, _24445_);
  or (_04943_, _04942_, _24594_);
  or (_04944_, _04943_, _24591_);
  and (_04945_, _26582_, _24546_);
  and (_04946_, _03275_, _24612_);
  or (_04947_, _04946_, _04945_);
  or (_04948_, _04947_, _04944_);
  or (_04949_, _04948_, _04941_);
  and (_04950_, _24613_, _24589_);
  and (_04952_, _26650_, _24556_);
  and (_04953_, _24598_, _24538_);
  and (_04955_, _04953_, _25667_);
  or (_04956_, _04955_, _04952_);
  or (_04957_, _04956_, _04950_);
  and (_04958_, _24593_, _26582_);
  and (_04959_, _04958_, _24471_);
  or (_04961_, _04959_, _24542_);
  and (_04962_, _24592_, _24448_);
  and (_04964_, _24556_, _24540_);
  or (_04965_, _04964_, _04962_);
  or (_04966_, _04965_, _04961_);
  or (_04967_, _04966_, _04957_);
  or (_04968_, _04967_, _04949_);
  or (_04969_, _26583_, _25639_);
  and (_04970_, _04953_, _24556_);
  or (_04972_, _04970_, _24558_);
  or (_04973_, _24618_, _24616_);
  and (_04974_, _04973_, _24556_);
  or (_04976_, _04974_, _04972_);
  or (_04977_, _04976_, _04969_);
  and (_04978_, _26589_, _24588_);
  and (_04979_, _24593_, _24445_);
  or (_04980_, _04979_, _04978_);
  and (_04981_, _24545_, _24448_);
  and (_04982_, _24589_, _26582_);
  or (_04983_, _04982_, _04981_);
  and (_04984_, _00234_, _26582_);
  or (_04985_, _04984_, _24559_);
  or (_04987_, _04985_, _04983_);
  or (_04989_, _04987_, _04980_);
  or (_04991_, _04989_, _04977_);
  or (_04992_, _04991_, _04968_);
  and (_04993_, _04992_, _22768_);
  and (_04994_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_04995_, _25638_);
  nor (_04996_, _24567_, _24447_);
  nor (_04998_, _04996_, _04995_);
  nor (_05000_, _04998_, _04981_);
  not (_05001_, _05000_);
  and (_05003_, _05001_, _25662_);
  or (_05005_, _05003_, _24572_);
  or (_05006_, _05005_, _04994_);
  or (_05007_, _05006_, _04993_);
  and (_26869_[0], _05007_, _22762_);
  and (_05008_, _25078_, _23754_);
  and (_05009_, _05008_, _23946_);
  not (_05011_, _05008_);
  and (_05012_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_23248_, _05012_, _05009_);
  and (_05013_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and (_05014_, _01967_, _23707_);
  or (_23255_, _05014_, _05013_);
  or (_05016_, _04980_, _04962_);
  or (_05017_, _26654_, _26620_);
  and (_05018_, _05017_, _24408_);
  or (_05019_, _05018_, _05016_);
  or (_05020_, _05019_, _04948_);
  or (_05022_, _24559_, _24548_);
  or (_05023_, _03312_, _26629_);
  or (_05024_, _05023_, _05022_);
  and (_05025_, _04953_, _24581_);
  or (_05026_, _02268_, _26661_);
  or (_05027_, _05026_, _05025_);
  and (_05028_, _26589_, _24598_);
  or (_05029_, _05028_, _24586_);
  or (_05030_, _05029_, _24542_);
  or (_05031_, _05030_, _05027_);
  or (_05032_, _05031_, _05024_);
  or (_05033_, _05032_, _05020_);
  or (_05034_, _05033_, _04977_);
  and (_05035_, _05034_, _22768_);
  and (_05036_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_05037_, _05036_, _05005_);
  or (_05038_, _05037_, _05035_);
  and (_26869_[1], _05038_, _22762_);
  and (_05039_, _04832_, _23946_);
  and (_05041_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_23297_, _05041_, _05039_);
  and (_05042_, _01809_, _23991_);
  and (_05044_, _05042_, _23778_);
  not (_05045_, _05042_);
  and (_05047_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_23300_, _05047_, _05044_);
  and (_05049_, _24639_, _23649_);
  and (_05050_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_23319_, _05050_, _05049_);
  and (_05052_, _02326_, _23707_);
  and (_05053_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_23328_, _05053_, _05052_);
  and (_05054_, _25618_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_05055_, _26645_, _24618_);
  and (_05057_, _05055_, _24448_);
  or (_05058_, _05057_, _04945_);
  or (_05060_, _05058_, _02381_);
  or (_05061_, _24616_, _24584_);
  and (_05063_, _05061_, _26589_);
  or (_05064_, _05063_, _24537_);
  or (_05065_, _05064_, _26581_);
  or (_05066_, _05065_, _05060_);
  or (_05067_, _04942_, _03274_);
  or (_05068_, _05067_, _04984_);
  and (_05070_, _24606_, _24448_);
  and (_05072_, _00234_, _24445_);
  or (_05073_, _05072_, _05070_);
  or (_05074_, _03317_, _02380_);
  and (_05075_, _24596_, _24584_);
  and (_05077_, _24616_, _26587_);
  or (_05079_, _05077_, _05075_);
  and (_05080_, _26587_, _24545_);
  and (_05081_, _24594_, _24538_);
  or (_05083_, _05081_, _05080_);
  or (_05085_, _05083_, _05079_);
  or (_05086_, _05085_, _05074_);
  and (_05087_, _24618_, _24556_);
  and (_05088_, _26645_, _26582_);
  or (_05089_, _05088_, _05087_);
  and (_05090_, _00234_, _24448_);
  or (_05091_, _05090_, _26668_);
  or (_05093_, _05091_, _05089_);
  or (_05095_, _05093_, _05086_);
  or (_05096_, _05095_, _05073_);
  or (_05097_, _05096_, _05068_);
  or (_05098_, _05097_, _05066_);
  and (_05099_, _05098_, _25644_);
  or (_26870_[0], _05099_, _05054_);
  and (_05100_, _05008_, _23824_);
  and (_05101_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_27060_, _05101_, _05100_);
  and (_05102_, _01808_, _01758_);
  and (_05104_, _05102_, _23707_);
  not (_05105_, _05102_);
  and (_05107_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_23388_, _05107_, _05104_);
  and (_05109_, _05102_, _24050_);
  and (_05110_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_27302_, _05110_, _05109_);
  and (_05111_, _05102_, _23946_);
  and (_05113_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_23406_, _05113_, _05111_);
  and (_05114_, _24356_, _23656_);
  and (_05116_, _05114_, _23898_);
  not (_05117_, _05114_);
  and (_05118_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_23410_, _05118_, _05116_);
  and (_05119_, _24370_, _24005_);
  and (_05120_, _05119_, _23946_);
  not (_05121_, _05119_);
  and (_05122_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or (_23426_, _05122_, _05120_);
  and (_05125_, _24282_, _23754_);
  and (_05126_, _05125_, _24050_);
  not (_05127_, _05125_);
  and (_05128_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  or (_23477_, _05128_, _05126_);
  and (_05129_, _05008_, _23778_);
  and (_05130_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_23504_, _05130_, _05129_);
  and (_05131_, _05102_, _23778_);
  and (_05132_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_23507_, _05132_, _05131_);
  and (_05133_, _05102_, _23898_);
  and (_05134_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_23513_, _05134_, _05133_);
  and (_05135_, _05125_, _23707_);
  and (_05137_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  or (_23517_, _05137_, _05135_);
  and (_05138_, _24852_, _23898_);
  and (_05139_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  or (_23554_, _05139_, _05138_);
  and (_05140_, _05102_, _23747_);
  and (_05141_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_23566_, _05141_, _05140_);
  nand (_05142_, _24299_, _23702_);
  not (_05143_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_05144_, _04864_, _24313_);
  nor (_05145_, _05144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_05146_, _05145_, _05143_);
  and (_05147_, _05145_, _05143_);
  or (_05148_, _05147_, _05146_);
  and (_05149_, _05148_, _04861_);
  and (_05151_, _04876_, _24310_);
  and (_05152_, _05151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_05153_, _05152_, _05143_);
  and (_05154_, _05152_, _05143_);
  or (_05156_, _05154_, _05153_);
  and (_05157_, _05156_, _24302_);
  and (_05158_, _24309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_05159_, _05158_, _26114_);
  and (_05160_, _05159_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_05161_, _05160_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_05162_, _05161_, _26110_);
  or (_05163_, _05162_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_05164_, _05158_, _26115_);
  and (_05165_, _05164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_05166_, _05165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_05167_, _05166_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_05168_, _05167_, _26097_);
  and (_05169_, _05168_, _05163_);
  or (_05170_, _05169_, _05157_);
  or (_05171_, _05170_, _05149_);
  or (_05172_, _05171_, _24299_);
  and (_05173_, _05172_, _24294_);
  and (_05174_, _05173_, _05142_);
  and (_05175_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_05176_, _05175_, _05174_);
  and (_23573_, _05176_, _22762_);
  and (_05177_, _05125_, _23649_);
  and (_05178_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or (_23586_, _05178_, _05177_);
  and (_05180_, _01809_, _23903_);
  and (_05181_, _05180_, _23649_);
  not (_05182_, _05180_);
  and (_05183_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_23620_, _05183_, _05181_);
  and (_05184_, _05114_, _23707_);
  and (_05186_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_23650_, _05186_, _05184_);
  and (_05187_, _25078_, _24356_);
  and (_05188_, _05187_, _23824_);
  not (_05189_, _05187_);
  and (_05190_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_23659_, _05190_, _05188_);
  and (_05191_, _25142_, _23824_);
  and (_05192_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  or (_23685_, _05192_, _05191_);
  and (_05193_, _24201_, _23911_);
  not (_05194_, _05193_);
  and (_05195_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  and (_05197_, _05193_, _23707_);
  or (_23698_, _05197_, _05195_);
  and (_05199_, _24282_, _24201_);
  not (_05200_, _05199_);
  and (_05201_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  and (_05203_, _05199_, _23898_);
  or (_23703_, _05203_, _05201_);
  and (_05204_, _02321_, _23778_);
  and (_05205_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  or (_23723_, _05205_, _05204_);
  nor (_26912_, _02387_, rst);
  and (_05206_, _24063_, _23073_);
  and (_05207_, _05206_, _25171_);
  and (_05208_, _05207_, _25926_);
  nand (_05209_, _05208_, _23702_);
  or (_05210_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_05211_, _05210_, _22762_);
  and (_26874_[7], _05211_, _05209_);
  and (_05212_, _05206_, _26683_);
  not (_05213_, _05212_);
  nor (_05214_, _05213_, _23702_);
  not (_05215_, _25926_);
  and (_05216_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_05217_, _05216_, _05215_);
  or (_05218_, _05217_, _05214_);
  or (_05219_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_05221_, _05219_, _22762_);
  and (_26875_[7], _05221_, _05218_);
  and (_05222_, _05206_, _02310_);
  and (_05223_, _05222_, _25926_);
  nand (_05224_, _05223_, _23702_);
  or (_05226_, _05223_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_05227_, _05226_, _22762_);
  and (_26876_[7], _05227_, _05224_);
  and (_05228_, _05206_, _24076_);
  and (_05229_, _05228_, _25926_);
  not (_05230_, _05229_);
  nor (_05231_, _05230_, _23702_);
  and (_05233_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_05234_, _05233_, _05231_);
  and (_26877_[7], _05234_, _22762_);
  and (_05235_, _02311_, _25171_);
  and (_05236_, _05235_, _25926_);
  and (_05237_, _05236_, _26750_);
  or (_05238_, _05222_, _05228_);
  or (_05239_, _05235_, _05238_);
  nor (_05240_, _05239_, _05212_);
  or (_05241_, _05240_, _05215_);
  or (_05242_, _05238_, _05212_);
  and (_05243_, _05242_, _25926_);
  or (_05244_, _05243_, _05241_);
  and (_05245_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or (_05246_, _05245_, _05237_);
  and (_26878_[7], _05246_, _22762_);
  and (_05247_, _02311_, _26683_);
  nor (_05248_, _05247_, _05235_);
  not (_05249_, _05248_);
  nor (_05250_, _05249_, _05238_);
  or (_05251_, _05250_, _05215_);
  or (_05252_, _05251_, _05239_);
  and (_05253_, _05252_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_05254_, _05247_, _25926_);
  not (_05255_, _05254_);
  nor (_05256_, _05255_, _23702_);
  or (_05257_, _05256_, _05253_);
  and (_26879_[7], _05257_, _22762_);
  nor (_05259_, _02315_, _23702_);
  and (_05260_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or (_05261_, _05260_, _05259_);
  and (_26880_[7], _05261_, _22762_);
  and (_05262_, _02311_, _24076_);
  and (_05263_, _05262_, _25926_);
  and (_05264_, _05263_, _26750_);
  nor (_05265_, _05262_, _02312_);
  and (_05266_, _05265_, _05248_);
  or (_05267_, _05266_, _05215_);
  not (_05268_, _02312_);
  nand (_05269_, _05248_, _05268_);
  and (_05270_, _05269_, _25926_);
  or (_05271_, _05270_, _05267_);
  and (_05272_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_05273_, _05272_, _05264_);
  and (_26881_[7], _05273_, _22762_);
  or (_05275_, _05223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  not (_05276_, _05223_);
  or (_05277_, _05276_, _23816_);
  and (_23763_, _05277_, _05275_);
  and (_05278_, _05223_, _23898_);
  and (_05279_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_23815_, _05279_, _05278_);
  and (_05281_, _23986_, _23754_);
  and (_05282_, _05281_, _23747_);
  not (_05283_, _05281_);
  and (_05284_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_23819_, _05284_, _05282_);
  and (_05285_, _05223_, _23778_);
  and (_05286_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_23826_, _05286_, _05285_);
  and (_05288_, _23911_, _23754_);
  and (_05289_, _05288_, _23649_);
  not (_05290_, _05288_);
  and (_05291_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  or (_23891_, _05291_, _05289_);
  and (_05292_, _05223_, _23946_);
  and (_05293_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_27278_, _05293_, _05292_);
  and (_05294_, _05223_, _23649_);
  and (_05295_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_23928_, _05295_, _05294_);
  and (_05296_, _05223_, _23747_);
  and (_05297_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_23931_, _05297_, _05296_);
  and (_05298_, _01758_, _23752_);
  and (_05299_, _05298_, _23824_);
  not (_05301_, _05298_);
  and (_05302_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_23996_, _05302_, _05299_);
  and (_05303_, _05298_, _23649_);
  and (_05304_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_23999_, _05304_, _05303_);
  and (_05305_, _05298_, _23747_);
  and (_05307_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_24002_, _05307_, _05305_);
  nor (_26897_[5], _00727_, rst);
  and (_05308_, _05288_, _23898_);
  and (_05309_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or (_24091_, _05309_, _05308_);
  and (_05310_, _05298_, _23707_);
  and (_05311_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_24097_, _05311_, _05310_);
  and (_05313_, _05298_, _24050_);
  and (_05314_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_24099_, _05314_, _05313_);
  and (_05315_, _05288_, _23707_);
  and (_05316_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or (_24106_, _05316_, _05315_);
  and (_05317_, _05288_, _24050_);
  and (_05318_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or (_27057_, _05318_, _05317_);
  and (_05319_, _01758_, _23656_);
  and (_05320_, _05319_, _23747_);
  not (_05322_, _05319_);
  and (_05323_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_24133_, _05323_, _05320_);
  and (_05324_, _05319_, _23946_);
  and (_05325_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_27234_, _05325_, _05324_);
  and (_05326_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  and (_05327_, _05199_, _23778_);
  or (_27230_, _05327_, _05326_);
  and (_05328_, _05319_, _23649_);
  and (_05329_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_24183_, _05329_, _05328_);
  and (_05330_, _05125_, _23778_);
  and (_05331_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  or (_24200_, _05331_, _05330_);
  and (_05332_, _05319_, _23707_);
  and (_05333_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_24202_, _05333_, _05332_);
  and (_05334_, _05298_, _23778_);
  and (_05335_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_24205_, _05335_, _05334_);
  and (_05336_, _23785_, _23662_);
  and (_05337_, _05336_, _24085_);
  not (_05338_, _05337_);
  and (_05339_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  and (_05340_, _05337_, _23649_);
  or (_24227_, _05340_, _05339_);
  and (_05342_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  and (_05343_, _05337_, _23747_);
  or (_24233_, _05343_, _05342_);
  and (_05344_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  and (_05345_, _05337_, _23824_);
  or (_24278_, _05345_, _05344_);
  and (_05346_, _01758_, _25078_);
  and (_05347_, _05346_, _24050_);
  not (_05348_, _05346_);
  and (_05349_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_24281_, _05349_, _05347_);
  and (_05350_, _01808_, _23754_);
  and (_05351_, _05350_, _23707_);
  not (_05352_, _05350_);
  and (_05353_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  or (_24298_, _05353_, _05351_);
  and (_05354_, _05336_, _24010_);
  not (_05355_, _05354_);
  and (_05356_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  and (_05357_, _05354_, _23778_);
  or (_24306_, _05357_, _05356_);
  and (_05358_, _05336_, _24275_);
  not (_05359_, _05358_);
  and (_05360_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  and (_05361_, _05358_, _23898_);
  or (_27105_, _05361_, _05360_);
  and (_05362_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  and (_05363_, _05358_, _24050_);
  or (_24311_, _05363_, _05362_);
  and (_05364_, _05319_, _23898_);
  and (_05365_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_24314_, _05365_, _05364_);
  and (_05366_, _05319_, _23778_);
  and (_05367_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_24321_, _05367_, _05366_);
  and (_05368_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  and (_05369_, _05358_, _23707_);
  or (_24327_, _05369_, _05368_);
  and (_05371_, _01809_, _23784_);
  and (_05372_, _05371_, _23778_);
  not (_05373_, _05371_);
  and (_05374_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_24330_, _05374_, _05372_);
  and (_05375_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  and (_05376_, _05337_, _23707_);
  or (_24355_, _05376_, _05375_);
  and (_05377_, _04797_, _23747_);
  and (_05378_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_24357_, _05378_, _05377_);
  and (_05379_, _01758_, _24282_);
  and (_05380_, _05379_, _23707_);
  not (_05381_, _05379_);
  and (_05382_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_24387_, _05382_, _05380_);
  and (_05384_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  and (_05385_, _05337_, _24050_);
  or (_24390_, _05385_, _05384_);
  and (_05387_, _05379_, _24050_);
  and (_05388_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_27204_, _05388_, _05387_);
  and (_05390_, _05379_, _23946_);
  and (_05391_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_24395_, _05391_, _05390_);
  and (_05392_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  and (_05393_, _05337_, _23946_);
  or (_24398_, _05393_, _05392_);
  and (_05394_, _05346_, _23747_);
  and (_05395_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_24410_, _05395_, _05394_);
  and (_05396_, _05346_, _23824_);
  and (_05397_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_24413_, _05397_, _05396_);
  and (_05398_, _05336_, _23784_);
  not (_05399_, _05398_);
  and (_05400_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_05401_, _05398_, _23649_);
  or (_24416_, _05401_, _05400_);
  and (_05402_, _05346_, _23898_);
  and (_05403_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_24419_, _05403_, _05402_);
  and (_05404_, _05346_, _23778_);
  and (_05405_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_24423_, _05405_, _05404_);
  and (_05407_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_05409_, _05398_, _23946_);
  or (_24433_, _05409_, _05407_);
  and (_05410_, _01808_, _23076_);
  and (_05411_, _05410_, _23649_);
  not (_05412_, _05410_);
  and (_05413_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  or (_24449_, _05413_, _05411_);
  and (_05414_, _05379_, _23778_);
  and (_05415_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_27203_, _05415_, _05414_);
  and (_05416_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_05417_, _05398_, _23707_);
  or (_24465_, _05417_, _05416_);
  and (_05419_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  and (_05420_, _05337_, _23778_);
  or (_24468_, _05420_, _05419_);
  and (_05422_, _05379_, _23747_);
  and (_05424_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_24496_, _05424_, _05422_);
  and (_05425_, _05379_, _23824_);
  and (_05426_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_24499_, _05426_, _05425_);
  and (_05427_, _05379_, _23898_);
  and (_05428_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_24502_, _05428_, _05427_);
  and (_05429_, _01758_, _23911_);
  and (_05430_, _05429_, _23824_);
  not (_05431_, _05429_);
  and (_05432_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_24547_, _05432_, _05430_);
  and (_05433_, _05429_, _23649_);
  and (_05434_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_24551_, _05434_, _05433_);
  and (_05435_, _05429_, _23747_);
  and (_05436_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_24557_, _05436_, _05435_);
  and (_05437_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  and (_05438_, _05358_, _23946_);
  or (_24571_, _05438_, _05437_);
  and (_05439_, _05371_, _23898_);
  and (_05440_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_24580_, _05440_, _05439_);
  and (_05441_, _05371_, _23747_);
  and (_05442_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_24583_, _05442_, _05441_);
  and (_05443_, _05429_, _24050_);
  and (_05444_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_24590_, _05444_, _05443_);
  and (_05445_, _01809_, _24085_);
  and (_05446_, _05445_, _23778_);
  not (_05447_, _05445_);
  and (_05448_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  or (_27106_, _05448_, _05446_);
  and (_05449_, _05371_, _24050_);
  and (_05450_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_24603_, _05450_, _05449_);
  and (_05452_, _05371_, _23707_);
  and (_05453_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_24609_, _05453_, _05452_);
  and (_05454_, _01758_, _24010_);
  and (_05455_, _05454_, _24050_);
  not (_05457_, _05454_);
  and (_05458_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_24638_, _05458_, _05455_);
  not (_05459_, _05208_);
  and (_05460_, _05459_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_05461_, _05208_, _24685_);
  or (_05462_, _05461_, _05460_);
  and (_26874_[0], _05462_, _22762_);
  or (_05463_, _05459_, _23892_);
  or (_05464_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_05466_, _05464_, _22762_);
  and (_26874_[1], _05466_, _05463_);
  or (_05467_, _05459_, _23816_);
  or (_05468_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_05469_, _05468_, _22762_);
  and (_26874_[2], _05469_, _05467_);
  or (_05470_, _05459_, _23738_);
  or (_05471_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_05472_, _05471_, _22762_);
  and (_26874_[3], _05472_, _05470_);
  or (_05474_, _05459_, _23642_);
  or (_05475_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_05477_, _05475_, _22762_);
  and (_26874_[4], _05477_, _05474_);
  or (_05478_, _05459_, _23939_);
  or (_05480_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_05481_, _05480_, _22762_);
  and (_26874_[5], _05481_, _05478_);
  or (_05482_, _05459_, _24043_);
  or (_05483_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_05484_, _05483_, _22762_);
  and (_26874_[6], _05484_, _05482_);
  nor (_05485_, _05215_, _23772_);
  and (_05486_, _05485_, _05212_);
  nand (_05487_, _05212_, _25926_);
  and (_05488_, _05487_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_05489_, _05488_, _05486_);
  and (_26875_[0], _05489_, _22762_);
  and (_05490_, _05212_, _23892_);
  and (_05491_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_05492_, _05491_, _05215_);
  or (_05493_, _05492_, _05490_);
  or (_05494_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_05495_, _05494_, _22762_);
  and (_26875_[1], _05495_, _05493_);
  and (_05496_, _05212_, _23816_);
  and (_05497_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_05499_, _05497_, _05215_);
  or (_05500_, _05499_, _05496_);
  or (_05501_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_05502_, _05501_, _22762_);
  and (_26875_[2], _05502_, _05500_);
  and (_05504_, _05212_, _23738_);
  and (_05505_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_05506_, _05505_, _05215_);
  or (_05507_, _05506_, _05504_);
  or (_05508_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_05509_, _05508_, _22762_);
  and (_26875_[3], _05509_, _05507_);
  and (_05510_, _05212_, _23642_);
  and (_05511_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_05512_, _05511_, _05215_);
  or (_05513_, _05512_, _05510_);
  or (_05514_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_05515_, _05514_, _22762_);
  and (_26875_[4], _05515_, _05513_);
  and (_05516_, _05212_, _23939_);
  and (_05517_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_05518_, _05517_, _05215_);
  or (_05519_, _05518_, _05516_);
  or (_05520_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_05521_, _05520_, _22762_);
  and (_26875_[5], _05521_, _05519_);
  and (_05522_, _05212_, _24043_);
  and (_05523_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_05524_, _05523_, _05215_);
  or (_05525_, _05524_, _05522_);
  or (_05526_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_05527_, _05526_, _22762_);
  and (_26875_[6], _05527_, _05525_);
  not (_05528_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_05529_, _05212_, _05207_);
  not (_05530_, _05222_);
  and (_05531_, _05530_, _05529_);
  nor (_05532_, _05531_, _05215_);
  nor (_05533_, _05532_, _05528_);
  nand (_05534_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_05535_, _05534_, _05529_);
  and (_05536_, _05223_, _24685_);
  or (_05537_, _05536_, _05535_);
  or (_05538_, _05537_, _05533_);
  and (_26876_[0], _05538_, _22762_);
  and (_05539_, _05223_, _23892_);
  and (_05540_, _05276_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_05541_, _05540_, _05539_);
  and (_26876_[1], _05541_, _22762_);
  or (_05544_, _05223_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_05545_, _05544_, _22762_);
  and (_26876_[2], _05545_, _05277_);
  or (_05547_, _05276_, _23738_);
  or (_05548_, _05223_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_05550_, _05548_, _22762_);
  and (_26876_[3], _05550_, _05547_);
  or (_05551_, _05276_, _23642_);
  or (_05552_, _05223_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_05553_, _05552_, _22762_);
  and (_26876_[4], _05553_, _05551_);
  and (_05554_, _05223_, _23939_);
  and (_05555_, _05276_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_05556_, _05555_, _05554_);
  and (_26876_[5], _05556_, _22762_);
  and (_05558_, _05223_, _24043_);
  and (_05559_, _05276_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_05560_, _05559_, _05558_);
  and (_26876_[6], _05560_, _22762_);
  and (_05561_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_05562_, _05485_, _05228_);
  or (_05563_, _05562_, _05561_);
  and (_26877_[0], _05563_, _22762_);
  and (_05564_, _05229_, _23892_);
  or (_05565_, _05230_, _05532_);
  and (_05566_, _05565_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_05567_, _05566_, _05564_);
  and (_26877_[1], _05567_, _22762_);
  and (_05569_, _05229_, _23816_);
  and (_05571_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_05572_, _05571_, _05569_);
  and (_26877_[2], _05572_, _22762_);
  and (_05574_, _05229_, _23738_);
  and (_05575_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_05576_, _05575_, _05574_);
  and (_26877_[3], _05576_, _22762_);
  and (_05578_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_05579_, _05229_, _23642_);
  or (_05580_, _05579_, _05578_);
  and (_26877_[4], _05580_, _22762_);
  and (_05581_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_05582_, _05229_, _23939_);
  or (_05583_, _05582_, _05581_);
  and (_26877_[5], _05583_, _22762_);
  and (_05585_, _05229_, _24043_);
  and (_05586_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_05588_, _05586_, _05585_);
  and (_26877_[6], _05588_, _22762_);
  and (_05590_, _05454_, _23946_);
  and (_05591_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_27172_, _05591_, _05590_);
  or (_05592_, _05242_, _05241_);
  and (_05593_, _05592_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_05594_, _05485_, _05235_);
  or (_05595_, _05594_, _05593_);
  and (_26878_[0], _05595_, _22762_);
  and (_05596_, _05236_, _23892_);
  and (_05597_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  or (_05599_, _05597_, _05596_);
  and (_26878_[1], _05599_, _22762_);
  and (_05600_, _05236_, _23816_);
  and (_05601_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or (_05602_, _05601_, _05600_);
  and (_26878_[2], _05602_, _22762_);
  and (_05603_, _05236_, _23738_);
  and (_05604_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or (_05605_, _05604_, _05603_);
  and (_26878_[3], _05605_, _22762_);
  and (_05606_, _05592_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_05607_, _05236_, _23642_);
  or (_05608_, _05607_, _05606_);
  and (_26878_[4], _05608_, _22762_);
  and (_05609_, _05236_, _23939_);
  and (_05610_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_05611_, _05610_, _05609_);
  and (_26878_[5], _05611_, _22762_);
  and (_05612_, _05236_, _24043_);
  and (_05613_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or (_05614_, _05613_, _05612_);
  and (_26878_[6], _05614_, _22762_);
  and (_05615_, _05252_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_05616_, _05485_, _05247_);
  or (_05617_, _05616_, _05615_);
  and (_26879_[0], _05617_, _22762_);
  and (_05618_, _05251_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_05619_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_05620_, _05619_, _05239_);
  and (_05621_, _05254_, _23892_);
  or (_05623_, _05621_, _05620_);
  or (_05624_, _05623_, _05618_);
  and (_26879_[1], _05624_, _22762_);
  and (_05626_, _05254_, _23816_);
  and (_05627_, _05255_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or (_05628_, _05627_, _05626_);
  and (_26879_[2], _05628_, _22762_);
  and (_05629_, _05254_, _23738_);
  and (_05630_, _05251_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_05631_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_05632_, _05631_, _05239_);
  or (_05634_, _05632_, _05630_);
  or (_05635_, _05634_, _05629_);
  and (_26879_[3], _05635_, _22762_);
  and (_05636_, _05254_, _23642_);
  and (_05637_, _05252_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or (_05638_, _05637_, _05636_);
  and (_26879_[4], _05638_, _22762_);
  and (_05640_, _05255_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_05641_, _05254_, _23939_);
  or (_05642_, _05641_, _05640_);
  and (_26879_[5], _05642_, _22762_);
  and (_05644_, _05254_, _24043_);
  and (_05645_, _05252_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or (_05646_, _05645_, _05644_);
  and (_26879_[6], _05646_, _22762_);
  and (_05647_, _05454_, _23649_);
  and (_05648_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_24681_, _05648_, _05647_);
  and (_05649_, _05485_, _02312_);
  and (_05650_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or (_05651_, _05650_, _05649_);
  and (_26880_[0], _05651_, _22762_);
  and (_05652_, _02313_, _23892_);
  and (_05653_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  or (_05654_, _05653_, _05652_);
  and (_26880_[1], _05654_, _22762_);
  and (_05655_, _02313_, _23816_);
  and (_05656_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or (_05657_, _05656_, _05655_);
  and (_26880_[2], _05657_, _22762_);
  and (_05658_, _02313_, _23738_);
  and (_05660_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or (_05662_, _05660_, _05658_);
  and (_26880_[3], _05662_, _22762_);
  and (_05663_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_05664_, _02313_, _23642_);
  or (_05665_, _05664_, _05663_);
  and (_26880_[4], _05665_, _22762_);
  and (_05666_, _02313_, _23939_);
  and (_05667_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_05668_, _05667_, _05666_);
  and (_26880_[5], _05668_, _22762_);
  and (_05669_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_05670_, _05669_, _02314_);
  and (_26880_[6], _05670_, _22762_);
  and (_05671_, _05485_, _05262_);
  and (_05672_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or (_05674_, _05672_, _05671_);
  and (_26881_[0], _05674_, _22762_);
  and (_05675_, _05263_, _23892_);
  and (_05676_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  or (_05677_, _05676_, _05675_);
  and (_26881_[1], _05677_, _22762_);
  and (_05679_, _05263_, _23816_);
  or (_05680_, _05267_, _05269_);
  and (_05681_, _05680_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_05682_, _05681_, _05679_);
  and (_26881_[2], _05682_, _22762_);
  and (_05683_, _05263_, _23738_);
  and (_05684_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or (_05685_, _05684_, _05683_);
  and (_26881_[3], _05685_, _22762_);
  and (_05686_, _05263_, _23642_);
  and (_05687_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_05688_, _05687_, _05686_);
  and (_26881_[4], _05688_, _22762_);
  and (_05690_, _05680_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_05691_, _05263_, _23939_);
  or (_05692_, _05691_, _05690_);
  and (_26881_[5], _05692_, _22762_);
  and (_05693_, _05263_, _24043_);
  and (_05694_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or (_05695_, _05694_, _05693_);
  and (_26881_[6], _05695_, _22762_);
  and (_05696_, _05410_, _23747_);
  and (_05697_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or (_24697_, _05697_, _05696_);
  and (_05698_, _25142_, _23898_);
  and (_05699_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or (_27200_, _05699_, _05698_);
  and (_05701_, _23991_, _23664_);
  and (_05702_, _05701_, _23898_);
  not (_05703_, _05701_);
  and (_05704_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_25107_, _05704_, _05702_);
  and (_05705_, _05336_, _23911_);
  not (_05706_, _05705_);
  and (_05708_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and (_05709_, _05705_, _23649_);
  or (_25124_, _05709_, _05708_);
  and (_05710_, _02325_, _23991_);
  and (_05711_, _05710_, _23649_);
  not (_05712_, _05710_);
  and (_05713_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  or (_27162_, _05713_, _05711_);
  and (_05714_, _02325_, _23903_);
  and (_05715_, _05714_, _23946_);
  not (_05716_, _05714_);
  and (_05717_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  or (_25147_, _05717_, _05715_);
  and (_05718_, _05701_, _23778_);
  and (_05719_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_25149_, _05719_, _05718_);
  and (_05720_, _05714_, _23778_);
  and (_05721_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  or (_25152_, _05721_, _05720_);
  and (_05722_, _04917_, _23946_);
  and (_05723_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_25177_, _05723_, _05722_);
  and (_05724_, _04917_, _23747_);
  and (_05725_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_25180_, _05725_, _05724_);
  not (_05726_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_05727_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and (_05728_, _05727_, _05726_);
  and (_05729_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _22762_);
  and (_27303_, _05729_, _05728_);
  nor (_05730_, _05728_, rst);
  nand (_05731_, _05727_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_05732_, _05727_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_05733_, _05732_, _05731_);
  and (_27304_[3], _05733_, _05730_);
  not (_05734_, _00014_);
  nor (_05735_, _05734_, _26817_);
  and (_05736_, _02397_, _26777_);
  and (_05737_, _05736_, _00037_);
  and (_05738_, _05737_, _05735_);
  not (_05739_, _00263_);
  nand (_05740_, _00451_, _05739_);
  and (_05741_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_05742_, _00267_, _00264_);
  not (_05743_, _05742_);
  nor (_05744_, _24291_, _23304_);
  nor (_05745_, _05744_, _04389_);
  nor (_05746_, _05745_, _05743_);
  nor (_05747_, _05746_, _05741_);
  nand (_05748_, _05747_, _05740_);
  nand (_05749_, _05748_, _00257_);
  nor (_05750_, _01061_, _00257_);
  not (_05751_, _05750_);
  nand (_05752_, _05751_, _05749_);
  nand (_05753_, _00545_, _05739_);
  and (_05755_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand (_05756_, _24118_, _23594_);
  or (_05757_, _24118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_05758_, _05757_, _05742_);
  and (_05759_, _05758_, _05756_);
  nor (_05760_, _05759_, _05755_);
  and (_05761_, _05760_, _00257_);
  and (_05762_, _05761_, _05753_);
  and (_05763_, _01129_, _00256_);
  nor (_05764_, _05763_, _05762_);
  nand (_05765_, _05764_, _05752_);
  or (_05766_, _05764_, _05752_);
  nand (_05767_, _05766_, _05765_);
  nand (_05768_, _26565_, _05739_);
  nor (_05770_, _24678_, _23387_);
  nor (_05771_, _05770_, _04418_);
  nor (_05772_, _05771_, _05743_);
  and (_05773_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_05774_, _05773_, _00256_);
  nor (_05775_, _05774_, _05772_);
  nand (_05776_, _05775_, _05768_);
  or (_05777_, _00930_, _00257_);
  and (_05778_, _05777_, _05776_);
  or (_05779_, _00372_, _00263_);
  nor (_05780_, _24067_, _23355_);
  nor (_05781_, _05780_, _04398_);
  nor (_05782_, _05781_, _05743_);
  and (_05783_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_05785_, _05783_, _00256_);
  nor (_05786_, _05785_, _05782_);
  nand (_05787_, _05786_, _05779_);
  and (_05789_, _00993_, _00256_);
  not (_05790_, _05789_);
  nand (_05791_, _05790_, _05787_);
  nand (_05792_, _05791_, _05778_);
  or (_05793_, _05791_, _05778_);
  nand (_05794_, _05793_, _05792_);
  nand (_05795_, _05794_, _05767_);
  or (_05796_, _05794_, _05767_);
  nand (_05797_, _05796_, _05795_);
  and (_05798_, _00620_, _05739_);
  nor (_05799_, _24296_, _23239_);
  or (_05800_, _05799_, _24745_);
  and (_05801_, _05800_, _05742_);
  and (_05802_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_05803_, _05802_, _00256_);
  or (_05805_, _05803_, _05801_);
  or (_05806_, _05805_, _05798_);
  or (_05807_, _01192_, _00257_);
  and (_05808_, _05807_, _05806_);
  and (_05809_, _00708_, _05739_);
  nand (_05810_, _24125_, _23594_);
  or (_05811_, _24125_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_05812_, _05811_, _05742_);
  and (_05813_, _05812_, _05810_);
  and (_05814_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_05816_, _05814_, _00256_);
  or (_05817_, _05816_, _05813_);
  or (_05818_, _05817_, _05809_);
  or (_05819_, _01255_, _00257_);
  and (_05820_, _05819_, _05818_);
  or (_05821_, _05820_, _05808_);
  nand (_05822_, _05820_, _05808_);
  nand (_05823_, _05822_, _05821_);
  or (_05824_, _00793_, _00263_);
  not (_05826_, _24705_);
  nor (_05827_, _05826_, _23594_);
  nor (_05828_, _24705_, _23166_);
  nor (_05829_, _05828_, _05827_);
  nor (_05830_, _05829_, _05743_);
  and (_05831_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_05832_, _05831_, _00256_);
  nor (_05833_, _05832_, _05830_);
  and (_05834_, _05833_, _05824_);
  and (_05835_, _01318_, _00256_);
  or (_05836_, _05835_, _05834_);
  and (_05837_, _00875_, _05739_);
  not (_05838_, _24654_);
  nor (_05839_, _05838_, _23594_);
  nor (_05840_, _24654_, _23126_);
  or (_05841_, _05840_, _05839_);
  and (_05843_, _05841_, _05742_);
  and (_05844_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_05845_, _05844_, _00256_);
  or (_05846_, _05845_, _05843_);
  or (_05847_, _05846_, _05837_);
  or (_05848_, _04299_, _00257_);
  and (_05850_, _05848_, _05847_);
  or (_05851_, _05850_, _05836_);
  nand (_05852_, _05850_, _05836_);
  and (_05853_, _05852_, _05851_);
  nand (_05855_, _05853_, _05823_);
  or (_05856_, _05853_, _05823_);
  nand (_05857_, _05856_, _05855_);
  nand (_05858_, _05857_, _05797_);
  or (_05859_, _05857_, _05797_);
  and (_05860_, _05859_, _05858_);
  nand (_05861_, _05860_, _00168_);
  and (_05863_, _00134_, _00099_);
  or (_05864_, _00168_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_05865_, _05864_, _05863_);
  and (_05866_, _05865_, _05861_);
  not (_05867_, _00134_);
  nor (_05868_, _05867_, _00099_);
  nor (_05869_, _00168_, _00527_);
  and (_05870_, _00168_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_05871_, _05870_, _05869_);
  and (_05872_, _05871_, _05868_);
  or (_05873_, _00168_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_05874_, _00134_, _00099_);
  not (_05876_, _00168_);
  or (_05877_, _05876_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_05878_, _05877_, _05874_);
  and (_05879_, _05878_, _05873_);
  or (_05880_, _00168_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_05881_, _05867_, _00099_);
  or (_05882_, _05876_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_05883_, _05882_, _05881_);
  and (_05884_, _05883_, _05880_);
  or (_05885_, _05884_, _05879_);
  or (_05886_, _05885_, _05872_);
  or (_05887_, _05886_, _05866_);
  and (_05888_, _05887_, _05738_);
  and (_05889_, _00175_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not (_05890_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_05891_, _00037_);
  and (_05892_, _00058_, _26777_);
  and (_05893_, _05892_, _05891_);
  and (_05894_, _05893_, _05735_);
  nor (_05895_, _05894_, _05890_);
  and (_05896_, _05892_, _00037_);
  not (_05897_, _05896_);
  nor (_05898_, _05897_, _05735_);
  and (_05900_, _26817_, _26777_);
  and (_05901_, _05900_, _05891_);
  or (_05903_, _05901_, _05737_);
  nor (_05904_, _05903_, _05898_);
  and (_05906_, _05904_, _05895_);
  nor (_05908_, _00014_, _26817_);
  and (_05909_, _05908_, _05737_);
  and (_05910_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_05911_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_05912_, _05911_, _05910_);
  and (_05913_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_05914_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_05916_, _05914_, _05913_);
  or (_05917_, _05916_, _05912_);
  and (_05918_, _05917_, _05876_);
  and (_05919_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_05920_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_05921_, _05920_, _05919_);
  and (_05922_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_05923_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_05924_, _05923_, _05922_);
  or (_05925_, _05924_, _05921_);
  and (_05926_, _05925_, _00168_);
  or (_05927_, _05926_, _05918_);
  and (_05928_, _05927_, _05909_);
  and (_05929_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_05930_, _05929_, _05876_);
  and (_05931_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_05932_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_05933_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_05934_, _05933_, _05932_);
  or (_05935_, _05934_, _05931_);
  or (_05936_, _05935_, _05930_);
  nor (_05937_, _00058_, _00014_);
  and (_05938_, _05937_, _05936_);
  and (_05939_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_05940_, _05939_, _00168_);
  and (_05941_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_05942_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_05943_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_05944_, _05943_, _05942_);
  or (_05945_, _05944_, _05941_);
  or (_05946_, _05945_, _05940_);
  and (_05947_, _05946_, _05901_);
  and (_05948_, _05947_, _05938_);
  or (_05950_, _05948_, _05928_);
  or (_05951_, _05950_, _05906_);
  or (_05952_, _05951_, _05889_);
  and (_05953_, _05734_, _26817_);
  and (_05954_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_05955_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_05957_, _05955_, _05954_);
  and (_05958_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_05959_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_05960_, _05959_, _05958_);
  or (_05961_, _05960_, _05957_);
  and (_05962_, _05961_, _05953_);
  and (_05963_, _00014_, _26817_);
  and (_05965_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_05966_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_05967_, _05966_, _05965_);
  and (_05969_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_05970_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_05972_, _05970_, _05969_);
  or (_05973_, _05972_, _05967_);
  and (_05975_, _05973_, _05963_);
  or (_05976_, _05975_, _05962_);
  and (_05977_, _05976_, _00168_);
  and (_05978_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_05979_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_05980_, _05979_, _05978_);
  and (_05981_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_05982_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_05983_, _05982_, _05981_);
  or (_05984_, _05983_, _05980_);
  and (_05985_, _05984_, _05963_);
  and (_05986_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_05988_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_05989_, _05988_, _05986_);
  and (_05990_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_05992_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_05993_, _05992_, _05990_);
  or (_05994_, _05993_, _05989_);
  and (_05996_, _05994_, _05953_);
  or (_05997_, _05996_, _05985_);
  and (_05998_, _05997_, _05876_);
  or (_05999_, _05998_, _05977_);
  and (_06000_, _05999_, _05893_);
  and (_06001_, _02397_, _00014_);
  and (_06002_, _06001_, _05901_);
  and (_06003_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_06004_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_06005_, _06004_, _06003_);
  and (_06006_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_06007_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_06008_, _06007_, _06006_);
  or (_06010_, _06008_, _06005_);
  and (_06011_, _06010_, _00168_);
  and (_06012_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_06013_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_06014_, _06013_, _06012_);
  and (_06015_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_06017_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_06018_, _06017_, _06015_);
  or (_06019_, _06018_, _06014_);
  and (_06020_, _06019_, _05876_);
  or (_06021_, _06020_, _06011_);
  and (_06022_, _06021_, _06002_);
  and (_06024_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_06025_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_06026_, _06025_, _06024_);
  and (_06027_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_06028_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_06029_, _06028_, _06027_);
  or (_06030_, _06029_, _06026_);
  and (_06032_, _06030_, _05876_);
  and (_06033_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_06034_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_06035_, _06034_, _06033_);
  and (_06036_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_06037_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_06038_, _06037_, _06036_);
  or (_06039_, _06038_, _06035_);
  and (_06040_, _06039_, _00168_);
  or (_06042_, _06040_, _06032_);
  and (_06043_, _06042_, _05894_);
  or (_06044_, _06043_, _06022_);
  and (_06045_, _05908_, _05896_);
  and (_06046_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_06047_, _06046_, _05876_);
  and (_06048_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_06049_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_06050_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_06052_, _06050_, _06049_);
  or (_06053_, _06052_, _06048_);
  or (_06054_, _06053_, _06047_);
  and (_06055_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_06056_, _06055_, _00168_);
  and (_06057_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_06058_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_06059_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_06060_, _06059_, _06058_);
  or (_06061_, _06060_, _06057_);
  or (_06062_, _06061_, _06056_);
  and (_06063_, _06062_, _06054_);
  and (_06064_, _06063_, _06045_);
  or (_06065_, _06064_, _06044_);
  or (_06066_, _06065_, _06000_);
  or (_06067_, _06066_, _05952_);
  or (_06068_, _04982_, _26662_);
  or (_06069_, _02254_, _26663_);
  or (_06070_, _06069_, _24591_);
  and (_06071_, _26625_, _24588_);
  or (_06072_, _06071_, _04978_);
  and (_06073_, _26625_, _24616_);
  or (_06074_, _06073_, _02262_);
  or (_06075_, _06074_, _06072_);
  or (_06076_, _06075_, _26615_);
  or (_06078_, _06076_, _06070_);
  or (_06079_, _26620_, _24617_);
  and (_06080_, _24618_, _24613_);
  or (_06081_, _05063_, _06080_);
  or (_06082_, _06081_, _06079_);
  or (_06083_, _06082_, _06078_);
  or (_06084_, _06083_, _06068_);
  or (_06086_, _06084_, _26659_);
  and (_06087_, _06086_, _26572_);
  or (_06089_, _06087_, p2_in[1]);
  not (_06090_, _06087_);
  or (_06091_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_06092_, _06091_, _06089_);
  and (_06094_, _06092_, _05881_);
  nor (_06095_, _06087_, p2_in[0]);
  and (_06096_, _06087_, _25336_);
  nor (_06097_, _06096_, _06095_);
  and (_06099_, _06097_, _05863_);
  or (_06101_, _06099_, _06094_);
  or (_06102_, _06087_, p2_in[2]);
  or (_06104_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_06105_, _06104_, _06102_);
  and (_06106_, _06105_, _05868_);
  or (_06107_, _06087_, p2_in[3]);
  or (_06108_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_06110_, _06108_, _06107_);
  and (_06111_, _06110_, _05874_);
  or (_06113_, _06111_, _06106_);
  or (_06114_, _06113_, _06101_);
  and (_06115_, _06114_, _05896_);
  or (_06117_, _06087_, p3_in[3]);
  or (_06118_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_06119_, _06118_, _06117_);
  and (_06120_, _06119_, _05874_);
  or (_06122_, _06087_, p3_in[1]);
  or (_06124_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_06125_, _06124_, _06122_);
  and (_06126_, _06125_, _05881_);
  or (_06127_, _06126_, _06120_);
  or (_06128_, _06087_, p3_in[2]);
  or (_06129_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_06130_, _06129_, _06128_);
  and (_06132_, _06130_, _05868_);
  nor (_06133_, _06087_, p3_in[0]);
  and (_06135_, _06087_, _25217_);
  nor (_06136_, _06135_, _06133_);
  and (_06137_, _06136_, _05863_);
  or (_06138_, _06137_, _06132_);
  or (_06139_, _06138_, _06127_);
  and (_06140_, _06139_, _05737_);
  or (_06142_, _06140_, _06115_);
  and (_06143_, _06142_, _00168_);
  nor (_06144_, _06087_, p3_in[6]);
  and (_06145_, _06087_, _25234_);
  nor (_06146_, _06145_, _06144_);
  and (_06147_, _06146_, _05868_);
  nor (_06148_, _06087_, p3_in[4]);
  not (_06149_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_06150_, _06087_, _06149_);
  nor (_06152_, _06150_, _06148_);
  and (_06153_, _06152_, _05863_);
  or (_06154_, _06153_, _06147_);
  or (_06155_, _06087_, p3_in[7]);
  or (_06156_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_06157_, _06156_, _06155_);
  and (_06158_, _06157_, _05874_);
  or (_06159_, _06087_, p3_in[5]);
  or (_06161_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_06162_, _06161_, _06159_);
  and (_06164_, _06162_, _05881_);
  or (_06165_, _06164_, _06158_);
  or (_06166_, _06165_, _06154_);
  and (_06167_, _06166_, _05737_);
  or (_06169_, _06087_, p2_in[5]);
  or (_06172_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_06173_, _06172_, _06169_);
  and (_06174_, _06173_, _05881_);
  nor (_06175_, _06087_, p2_in[4]);
  and (_06177_, _06087_, _25300_);
  nor (_06179_, _06177_, _06175_);
  and (_06181_, _06179_, _05863_);
  or (_06182_, _06181_, _06174_);
  nor (_06183_, _06087_, p2_in[6]);
  not (_06185_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_06186_, _06087_, _06185_);
  nor (_06187_, _06186_, _06183_);
  and (_06188_, _06187_, _05868_);
  or (_06189_, _06087_, p2_in[7]);
  or (_06190_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_06191_, _06190_, _06189_);
  and (_06192_, _06191_, _05874_);
  or (_06193_, _06192_, _06188_);
  or (_06194_, _06193_, _06182_);
  and (_06195_, _06194_, _05896_);
  or (_06196_, _06195_, _06167_);
  and (_06197_, _06196_, _05876_);
  or (_06198_, _06197_, _06143_);
  and (_06199_, _06198_, _05953_);
  or (_06200_, _06087_, p0_in[1]);
  or (_06201_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_06202_, _06201_, _06200_);
  and (_06203_, _06202_, _05881_);
  nor (_06204_, _06087_, p0_in[0]);
  and (_06206_, _06087_, _25483_);
  nor (_06207_, _06206_, _06204_);
  and (_06208_, _06207_, _05863_);
  or (_06209_, _06208_, _06203_);
  or (_06210_, _06087_, p0_in[2]);
  or (_06211_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_06212_, _06211_, _06210_);
  and (_06213_, _06212_, _05868_);
  or (_06214_, _06087_, p0_in[3]);
  or (_06215_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_06216_, _06215_, _06214_);
  and (_06217_, _06216_, _05874_);
  or (_06218_, _06217_, _06213_);
  or (_06219_, _06218_, _06209_);
  and (_06220_, _06219_, _05896_);
  or (_06221_, _06087_, p1_in[2]);
  or (_06222_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_06223_, _06222_, _06221_);
  and (_06224_, _06223_, _05868_);
  or (_06225_, _06087_, p1_in[3]);
  or (_06226_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_06227_, _06226_, _06225_);
  and (_06228_, _06227_, _05874_);
  or (_06229_, _06228_, _06224_);
  or (_06230_, _06087_, p1_in[1]);
  or (_06231_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_06232_, _06231_, _06230_);
  and (_06234_, _06232_, _05881_);
  nor (_06235_, _06087_, p1_in[0]);
  and (_06236_, _06087_, _25400_);
  nor (_06237_, _06236_, _06235_);
  and (_06238_, _06237_, _05863_);
  or (_06239_, _06238_, _06234_);
  or (_06240_, _06239_, _06229_);
  and (_06241_, _06240_, _05737_);
  or (_06242_, _06241_, _06220_);
  and (_06243_, _06242_, _00168_);
  or (_06244_, _06087_, p1_in[5]);
  or (_06245_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_06246_, _06245_, _06244_);
  and (_06247_, _06246_, _05881_);
  nor (_06248_, _06087_, p1_in[4]);
  not (_06249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_06250_, _06087_, _06249_);
  nor (_06251_, _06250_, _06248_);
  and (_06252_, _06251_, _05863_);
  or (_06253_, _06252_, _06247_);
  nor (_06255_, _06087_, p1_in[6]);
  and (_06256_, _06087_, _25418_);
  nor (_06258_, _06256_, _06255_);
  and (_06259_, _06258_, _05868_);
  or (_06260_, _06087_, p1_in[7]);
  or (_06261_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_06262_, _06261_, _06260_);
  and (_06263_, _06262_, _05874_);
  or (_06265_, _06263_, _06259_);
  or (_06266_, _06265_, _06253_);
  and (_06268_, _06266_, _05737_);
  or (_06269_, _06087_, p0_in[5]);
  or (_06270_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_06272_, _06270_, _06269_);
  and (_06274_, _06272_, _05881_);
  nor (_06275_, _06087_, p0_in[4]);
  and (_06277_, _06087_, _25531_);
  nor (_06278_, _06277_, _06275_);
  and (_06279_, _06278_, _05863_);
  or (_06281_, _06279_, _06274_);
  nor (_06282_, _06087_, p0_in[6]);
  and (_06283_, _06087_, _25517_);
  nor (_06284_, _06283_, _06282_);
  and (_06285_, _06284_, _05868_);
  or (_06286_, _06087_, p0_in[7]);
  or (_06287_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_06288_, _06287_, _06286_);
  and (_06290_, _06288_, _05874_);
  or (_06291_, _06290_, _06285_);
  or (_06292_, _06291_, _06281_);
  and (_06294_, _06292_, _05896_);
  or (_06295_, _06294_, _06268_);
  and (_06296_, _06295_, _05876_);
  or (_06297_, _06296_, _06243_);
  and (_06298_, _06297_, _05963_);
  or (_06299_, _06298_, _06199_);
  or (_06300_, _06299_, _06067_);
  or (_06301_, _06300_, _05888_);
  and (_06302_, _06045_, _00260_);
  nor (_06303_, _06302_, _00184_);
  nand (_06304_, _05889_, _23594_);
  and (_06305_, _06304_, _06303_);
  and (_06306_, _06305_, _06301_);
  and (_06307_, _05868_, _23816_);
  or (_06308_, _06307_, _05876_);
  and (_06309_, _05863_, _24685_);
  and (_06310_, _05881_, _23892_);
  and (_06311_, _05874_, _23738_);
  or (_06312_, _06311_, _06310_);
  or (_06313_, _06312_, _06309_);
  or (_06314_, _06313_, _06308_);
  and (_06315_, _05868_, _24043_);
  or (_06316_, _06315_, _00168_);
  and (_06317_, _05863_, _23642_);
  and (_06318_, _05881_, _23939_);
  and (_06319_, _05874_, _26750_);
  or (_06320_, _06319_, _06318_);
  or (_06321_, _06320_, _06317_);
  or (_06322_, _06321_, _06316_);
  nand (_06323_, _06322_, _06314_);
  nor (_06324_, _06323_, _06303_);
  or (_06325_, _06324_, _06306_);
  and (_27305_, _06325_, _22762_);
  nor (_06327_, _26817_, _02444_);
  and (_06328_, _00168_, _00037_);
  and (_06329_, _06328_, _05863_);
  nor (_06330_, _02397_, _00014_);
  and (_06331_, _06330_, _06329_);
  and (_06333_, _06331_, _06327_);
  and (_06334_, _06333_, _00260_);
  not (_06335_, _24646_);
  and (_06336_, _05874_, _05876_);
  nor (_06337_, _06336_, _06335_);
  and (_06339_, _06337_, _00065_);
  nor (_06340_, _06339_, _06334_);
  and (_06341_, _06340_, _00178_);
  and (_06343_, _00259_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_06344_, _05963_, _05892_);
  and (_06345_, _06328_, _05874_);
  and (_06346_, _06345_, _06344_);
  and (_06347_, _06346_, _06343_);
  not (_06348_, _06347_);
  and (_06349_, _06333_, _00256_);
  and (_06350_, _06329_, _06001_);
  and (_06351_, _06350_, _06327_);
  and (_06352_, _06351_, _00278_);
  nor (_06353_, _06352_, _06349_);
  and (_06354_, _06353_, _06348_);
  nor (_06355_, _06354_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_06356_, _06355_);
  and (_06357_, _06356_, _06341_);
  and (_06358_, _06344_, _05868_);
  and (_06359_, _06358_, _06328_);
  and (_06361_, _06359_, _06343_);
  or (_06362_, _06361_, rst);
  nor (_27306_, _06362_, _06357_);
  and (_06363_, _05892_, _05735_);
  and (_06365_, _00168_, _05891_);
  and (_06366_, _06365_, _05863_);
  and (_06367_, _06366_, _06363_);
  nor (_06369_, _00168_, _00037_);
  and (_06371_, _06369_, _05863_);
  and (_06372_, _06371_, _06363_);
  or (_06373_, _06372_, _06367_);
  and (_06374_, _06365_, _05868_);
  and (_06375_, _06374_, _06363_);
  and (_06376_, _06369_, _05881_);
  and (_06377_, _06376_, _06363_);
  or (_06378_, _06377_, _06375_);
  nor (_06379_, _06378_, _06373_);
  and (_06380_, _06330_, _05900_);
  and (_06381_, _06380_, _06366_);
  and (_06382_, _06336_, _00037_);
  and (_06383_, _05937_, _05900_);
  and (_06384_, _06383_, _06382_);
  nor (_06385_, _06384_, _06381_);
  and (_06387_, _06366_, _06344_);
  and (_06388_, _06365_, _05874_);
  and (_06389_, _06388_, _06363_);
  nor (_06390_, _06389_, _06387_);
  and (_06392_, _06390_, _06385_);
  and (_06393_, _06392_, _06379_);
  and (_06394_, _06388_, _06344_);
  and (_06396_, _06365_, _05881_);
  and (_06397_, _06396_, _06344_);
  nor (_06399_, _06397_, _06394_);
  and (_06400_, _06376_, _06344_);
  and (_06402_, _06374_, _06344_);
  nor (_06404_, _06402_, _06400_);
  and (_06405_, _06404_, _06399_);
  and (_06406_, _06371_, _06344_);
  and (_06407_, _06382_, _06344_);
  nor (_06408_, _06407_, _06406_);
  and (_06409_, _05963_, _05736_);
  and (_06410_, _06409_, _06396_);
  and (_06411_, _06409_, _06366_);
  nor (_06412_, _06411_, _06410_);
  and (_06413_, _06412_, _06408_);
  and (_06414_, _06413_, _06405_);
  and (_06416_, _06414_, _06393_);
  or (_06417_, _06351_, _06333_);
  and (_06418_, _06329_, _05900_);
  or (_06419_, _06359_, _06346_);
  and (_06420_, _06344_, _05881_);
  and (_06421_, _06420_, _06328_);
  and (_06422_, _05937_, _06327_);
  and (_06423_, _06422_, _06329_);
  or (_06424_, _06423_, _06421_);
  or (_06425_, _06424_, _06419_);
  or (_06426_, _06425_, _06418_);
  nor (_06427_, _06426_, _06417_);
  and (_06428_, _06427_, _06416_);
  not (_06429_, _06428_);
  and (_06431_, _06429_, _06357_);
  not (_06432_, _06431_);
  and (_06433_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_06434_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_06435_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_06436_, _06435_, _06434_);
  and (_06437_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_06438_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_06439_, _06438_, _06437_);
  or (_06441_, _06439_, _06436_);
  and (_06442_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_06443_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_06444_, _06443_, _06442_);
  and (_06445_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_06447_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_06448_, _06447_, _06445_);
  or (_06449_, _06448_, _06444_);
  or (_06451_, _06449_, _06441_);
  and (_06452_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_06453_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_06454_, _06453_, _06452_);
  and (_06455_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_06456_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_06458_, _06456_, _06455_);
  or (_06459_, _06458_, _06454_);
  and (_06460_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_06462_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_06463_, _06462_, _06460_);
  and (_06464_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_06465_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_06466_, _06465_, _06464_);
  or (_06467_, _06466_, _06463_);
  or (_06469_, _06467_, _06459_);
  or (_06471_, _06469_, _06451_);
  and (_06472_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_06474_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_06475_, _06474_, _06472_);
  and (_06476_, _06421_, _26727_);
  and (_06477_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_06478_, _06477_, _06476_);
  or (_06479_, _06478_, _06475_);
  and (_06480_, _06418_, _05937_);
  and (_06481_, _06480_, _06157_);
  and (_06482_, _06331_, _05900_);
  and (_06483_, _06482_, _06191_);
  or (_06485_, _06483_, _06481_);
  and (_06486_, _06344_, _06329_);
  and (_06487_, _06486_, _06288_);
  and (_06488_, _06409_, _06329_);
  and (_06489_, _06488_, _06262_);
  or (_06490_, _06489_, _06487_);
  or (_06491_, _06490_, _06485_);
  or (_06493_, _06491_, _06479_);
  and (_06494_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_06495_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_06496_, _06495_, _06494_);
  or (_06497_, _06496_, _06493_);
  or (_06498_, _06497_, _06471_);
  and (_06499_, _06498_, _06357_);
  or (_06500_, _06499_, _06361_);
  or (_06501_, _06500_, _06433_);
  not (_06502_, _06361_);
  or (_06503_, _06502_, _00875_);
  and (_06504_, _06503_, _22762_);
  and (_27307_[7], _06504_, _06501_);
  and (_06505_, _23753_, _22946_);
  and (_06506_, _06505_, _23661_);
  and (_06507_, _06506_, _24010_);
  not (_06508_, _06507_);
  and (_06509_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and (_06510_, _06507_, _23898_);
  or (_25285_, _06510_, _06509_);
  and (_06511_, _02325_, _23656_);
  and (_06513_, _06511_, _24050_);
  not (_06514_, _06511_);
  and (_06515_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_25288_, _06515_, _06513_);
  and (_06517_, _02325_, _25078_);
  and (_06518_, _06517_, _23824_);
  not (_06520_, _06517_);
  and (_06522_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_27151_, _06522_, _06518_);
  and (_06524_, _02325_, _24282_);
  and (_06525_, _06524_, _23649_);
  not (_06527_, _06524_);
  and (_06529_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  or (_25295_, _06529_, _06525_);
  and (_06530_, _02325_, _23911_);
  and (_06531_, _06530_, _23898_);
  not (_06532_, _06530_);
  and (_06533_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  or (_25298_, _06533_, _06531_);
  and (_06534_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_06536_, _05705_, _23747_);
  or (_25344_, _06536_, _06534_);
  and (_06538_, _05429_, _23778_);
  and (_06539_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_25347_, _06539_, _06538_);
  and (_06540_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and (_06541_, _05705_, _23824_);
  or (_25351_, _06541_, _06540_);
  and (_06544_, _02325_, _24010_);
  and (_06545_, _06544_, _23946_);
  not (_06547_, _06544_);
  and (_06548_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_25357_, _06548_, _06545_);
  and (_06550_, _06544_, _23778_);
  and (_06551_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_25366_, _06551_, _06550_);
  and (_06552_, _02325_, _24085_);
  and (_06553_, _06552_, _23898_);
  not (_06554_, _06552_);
  and (_06555_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_27143_, _06555_, _06553_);
  and (_06557_, _05454_, _23778_);
  and (_06558_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_25392_, _06558_, _06557_);
  and (_06559_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_06561_, _05705_, _23707_);
  or (_25413_, _06561_, _06559_);
  and (_06563_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_06564_, _05705_, _24050_);
  or (_25424_, _06564_, _06563_);
  and (_06566_, _24581_, _26650_);
  or (_06567_, _02261_, _23950_);
  or (_06568_, _06567_, _06566_);
  nor (_06569_, _06568_, _24595_);
  nand (_06570_, _06569_, _24543_);
  or (_06572_, _05087_, _05090_);
  or (_06573_, _06572_, _26662_);
  or (_06574_, _06573_, _06570_);
  or (_06575_, _26654_, _26644_);
  or (_06576_, _06575_, _04952_);
  or (_06577_, _03276_, _26651_);
  and (_06578_, _26645_, _24448_);
  or (_06579_, _06578_, _04959_);
  or (_06580_, _06579_, _06577_);
  or (_06581_, _06580_, _06576_);
  or (_06582_, _06581_, _06574_);
  or (_06583_, _06582_, _04989_);
  or (_06584_, _24559_, _26572_);
  or (_06586_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _22766_);
  and (_06587_, _06586_, _22762_);
  and (_06588_, _06587_, _06584_);
  and (_26871_[0], _06588_, _06583_);
  and (_06589_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_06590_, _05705_, _23946_);
  or (_25428_, _06590_, _06589_);
  and (_06592_, _05454_, _23824_);
  and (_06593_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_25436_, _06593_, _06592_);
  and (_06594_, _05042_, _23747_);
  and (_06596_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_25440_, _06596_, _06594_);
  nor (_26897_[3], _00566_, rst);
  and (_06597_, _05454_, _23898_);
  and (_06598_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_25452_, _06598_, _06597_);
  and (_06599_, _23778_, _23665_);
  and (_06600_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or (_25454_, _06600_, _06599_);
  and (_06602_, _02325_, _23069_);
  and (_06603_, _06602_, _23649_);
  not (_06604_, _06602_);
  and (_06605_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  or (_25457_, _06605_, _06603_);
  and (_06606_, _06602_, _23898_);
  and (_06607_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  or (_25458_, _06607_, _06606_);
  and (_06608_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  and (_06609_, _05354_, _23747_);
  or (_25463_, _06609_, _06608_);
  and (_06610_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  and (_06612_, _05354_, _23946_);
  or (_25465_, _06612_, _06610_);
  and (_06613_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  and (_06614_, _05354_, _23649_);
  or (_25471_, _06614_, _06613_);
  and (_06615_, _01758_, _24085_);
  and (_06616_, _06615_, _23649_);
  not (_06618_, _06615_);
  and (_06619_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_25478_, _06619_, _06616_);
  and (_06620_, _06615_, _23747_);
  and (_06621_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_25487_, _06621_, _06620_);
  and (_06622_, _02326_, _24050_);
  and (_06623_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_25492_, _06623_, _06622_);
  and (_06624_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  and (_06625_, _05354_, _23707_);
  or (_25513_, _06625_, _06624_);
  nor (_26887_[6], _26811_, rst);
  and (_06626_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_06627_, _05705_, _23778_);
  or (_25522_, _06627_, _06626_);
  and (_06628_, _06615_, _24050_);
  and (_06629_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_27082_, _06629_, _06628_);
  and (_06630_, _06615_, _23946_);
  and (_06632_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_25535_, _06632_, _06630_);
  or (_06634_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_26915_, _06634_, _05209_);
  and (_06636_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  and (_06637_, _05354_, _23898_);
  or (_25567_, _06637_, _06636_);
  and (_06639_, _02325_, _24275_);
  and (_06641_, _06639_, _23747_);
  not (_06643_, _06639_);
  and (_06644_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_25569_, _06644_, _06641_);
  and (_06646_, _02325_, _24005_);
  and (_06647_, _06646_, _23747_);
  not (_06649_, _06646_);
  and (_06650_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_25575_, _06650_, _06647_);
  nor (_26897_[6], _00814_, rst);
  and (_06651_, _02325_, _23752_);
  and (_06652_, _06651_, _23946_);
  not (_06653_, _06651_);
  and (_06654_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  or (_25578_, _06654_, _06652_);
  and (_06655_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  and (_06656_, _04748_, _23824_);
  or (_25580_, _06656_, _06655_);
  and (_06657_, _24852_, _23747_);
  and (_06658_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or (_27205_, _06658_, _06657_);
  and (_06659_, _06615_, _23778_);
  and (_06661_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_25585_, _06661_, _06659_);
  and (_06662_, _06511_, _23778_);
  and (_06663_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_25589_, _06663_, _06662_);
  and (_06665_, _24275_, _23664_);
  and (_06666_, _06665_, _23824_);
  not (_06667_, _06665_);
  and (_06668_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  or (_27088_, _06668_, _06666_);
  and (_06669_, _06665_, _23898_);
  and (_06670_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  or (_25600_, _06670_, _06669_);
  and (_06671_, _06665_, _23778_);
  and (_06672_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or (_25606_, _06672_, _06671_);
  or (_06673_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_25614_, _06673_, _05467_);
  or (_06674_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_25617_, _06674_, _05463_);
  and (_06675_, _24593_, _24448_);
  or (_06676_, _04978_, _24591_);
  or (_06677_, _06676_, _05067_);
  or (_06678_, _06677_, _06675_);
  or (_06680_, _26652_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_06681_, _06680_, _24587_);
  or (_06682_, _26665_, _24559_);
  or (_06683_, _06682_, _06681_);
  or (_06685_, _06683_, _06678_);
  and (_06686_, _04973_, _24445_);
  and (_06687_, _24606_, _24447_);
  or (_06688_, _06687_, _04970_);
  or (_06690_, _06688_, _06686_);
  or (_06691_, _06690_, _06068_);
  or (_06692_, _06691_, _06685_);
  and (_06693_, _26614_, _24556_);
  or (_06694_, _06693_, _03316_);
  or (_06696_, _06694_, _05088_);
  or (_06697_, _26599_, _24617_);
  or (_06698_, _04969_, _04947_);
  or (_06699_, _06698_, _06697_);
  or (_06700_, _06699_, _06696_);
  or (_06701_, _06700_, _06692_);
  or (_06703_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _22766_);
  and (_06704_, _06703_, _22762_);
  and (_06706_, _06704_, _06584_);
  and (_26871_[1], _06706_, _06701_);
  and (_06708_, _25733_, _23898_);
  and (_06710_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_25628_, _06710_, _06708_);
  and (_06712_, _05042_, _23707_);
  and (_06713_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_25632_, _06713_, _06712_);
  and (_06715_, _06665_, _23946_);
  and (_06716_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or (_25637_, _06716_, _06715_);
  and (_06717_, _06665_, _23649_);
  and (_06718_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  or (_25643_, _06718_, _06717_);
  or (_06719_, _03274_, _26665_);
  or (_06720_, _05089_, _02381_);
  or (_06722_, _06720_, _06719_);
  or (_06723_, _04982_, _24617_);
  or (_06724_, _06723_, _06676_);
  and (_06725_, _24616_, _24448_);
  or (_06726_, _26661_, _24585_);
  or (_06727_, _06726_, _06725_);
  or (_06728_, _06727_, _06724_);
  or (_06729_, _06728_, _06690_);
  or (_06730_, _06729_, _06694_);
  or (_06731_, _06730_, _06722_);
  and (_06732_, _06731_, _22768_);
  and (_06733_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06734_, _24558_, _22766_);
  or (_06735_, _06734_, _06733_);
  or (_06736_, _06735_, _06732_);
  and (_26871_[2], _06736_, _22762_);
  or (_06737_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_25648_, _06737_, _05478_);
  and (_06738_, _02326_, _23946_);
  and (_06739_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_27153_, _06739_, _06738_);
  and (_06740_, _06665_, _23747_);
  and (_06741_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  or (_25655_, _06741_, _06740_);
  or (_06743_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_25658_, _06743_, _05474_);
  and (_06746_, _05701_, _23649_);
  and (_06747_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_25670_, _06747_, _06746_);
  and (_06749_, _05714_, _24050_);
  and (_06750_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  or (_25673_, _06750_, _06749_);
  and (_06751_, _23898_, _23665_);
  and (_06753_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  or (_25732_, _06753_, _06751_);
  and (_06755_, _02325_, _23986_);
  and (_06756_, _06755_, _23778_);
  not (_06757_, _06755_);
  and (_06759_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_25747_, _06759_, _06756_);
  and (_06761_, _02359_, _23824_);
  and (_06763_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  or (_25758_, _06763_, _06761_);
  and (_06764_, _05701_, _23707_);
  and (_06766_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_25767_, _06766_, _06764_);
  and (_06768_, _05701_, _24050_);
  and (_06769_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_25768_, _06769_, _06768_);
  and (_06771_, _06651_, _24050_);
  and (_06772_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  or (_25771_, _06772_, _06771_);
  not (_06773_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_06774_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not (_06775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor (_06776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_06778_, _06776_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_06779_, _06778_, _06775_);
  and (_06780_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _04488_);
  or (_06781_, _06780_, _06779_);
  nor (_06783_, _06781_, _06774_);
  nand (_06785_, _06783_, _06773_);
  nor (_06786_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor (_06788_, _06786_, _06783_);
  nand (_06789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_06791_, _06789_, _06788_);
  and (_06792_, _06791_, _22762_);
  and (_25778_, _06792_, _06785_);
  not (_06795_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and (_06796_, _04449_, _06795_);
  and (_06797_, _04567_, _04454_);
  and (_06798_, _06797_, _06796_);
  and (_06799_, _06798_, _04563_);
  not (_06800_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or (_06801_, _04569_, _06800_);
  nor (_06803_, _06801_, _06799_);
  or (_06804_, _06803_, _04462_);
  and (_25781_, _06804_, _22762_);
  nand (_06805_, _24504_, _24399_);
  nor (_06806_, _06805_, _24461_);
  and (_06807_, _22765_, _23839_);
  nand (_06808_, _06807_, _25644_);
  nor (_06809_, _06808_, _23863_);
  and (_06810_, _24526_, _24482_);
  and (_06811_, _06810_, _06809_);
  and (_06813_, _24431_, _24349_);
  and (_06814_, _06813_, _06811_);
  and (_26898_, _06814_, _06806_);
  and (_25786_, _06788_, _22762_);
  and (_06815_, _05410_, _24050_);
  and (_06816_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  or (_25792_, _06816_, _06815_);
  and (_06817_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  or (_06818_, _06817_, _04462_);
  nor (_06819_, _04490_, rst);
  and (_25796_, _06819_, _06818_);
  or (_06820_, _04780_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_06821_, _04780_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_06822_, _06821_, _06820_);
  nand (_06823_, _06822_, _22762_);
  nor (_25800_, _06823_, _04462_);
  not (_06825_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_06826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_06827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_06828_, _06778_, _06827_);
  or (_06829_, _06828_, _06780_);
  nor (_06830_, _06829_, _06826_);
  nand (_06832_, _06830_, _06825_);
  nor (_06834_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor (_06835_, _06834_, _06830_);
  nand (_06836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_06838_, _06836_, _06835_);
  and (_06839_, _06838_, _22762_);
  and (_25814_, _06839_, _06832_);
  and (_25815_, _06835_, _22762_);
  and (_06840_, _06665_, _23707_);
  and (_06841_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or (_25819_, _06841_, _06840_);
  and (_06842_, _04917_, _23898_);
  and (_06843_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_27108_, _06843_, _06842_);
  not (_06845_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_06846_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_06847_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _06846_);
  not (_06848_, _06847_);
  nor (_06849_, _04376_, _04609_);
  and (_06850_, _06849_, _06848_);
  and (_06851_, _06850_, _04628_);
  nor (_06852_, _06851_, _06845_);
  and (_06853_, _06851_, rxd_i);
  or (_06854_, _06853_, rst);
  or (_25872_, _06854_, _06852_);
  or (_06855_, _04605_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_06856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_06857_, _06856_, _04376_);
  or (_06858_, _06857_, _04579_);
  nand (_06860_, _06858_, _06855_);
  nand (_25874_, _06860_, _02066_);
  and (_06861_, _25618_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_06862_, _26599_, _26583_);
  or (_06863_, _06862_, _02380_);
  or (_06865_, _06863_, _06572_);
  or (_06867_, _04958_, _05080_);
  or (_06868_, _04979_, _04943_);
  or (_06870_, _06868_, _06867_);
  or (_06871_, _05070_, _26635_);
  or (_06872_, _06871_, _25622_);
  or (_06873_, _06872_, _05060_);
  or (_06874_, _06873_, _06870_);
  or (_06875_, _06874_, _06865_);
  and (_06876_, _06875_, _25644_);
  or (_26872_[0], _06876_, _06861_);
  and (_06877_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_06878_, _05398_, _23824_);
  or (_25944_, _06878_, _06877_);
  and (_06879_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_06880_, _05398_, _23898_);
  or (_25951_, _06880_, _06879_);
  and (_06881_, _05410_, _23707_);
  and (_06882_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  or (_25972_, _06882_, _06881_);
  and (_06883_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_06884_, _05398_, _23747_);
  or (_25999_, _06884_, _06883_);
  nor (_26897_[4], _00640_, rst);
  and (_06886_, _23785_, _23753_);
  and (_06888_, _06886_, _24005_);
  not (_06889_, _06888_);
  and (_06890_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  and (_06892_, _06888_, _23946_);
  or (_27014_, _06892_, _06890_);
  and (_06894_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  and (_06895_, _06888_, _23649_);
  or (_26025_, _06895_, _06894_);
  and (_06896_, _24766_, _24010_);
  not (_06897_, _06896_);
  and (_06898_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_06899_, _06896_, _23778_);
  or (_26050_, _06899_, _06898_);
  and (_06900_, _24766_, _24085_);
  not (_06902_, _06900_);
  and (_06903_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_06904_, _06900_, _23824_);
  or (_26054_, _06904_, _06903_);
  and (_06905_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_06906_, _06900_, _23747_);
  or (_26057_, _06906_, _06905_);
  and (_06907_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_06908_, _06900_, _23946_);
  or (_26059_, _06908_, _06907_);
  and (_06910_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_06912_, _06900_, _24050_);
  or (_26066_, _06912_, _06910_);
  and (_06914_, _04811_, _23824_);
  and (_06916_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or (_26068_, _06916_, _06914_);
  and (_06918_, _06886_, _23903_);
  not (_06919_, _06918_);
  and (_06920_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_06921_, _06918_, _24050_);
  or (_26071_, _06921_, _06920_);
  and (_06922_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_06924_, _06918_, _23707_);
  or (_27017_, _06924_, _06922_);
  and (_06927_, _06886_, _23991_);
  not (_06928_, _06927_);
  and (_06930_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and (_06931_, _06927_, _23898_);
  or (_26081_, _06931_, _06930_);
  and (_06933_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_06935_, _06927_, _23824_);
  or (_26087_, _06935_, _06933_);
  and (_06936_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_06937_, _06927_, _23946_);
  or (_26093_, _06937_, _06936_);
  nor (_27304_[0], \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_06940_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor (_06941_, _05727_, rst);
  and (_27304_[1], _06941_, _06940_);
  nor (_06942_, _05727_, _05726_);
  or (_06943_, _06942_, _05728_);
  and (_06944_, _05731_, _22762_);
  and (_27304_[2], _06944_, _06943_);
  nand (_06945_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_06946_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_06947_, _06946_, _06945_);
  nand (_06948_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_06949_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_06950_, _06949_, _06948_);
  and (_06951_, _06950_, _06947_);
  nand (_06952_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_06953_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_06954_, _06953_, _06952_);
  nand (_06955_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_06956_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_06957_, _06956_, _06955_);
  and (_06958_, _06957_, _06954_);
  and (_06959_, _06958_, _06951_);
  nand (_06961_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_06962_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_06963_, _06962_, _06961_);
  nand (_06964_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_06966_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_06967_, _06966_, _06964_);
  and (_06968_, _06967_, _06963_);
  nand (_06970_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand (_06971_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_06973_, _06971_, _06970_);
  nand (_06975_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand (_06976_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_06978_, _06976_, _06975_);
  and (_06979_, _06978_, _06973_);
  and (_06980_, _06979_, _06968_);
  and (_06981_, _06980_, _06959_);
  nand (_06982_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand (_06983_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_06984_, _06983_, _06982_);
  nand (_06985_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_06987_, _06421_, _00113_);
  and (_06988_, _06987_, _06985_);
  and (_06989_, _06988_, _06984_);
  nand (_06990_, _06480_, _06136_);
  nand (_06991_, _06482_, _06097_);
  and (_06992_, _06991_, _06990_);
  nand (_06993_, _06486_, _06207_);
  nand (_06995_, _06488_, _06237_);
  and (_06996_, _06995_, _06993_);
  and (_06997_, _06996_, _06992_);
  and (_06998_, _06997_, _06989_);
  not (_07000_, _06351_);
  or (_07001_, _07000_, _05860_);
  nand (_07002_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_07003_, _07002_, _07001_);
  and (_07004_, _07003_, _06998_);
  nand (_07005_, _07004_, _06981_);
  and (_07006_, _07005_, _06357_);
  nand (_07007_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_07008_, _07007_, _06502_);
  or (_07009_, _07008_, _07006_);
  or (_07010_, _06502_, _26565_);
  and (_07012_, _07010_, _22762_);
  and (_27307_[0], _07012_, _07009_);
  and (_07014_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_07015_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_07016_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_07017_, _07016_, _07015_);
  and (_07019_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_07020_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_07021_, _07020_, _07019_);
  or (_07023_, _07021_, _07017_);
  and (_07024_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_07025_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_07026_, _07025_, _07024_);
  and (_07027_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_07028_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_07029_, _07028_, _07027_);
  or (_07030_, _07029_, _07026_);
  or (_07031_, _07030_, _07023_);
  and (_07032_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_07033_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_07035_, _07033_, _07032_);
  and (_07036_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_07037_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_07038_, _07037_, _07036_);
  or (_07039_, _07038_, _07035_);
  and (_07040_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_07041_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_07042_, _07041_, _07040_);
  and (_07043_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_07044_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_07045_, _07044_, _07043_);
  or (_07046_, _07045_, _07042_);
  or (_07047_, _07046_, _07039_);
  or (_07048_, _07047_, _07031_);
  and (_07049_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_07050_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_07051_, _07050_, _07049_);
  and (_07052_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_07054_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_07056_, _07054_, _07052_);
  and (_07057_, _06421_, _00078_);
  and (_07058_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_07059_, _07058_, _07057_);
  or (_07060_, _07059_, _07056_);
  and (_07062_, _06480_, _06125_);
  and (_07063_, _06482_, _06092_);
  or (_07064_, _07063_, _07062_);
  and (_07065_, _06486_, _06202_);
  and (_07066_, _06488_, _06232_);
  or (_07067_, _07066_, _07065_);
  or (_07068_, _07067_, _07064_);
  or (_07069_, _07068_, _07060_);
  or (_07070_, _07069_, _07051_);
  or (_07071_, _07070_, _07048_);
  and (_07072_, _07071_, _06357_);
  or (_07073_, _07072_, _06361_);
  or (_07074_, _07073_, _07014_);
  nand (_07075_, _06361_, _00372_);
  and (_07076_, _07075_, _22762_);
  and (_27307_[1], _07076_, _07074_);
  and (_07077_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_07078_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_07079_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_07080_, _07079_, _07078_);
  and (_07082_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_07083_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_07084_, _07083_, _07082_);
  or (_07085_, _07084_, _07080_);
  and (_07087_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_07088_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_07090_, _07088_, _07087_);
  and (_07091_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_07093_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_07094_, _07093_, _07091_);
  or (_07095_, _07094_, _07090_);
  or (_07096_, _07095_, _07085_);
  and (_07097_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_07099_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or (_07100_, _07099_, _07097_);
  and (_07101_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_07102_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_07103_, _07102_, _07101_);
  or (_07104_, _07103_, _07100_);
  and (_07105_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_07107_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_07108_, _07107_, _07105_);
  and (_07109_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_07111_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_07112_, _07111_, _07109_);
  or (_07113_, _07112_, _07108_);
  or (_07114_, _07113_, _07104_);
  or (_07115_, _07114_, _07096_);
  and (_07116_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_07117_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_07118_, _07117_, _07116_);
  and (_07119_, _06421_, _00148_);
  and (_07120_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_07121_, _07120_, _07119_);
  or (_07122_, _07121_, _07118_);
  and (_07123_, _06480_, _06130_);
  and (_07124_, _06482_, _06105_);
  or (_07125_, _07124_, _07123_);
  and (_07126_, _06486_, _06212_);
  and (_07127_, _06488_, _06223_);
  or (_07128_, _07127_, _07126_);
  or (_07129_, _07128_, _07125_);
  or (_07130_, _07129_, _07122_);
  and (_07131_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_07132_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_07133_, _07132_, _07131_);
  or (_07134_, _07133_, _07130_);
  or (_07135_, _07134_, _07115_);
  and (_07136_, _07135_, _06357_);
  or (_07137_, _07136_, _06361_);
  or (_07138_, _07137_, _07077_);
  or (_07139_, _06502_, _00451_);
  and (_07140_, _07139_, _22762_);
  and (_27307_[2], _07140_, _07138_);
  and (_07141_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_07142_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_07143_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_07144_, _07143_, _07142_);
  and (_07145_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_07146_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_07147_, _07146_, _07145_);
  or (_07148_, _07147_, _07144_);
  and (_07149_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_07151_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_07152_, _07151_, _07149_);
  and (_07153_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_07154_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_07155_, _07154_, _07153_);
  or (_07156_, _07155_, _07152_);
  or (_07157_, _07156_, _07148_);
  and (_07158_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_07159_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or (_07160_, _07159_, _07158_);
  and (_07161_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_07162_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_07163_, _07162_, _07161_);
  or (_07164_, _07163_, _07160_);
  and (_07165_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_07166_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_07167_, _07166_, _07165_);
  and (_07168_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_07169_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_07170_, _07169_, _07168_);
  or (_07171_, _07170_, _07167_);
  or (_07172_, _07171_, _07164_);
  or (_07174_, _07172_, _07157_);
  and (_07175_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_07176_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_07177_, _07176_, _07175_);
  and (_07178_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_07179_, _06421_, _00030_);
  or (_07180_, _07179_, _07178_);
  or (_07181_, _07180_, _07177_);
  and (_07182_, _06480_, _06119_);
  and (_07183_, _06482_, _06110_);
  or (_07184_, _07183_, _07182_);
  and (_07186_, _06486_, _06216_);
  and (_07187_, _06488_, _06227_);
  or (_07188_, _07187_, _07186_);
  or (_07189_, _07188_, _07184_);
  or (_07190_, _07189_, _07181_);
  and (_07192_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_07193_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_07194_, _07193_, _07192_);
  or (_07196_, _07194_, _07190_);
  or (_07197_, _07196_, _07174_);
  and (_07198_, _07197_, _06357_);
  or (_07199_, _07198_, _06361_);
  or (_07200_, _07199_, _07141_);
  or (_07201_, _06502_, _00545_);
  and (_07202_, _07201_, _22762_);
  and (_27307_[3], _07202_, _07200_);
  and (_07204_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_07205_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand (_07206_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_07207_, _07206_, _07205_);
  nand (_07209_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand (_07210_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_07211_, _07210_, _07209_);
  and (_07212_, _07211_, _07207_);
  nand (_07213_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nand (_07214_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_07215_, _07214_, _07213_);
  nand (_07216_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand (_07217_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_07219_, _07217_, _07216_);
  and (_07220_, _07219_, _07215_);
  and (_07221_, _07220_, _07212_);
  nand (_07223_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand (_07224_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_07225_, _07224_, _07223_);
  nand (_07227_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_07229_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_07230_, _07229_, _07227_);
  and (_07232_, _07230_, _07225_);
  nand (_07233_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  nand (_07235_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_07236_, _07235_, _07233_);
  nand (_07238_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  nand (_07239_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_07240_, _07239_, _07238_);
  and (_07242_, _07240_, _07236_);
  and (_07243_, _07242_, _07232_);
  and (_07245_, _07243_, _07221_);
  nand (_07247_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_07248_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_07249_, _07248_, _07247_);
  nand (_07251_, _06421_, _00047_);
  nand (_07252_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_07254_, _07252_, _07251_);
  and (_07255_, _07254_, _07249_);
  nand (_07256_, _06480_, _06152_);
  nand (_07257_, _06482_, _06179_);
  and (_07258_, _07257_, _07256_);
  nand (_07259_, _06486_, _06278_);
  nand (_07260_, _06488_, _06251_);
  and (_07261_, _07260_, _07259_);
  and (_07262_, _07261_, _07258_);
  and (_07263_, _07262_, _07255_);
  nand (_07264_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nand (_07265_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_07266_, _07265_, _07264_);
  and (_07267_, _07266_, _07263_);
  and (_07268_, _07267_, _07245_);
  nor (_07269_, _06341_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_07270_, _07269_, _06355_);
  nor (_07271_, _07270_, _07268_);
  or (_07272_, _07271_, _06361_);
  or (_07273_, _07272_, _07204_);
  or (_07274_, _06502_, _00620_);
  and (_07275_, _07274_, _22762_);
  and (_27307_[4], _07275_, _07273_);
  and (_07276_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_07277_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_07279_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_07280_, _07279_, _07277_);
  and (_07283_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_07284_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_07285_, _07284_, _07283_);
  or (_07286_, _07285_, _07280_);
  and (_07288_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_07289_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_07291_, _07289_, _07288_);
  and (_07292_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_07293_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_07294_, _07293_, _07292_);
  or (_07295_, _07294_, _07291_);
  or (_07296_, _07295_, _07286_);
  and (_07297_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_07298_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_07299_, _07298_, _07297_);
  and (_07301_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_07302_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_07303_, _07302_, _07301_);
  or (_07304_, _07303_, _07299_);
  and (_07306_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_07307_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_07308_, _07307_, _07306_);
  and (_07309_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_07311_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_07312_, _07311_, _07309_);
  or (_07313_, _07312_, _07308_);
  or (_07314_, _07313_, _07304_);
  or (_07315_, _07314_, _07296_);
  and (_07316_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_07317_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_07318_, _07317_, _07316_);
  and (_07319_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_07320_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_07321_, _07320_, _07319_);
  not (_07322_, _26826_);
  and (_07323_, _06421_, _07322_);
  and (_07324_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_07325_, _07324_, _07323_);
  or (_07326_, _07325_, _07321_);
  and (_07327_, _06480_, _06162_);
  and (_07328_, _06482_, _06173_);
  or (_07329_, _07328_, _07327_);
  and (_07330_, _06486_, _06272_);
  and (_07331_, _06488_, _06246_);
  or (_07332_, _07331_, _07330_);
  or (_07333_, _07332_, _07329_);
  or (_07334_, _07333_, _07326_);
  or (_07335_, _07334_, _07318_);
  or (_07336_, _07335_, _07315_);
  and (_07337_, _07336_, _06357_);
  or (_07339_, _07337_, _06361_);
  or (_07340_, _07339_, _07276_);
  or (_07341_, _06502_, _00708_);
  and (_07343_, _07341_, _22762_);
  and (_27307_[5], _07343_, _07340_);
  and (_07344_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_07345_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand (_07346_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_07347_, _07346_, _07345_);
  nand (_07348_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nand (_07349_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_07350_, _07349_, _07348_);
  and (_07351_, _07350_, _07347_);
  nand (_07352_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nand (_07353_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_07354_, _07353_, _07352_);
  and (_07355_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_07356_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nor (_07357_, _07356_, _07355_);
  and (_07358_, _07357_, _07354_);
  and (_07360_, _07358_, _07351_);
  nand (_07361_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  nand (_07362_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_07364_, _07362_, _07361_);
  nand (_07365_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  nand (_07366_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_07367_, _07366_, _07365_);
  and (_07368_, _07367_, _07364_);
  nand (_07369_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_07370_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_07371_, _07370_, _07369_);
  nand (_07372_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_07373_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_07374_, _07373_, _07372_);
  and (_07375_, _07374_, _07371_);
  and (_07376_, _07375_, _07368_);
  and (_07377_, _07376_, _07360_);
  nand (_07378_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand (_07379_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_07380_, _07379_, _07378_);
  not (_07381_, _26788_);
  nand (_07382_, _06421_, _07381_);
  nand (_07383_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_07384_, _07383_, _07382_);
  and (_07385_, _07384_, _07380_);
  nand (_07386_, _06480_, _06146_);
  nand (_07387_, _06482_, _06187_);
  and (_07388_, _07387_, _07386_);
  nand (_07389_, _06486_, _06284_);
  nand (_07391_, _06488_, _06258_);
  and (_07392_, _07391_, _07389_);
  and (_07393_, _07392_, _07388_);
  and (_07394_, _07393_, _07385_);
  nand (_07395_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand (_07397_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_07398_, _07397_, _07395_);
  and (_07399_, _07398_, _07394_);
  and (_07400_, _07399_, _07377_);
  nor (_07401_, _06341_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or (_07403_, _07401_, _06355_);
  nor (_07404_, _07403_, _07400_);
  or (_07405_, _07404_, _06361_);
  or (_07406_, _07405_, _07344_);
  nand (_07407_, _06361_, _00793_);
  and (_07409_, _07407_, _22762_);
  and (_27307_[6], _07409_, _07406_);
  and (_07410_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_07411_, _06927_, _24050_);
  or (_26132_, _07411_, _07410_);
  or (_07412_, _04891_, _23642_);
  nand (_07413_, _04882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_07414_, _04882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_07415_, _07414_, _26097_);
  and (_07417_, _07415_, _07413_);
  and (_07418_, _04864_, _24309_);
  or (_07419_, _07418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_07420_, _05158_, _04864_);
  not (_07421_, _07420_);
  and (_07422_, _07421_, _04860_);
  and (_07423_, _07422_, _07419_);
  and (_07424_, _04876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_07426_, _07424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_07427_, _07424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_07429_, _07427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_07430_, _07429_, _07426_);
  or (_07431_, _07430_, _07423_);
  or (_07432_, _07431_, _07417_);
  or (_07433_, _07432_, _24299_);
  and (_07434_, _07433_, _24294_);
  and (_07436_, _07434_, _07412_);
  and (_07437_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_07438_, _07437_, _07436_);
  and (_26617_, _07438_, _22762_);
  and (_07439_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  and (_07440_, _02298_, _23747_);
  or (_26642_, _07440_, _07439_);
  and (_07442_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  and (_07443_, _02298_, _23649_);
  or (_26649_, _07443_, _07442_);
  and (_07444_, _04917_, _23778_);
  and (_07446_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_26664_, _07446_, _07444_);
  and (_07447_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  and (_07448_, _02298_, _23946_);
  or (_26667_, _07448_, _07447_);
  or (_07449_, _04891_, _23939_);
  not (_07450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_07451_, _07420_, _26099_);
  nor (_07452_, _07451_, _07450_);
  and (_07454_, _07451_, _07450_);
  or (_07455_, _07454_, _07452_);
  and (_07456_, _07455_, _04861_);
  and (_07457_, _05158_, _24300_);
  or (_07458_, _07457_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_07459_, _07458_, _24302_);
  nor (_07460_, _07459_, _05151_);
  or (_07461_, _05164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_07462_, _05165_, _26098_);
  and (_07463_, _07462_, _07461_);
  or (_07464_, _07463_, _07460_);
  or (_07465_, _07464_, _07456_);
  or (_07466_, _07465_, _24299_);
  and (_07467_, _07466_, _24294_);
  and (_07468_, _07467_, _07449_);
  and (_07469_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_07470_, _07469_, _07468_);
  and (_26690_, _07470_, _22762_);
  and (_07471_, _01809_, _24010_);
  and (_07472_, _07471_, _23946_);
  not (_07473_, _07471_);
  and (_07474_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  or (_27107_, _07474_, _07472_);
  and (_07475_, _04811_, _23707_);
  and (_07476_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or (_26706_, _07476_, _07475_);
  and (_07477_, _07471_, _23649_);
  and (_07478_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or (_26720_, _07478_, _07477_);
  and (_07479_, _07471_, _23824_);
  and (_07480_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or (_26726_, _07480_, _07479_);
  and (_07482_, _07471_, _23778_);
  and (_07483_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or (_26731_, _07483_, _07482_);
  and (_07484_, _05445_, _24050_);
  and (_07486_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  or (_26748_, _07486_, _07484_);
  and (_07488_, _05445_, _23946_);
  and (_07489_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or (_26764_, _07489_, _07488_);
  and (_07492_, _24329_, _24201_);
  not (_07493_, _07492_);
  and (_07494_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and (_07496_, _07492_, _24050_);
  or (_26769_, _07496_, _07494_);
  and (_07497_, _25142_, _23649_);
  and (_07499_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  or (_26771_, _07499_, _07497_);
  and (_07500_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_07501_, _24128_, _24043_);
  not (_07502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_07503_, _25684_, _07502_);
  and (_07504_, _25684_, _07502_);
  or (_07505_, _07504_, _07503_);
  or (_07506_, _07505_, _24127_);
  and (_07508_, _07506_, _24166_);
  and (_07509_, _07508_, _07501_);
  or (_26774_, _07509_, _07500_);
  and (_07510_, _25733_, _23824_);
  and (_07511_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_26780_, _07511_, _07510_);
  and (_26860_[1], _23866_, _22762_);
  and (_07513_, _04760_, _23069_);
  not (_07514_, _07513_);
  and (_07515_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and (_07516_, _07513_, _23898_);
  or (_26963_, _07516_, _07515_);
  and (_26860_[2], _24436_, _22762_);
  and (_07517_, _05445_, _23747_);
  and (_07518_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or (_26805_, _07518_, _07517_);
  and (_07519_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and (_07521_, _07492_, _23946_);
  or (_26828_, _07521_, _07519_);
  and (_07522_, _05445_, _23898_);
  and (_07524_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  or (_26834_, _07524_, _07522_);
  and (_07525_, _06886_, _24275_);
  not (_07526_, _07525_);
  and (_07527_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  and (_07530_, _07525_, _23778_);
  or (_00090_, _07530_, _07527_);
  and (_26910_, _02443_, _22762_);
  and (_26911_[7], _23706_, _22762_);
  nor (_26913_[2], _00168_, rst);
  and (_07533_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  and (_07534_, _07525_, _23898_);
  or (_00200_, _07534_, _07533_);
  and (_07536_, _01809_, _25078_);
  and (_07537_, _07536_, _23778_);
  not (_07539_, _07536_);
  and (_07541_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or (_00203_, _07541_, _07537_);
  and (_07542_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  and (_07543_, _07525_, _23649_);
  or (_00206_, _07543_, _07542_);
  and (_07544_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  and (_07545_, _07525_, _23946_);
  or (_00269_, _07545_, _07544_);
  and (_07547_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  and (_07550_, _07525_, _23707_);
  or (_00275_, _07550_, _07547_);
  and (_07551_, _24766_, _23784_);
  not (_07552_, _07551_);
  and (_07553_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  and (_07554_, _07551_, _23778_);
  or (_00279_, _07554_, _07553_);
  nor (_26887_[2], _00163_, rst);
  and (_07555_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  and (_07556_, _07551_, _23824_);
  or (_00296_, _07556_, _07555_);
  and (_07557_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and (_07558_, _07551_, _23649_);
  or (_00299_, _07558_, _07557_);
  and (_07559_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  and (_07560_, _07551_, _24050_);
  or (_00309_, _07560_, _07559_);
  and (_26911_[0], _23777_, _22762_);
  and (_26911_[1], _23897_, _22762_);
  and (_26911_[2], _23823_, _22762_);
  and (_26911_[3], _23746_, _22762_);
  and (_26911_[4], _23648_, _22762_);
  and (_26911_[5], _23945_, _22762_);
  and (_26911_[6], _24049_, _22762_);
  and (_07562_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  and (_07563_, _07551_, _23707_);
  or (_00385_, _07563_, _07562_);
  nor (_26913_[0], _00134_, rst);
  nor (_26913_[1], _00099_, rst);
  nor (_07566_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_07568_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _23978_);
  nor (_07570_, _07568_, _07566_);
  not (_07572_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_07574_, _00587_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_07576_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _23978_);
  nor (_07577_, _07576_, _07574_);
  and (_07578_, _07577_, _07572_);
  nor (_07580_, _07577_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_07581_, _07580_, _07578_);
  not (_07582_, _07581_);
  nor (_07583_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_07584_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _23978_);
  nor (_07585_, _07584_, _07583_);
  not (_07586_, _07585_);
  nor (_07588_, _00495_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_07589_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _23978_);
  nor (_07590_, _07589_, _07588_);
  and (_07591_, _07590_, _07586_);
  nand (_07592_, _07591_, _07582_);
  and (_07594_, _07592_, _07570_);
  nor (_07597_, _07590_, _07586_);
  not (_07599_, _07597_);
  not (_07600_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_07601_, _07577_, _07600_);
  and (_07603_, _07577_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_07605_, _07603_, _07601_);
  nor (_07606_, _07605_, _07599_);
  and (_07608_, _07590_, _07585_);
  not (_07610_, _07608_);
  not (_07612_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_07613_, _07577_, _07612_);
  nor (_07615_, _07577_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_07616_, _07615_, _07613_);
  nor (_07618_, _07616_, _07610_);
  nor (_07619_, _07618_, _07606_);
  not (_07621_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_07623_, _07577_, _07621_);
  nor (_07624_, _07590_, _07585_);
  not (_07626_, _07624_);
  nor (_07628_, _07577_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_07631_, _07628_, _07626_);
  or (_07632_, _07631_, _07623_);
  and (_07634_, _07632_, _07619_);
  and (_07636_, _07634_, _07594_);
  not (_07637_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_07639_, _07577_, _07637_);
  nor (_07641_, _07577_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_07642_, _07641_, _07639_);
  nor (_07643_, _07642_, _07610_);
  nor (_07645_, _07643_, _07570_);
  and (_07647_, _07577_, \oc8051_symbolic_cxrom1.regvalid [12]);
  not (_07648_, _07577_);
  and (_07649_, _07648_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_07650_, _07649_, _07647_);
  not (_07652_, _07650_);
  nand (_07653_, _07652_, _07591_);
  and (_07655_, _07577_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_07657_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_07659_, _07577_, _07657_);
  nor (_07660_, _07659_, _07655_);
  nor (_07662_, _07660_, _07599_);
  nor (_07663_, _07577_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not (_07664_, _07663_);
  not (_07665_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_07666_, _07577_, _07665_);
  nor (_07667_, _07666_, _07626_);
  and (_07668_, _07667_, _07664_);
  nor (_07669_, _07668_, _07662_);
  and (_07670_, _07669_, _07653_);
  and (_07671_, _07670_, _07645_);
  nor (_07672_, _07671_, _07636_);
  not (_07673_, _07672_);
  and (_07674_, _07673_, word_in[7]);
  not (_07675_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_07676_, _07570_, _07675_);
  or (_07677_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_07678_, _07677_, _07676_);
  and (_07679_, _07678_, _07624_);
  or (_07681_, _07679_, _07577_);
  not (_07682_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_07684_, _07570_, _07682_);
  or (_07685_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_07686_, _07685_, _07684_);
  and (_07687_, _07686_, _07608_);
  not (_07689_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_07691_, _07570_, _07689_);
  or (_07692_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_07693_, _07692_, _07691_);
  and (_07695_, _07693_, _07591_);
  not (_07696_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_07698_, _07570_, _07696_);
  or (_07700_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_07701_, _07700_, _07698_);
  and (_07703_, _07701_, _07597_);
  or (_07704_, _07703_, _07695_);
  or (_07706_, _07704_, _07687_);
  or (_07707_, _07706_, _07681_);
  not (_07709_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_07710_, _07570_, _07709_);
  or (_07711_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_07713_, _07711_, _07710_);
  and (_07714_, _07713_, _07624_);
  or (_07715_, _07714_, _07648_);
  not (_07717_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_07718_, _07570_, _07717_);
  or (_07720_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_07721_, _07720_, _07718_);
  and (_07722_, _07721_, _07591_);
  not (_07723_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_07725_, _07570_, _07723_);
  or (_07726_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_07727_, _07726_, _07725_);
  and (_07728_, _07727_, _07608_);
  or (_07730_, _07728_, _07722_);
  not (_07731_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_07732_, _07570_, _07731_);
  or (_07733_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_07734_, _07733_, _07732_);
  and (_07735_, _07734_, _07597_);
  or (_07736_, _07735_, _07730_);
  or (_07738_, _07736_, _07715_);
  and (_07740_, _07738_, _07707_);
  and (_07742_, _07740_, _07672_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _07742_, _07674_);
  and (_07743_, _24085_, _23664_);
  and (_07745_, _07743_, _23898_);
  not (_07747_, _07743_);
  and (_07748_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  or (_27072_, _07748_, _07745_);
  not (_07749_, _07570_);
  and (_07751_, _07585_, _07749_);
  not (_07753_, _07751_);
  and (_07754_, _07585_, _07570_);
  and (_07755_, _07754_, _07590_);
  nor (_07756_, _07754_, _07590_);
  nor (_07757_, _07756_, _07755_);
  not (_07758_, _07757_);
  nor (_07759_, _07758_, _07616_);
  nor (_07760_, _07755_, _07648_);
  not (_07761_, _07590_);
  nor (_07762_, _07761_, _07577_);
  and (_07763_, _07754_, _07762_);
  nor (_07764_, _07763_, _07760_);
  and (_07766_, _07764_, _07758_);
  and (_07768_, _07766_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_07770_, _07764_, _07757_);
  and (_07772_, _07770_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_07774_, _07772_, _07768_);
  nor (_07776_, _07774_, _07759_);
  nor (_07778_, _07776_, _07753_);
  nor (_07780_, _07585_, _07570_);
  not (_07782_, _07780_);
  nor (_07783_, _07758_, _07581_);
  and (_07784_, _07766_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_07785_, _07770_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_07786_, _07785_, _07784_);
  nor (_07787_, _07786_, _07783_);
  nor (_07788_, _07787_, _07782_);
  nor (_07789_, _07788_, _07778_);
  and (_07790_, _07586_, _07570_);
  not (_07791_, _07790_);
  nor (_07792_, _07758_, _07642_);
  and (_07793_, _07766_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_07794_, _07770_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_07795_, _07794_, _07793_);
  nor (_07796_, _07795_, _07792_);
  nor (_07798_, _07796_, _07791_);
  not (_07799_, _07754_);
  nor (_07801_, _07758_, _07650_);
  and (_07803_, _07766_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_07804_, _07770_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_07806_, _07804_, _07803_);
  nor (_07807_, _07806_, _07801_);
  nor (_07808_, _07807_, _07799_);
  nor (_07809_, _07808_, _07798_);
  and (_07810_, _07809_, _07789_);
  or (_07811_, _07780_, _07754_);
  not (_07812_, _07811_);
  not (_07813_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_07814_, _07570_, _07813_);
  or (_07815_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_07816_, _07815_, _07814_);
  and (_07817_, _07816_, _07812_);
  not (_07819_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_07821_, _07570_, _07819_);
  or (_07822_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_07824_, _07822_, _07821_);
  and (_07825_, _07824_, _07811_);
  or (_07826_, _07825_, _07817_);
  and (_07827_, _07826_, _07770_);
  not (_07829_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_07831_, _07570_, _07829_);
  or (_07833_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_07835_, _07833_, _07831_);
  and (_07836_, _07835_, _07812_);
  not (_07837_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_07839_, _07570_, _07837_);
  or (_07840_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_07841_, _07840_, _07839_);
  and (_07842_, _07841_, _07811_);
  or (_07843_, _07842_, _07836_);
  and (_07844_, _07843_, _07766_);
  and (_07845_, _07757_, _07648_);
  not (_07846_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_07847_, _07570_, _07846_);
  or (_07848_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_07849_, _07848_, _07847_);
  and (_07850_, _07849_, _07812_);
  not (_07852_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_07853_, _07570_, _07852_);
  or (_07855_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_07856_, _07855_, _07853_);
  and (_07857_, _07856_, _07811_);
  or (_07858_, _07857_, _07850_);
  and (_07859_, _07858_, _07845_);
  and (_07860_, _07757_, _07577_);
  not (_07861_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_07862_, _07570_, _07861_);
  or (_07863_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_07864_, _07863_, _07862_);
  and (_07865_, _07864_, _07812_);
  not (_07866_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_07867_, _07570_, _07866_);
  or (_07868_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_07869_, _07868_, _07867_);
  and (_07870_, _07869_, _07811_);
  or (_07871_, _07870_, _07865_);
  and (_07872_, _07871_, _07860_);
  or (_07873_, _07872_, _07859_);
  or (_07874_, _07873_, _07844_);
  nor (_07875_, _07874_, _07827_);
  nor (_07876_, _07875_, _07810_);
  and (_07877_, _07810_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _07877_, _07876_);
  nor (_07878_, _07608_, _07624_);
  and (_07879_, _07608_, _07577_);
  nor (_07880_, _07608_, _07577_);
  nor (_07881_, _07880_, _07879_);
  nor (_07882_, _07881_, _07878_);
  and (_07883_, _07882_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_07884_, _07883_);
  not (_07885_, _07878_);
  nor (_07886_, _07885_, _07581_);
  and (_07887_, _07881_, _07885_);
  and (_07888_, _07887_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_07889_, _07888_, _07886_);
  and (_07890_, _07889_, _07884_);
  nor (_07891_, _07890_, _07799_);
  nor (_07892_, _07885_, _07616_);
  and (_07893_, _07887_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_07895_, _07882_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_07896_, _07895_, _07893_);
  nor (_07897_, _07896_, _07892_);
  nor (_07898_, _07897_, _07791_);
  nor (_07899_, _07898_, _07891_);
  nor (_07900_, _07885_, _07642_);
  and (_07901_, _07882_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_07902_, _07887_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_07903_, _07902_, _07901_);
  nor (_07904_, _07903_, _07900_);
  nor (_07905_, _07904_, _07782_);
  and (_07906_, _07882_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not (_07907_, _07906_);
  nor (_07908_, _07885_, _07650_);
  and (_07909_, _07887_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_07910_, _07909_, _07908_);
  and (_07911_, _07910_, _07907_);
  nor (_07912_, _07911_, _07753_);
  nor (_07913_, _07912_, _07905_);
  and (_07914_, _07913_, _07899_);
  not (_07915_, _07881_);
  and (_07916_, _07686_, _07591_);
  and (_07917_, _07678_, _07577_);
  or (_07918_, _07917_, _07916_);
  and (_07919_, _07693_, _07597_);
  and (_07920_, _07701_, _07624_);
  or (_07921_, _07920_, _07919_);
  or (_07922_, _07921_, _07918_);
  and (_07923_, _07922_, _07915_);
  and (_07924_, _07721_, _07597_);
  and (_07926_, _07734_, _07624_);
  or (_07927_, _07926_, _07924_);
  and (_07928_, _07727_, _07591_);
  and (_07929_, _07713_, _07608_);
  or (_07930_, _07929_, _07928_);
  or (_07931_, _07930_, _07927_);
  and (_07932_, _07931_, _07881_);
  nor (_07933_, _07932_, _07923_);
  nor (_07934_, _07933_, _07914_);
  and (_07935_, _07914_, word_in[23]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _07935_, _07934_);
  and (_07936_, _05281_, _23824_);
  and (_07937_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_00562_, _07937_, _07936_);
  nor (_07938_, _07782_, _07590_);
  and (_07939_, _07938_, _07601_);
  not (_07940_, _07938_);
  nand (_07941_, _07782_, _07590_);
  and (_07942_, _07941_, _07940_);
  not (_07943_, _07942_);
  nor (_07945_, _07943_, _07581_);
  nor (_07946_, _07941_, _07577_);
  and (_07947_, _07941_, _07577_);
  nor (_07948_, _07947_, _07946_);
  and (_07949_, _07948_, _07943_);
  and (_07950_, _07949_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_07951_, _07948_, _07942_);
  and (_07952_, _07951_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_07953_, _07952_, _07950_);
  nor (_07954_, _07953_, _07945_);
  nor (_07955_, _07954_, _07753_);
  nor (_07956_, _07955_, _07939_);
  nor (_07957_, _07943_, _07616_);
  and (_07958_, _07951_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_07959_, _07958_, _07957_);
  nor (_07960_, _07959_, _07782_);
  nor (_07961_, _07943_, _07642_);
  and (_07962_, _07949_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_07963_, _07951_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_07964_, _07963_, _07962_);
  nor (_07965_, _07964_, _07961_);
  nor (_07966_, _07965_, _07799_);
  nor (_07967_, _07943_, _07650_);
  and (_07968_, _07949_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_07969_, _07951_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_07970_, _07969_, _07968_);
  nor (_07971_, _07970_, _07967_);
  nor (_07972_, _07971_, _07791_);
  or (_07973_, _07972_, _07966_);
  nor (_07974_, _07973_, _07960_);
  and (_07975_, _07974_, _07956_);
  and (_07976_, _07824_, _07812_);
  and (_07977_, _07816_, _07811_);
  or (_07978_, _07977_, _07976_);
  and (_07979_, _07978_, _07951_);
  and (_07980_, _07841_, _07812_);
  and (_07981_, _07835_, _07811_);
  or (_07982_, _07981_, _07980_);
  and (_07983_, _07982_, _07949_);
  and (_07984_, _07942_, _07648_);
  and (_07985_, _07856_, _07812_);
  and (_07986_, _07849_, _07811_);
  or (_07987_, _07986_, _07985_);
  and (_07988_, _07987_, _07984_);
  and (_07989_, _07869_, _07812_);
  and (_07990_, _07864_, _07811_);
  or (_07991_, _07990_, _07989_);
  and (_07992_, _07947_, _07940_);
  and (_07993_, _07992_, _07991_);
  or (_07994_, _07993_, _07988_);
  or (_07996_, _07994_, _07983_);
  nor (_07997_, _07996_, _07979_);
  nor (_07998_, _07997_, _07975_);
  and (_07999_, _07975_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _07999_, _07998_);
  and (_08000_, _07590_, _07577_);
  or (_08001_, _08000_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_26842_[15], _08001_, _22762_);
  and (_08002_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_08003_, _06896_, _23824_);
  or (_00617_, _08003_, _08002_);
  and (_08004_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_08005_, _06896_, _23649_);
  or (_00626_, _08005_, _08004_);
  and (_08006_, _07914_, _22762_);
  and (_08007_, _08006_, _07878_);
  and (_08008_, _08007_, _07881_);
  and (_08009_, _08008_, _07790_);
  and (_08010_, _07810_, _22762_);
  and (_08011_, _08010_, _07751_);
  and (_08012_, _08011_, _07860_);
  and (_08013_, _07636_, _22762_);
  and (_08014_, _08013_, _07585_);
  nor (_08015_, _07672_, rst);
  and (_08016_, _08015_, _08000_);
  and (_08017_, _08016_, _08014_);
  nor (_08018_, _08017_, _07723_);
  and (_08019_, _08015_, word_in[7]);
  and (_08020_, _08019_, _08017_);
  or (_08021_, _08020_, _08018_);
  or (_08022_, _08021_, _08012_);
  not (_08023_, _08012_);
  or (_08024_, _08023_, word_in[15]);
  and (_08025_, _08024_, _08022_);
  or (_08026_, _08025_, _08009_);
  and (_08027_, _08000_, _07780_);
  and (_08028_, _07975_, _22762_);
  and (_08029_, _08028_, _08027_);
  not (_08030_, _08029_);
  not (_08031_, _08009_);
  and (_08033_, _08006_, word_in[23]);
  or (_08034_, _08033_, _08031_);
  and (_08035_, _08034_, _08030_);
  and (_08036_, _08035_, _08026_);
  and (_08037_, _08029_, word_in[31]);
  or (_26849_[7], _08037_, _08036_);
  or (_08038_, _07949_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_26859_, _08038_, _22762_);
  not (_08039_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08040_, _07626_, _07577_);
  nand (_08041_, _08040_, _08039_);
  or (_08042_, _08041_, _07879_);
  and (_26842_[1], _08042_, _22762_);
  and (_08043_, _24329_, _23076_);
  and (_08044_, _08043_, _24050_);
  not (_08045_, _08043_);
  and (_08046_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_27212_, _08046_, _08044_);
  and (_08047_, _05410_, _23778_);
  and (_08048_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or (_27213_, _08048_, _08047_);
  and (_08050_, _07755_, _07577_);
  not (_08051_, _08040_);
  nor (_08052_, _08051_, _08050_);
  and (_08053_, _07984_, _07751_);
  nor (_08054_, _08053_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_08055_, _08054_, _08052_);
  and (_26842_[2], _08055_, _22762_);
  not (_08056_, _07766_);
  and (_08057_, _07984_, _07754_);
  or (_08058_, _07590_, _07577_);
  or (_08059_, _08058_, _07751_);
  and (_08060_, _08059_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_08061_, _08060_, _08057_);
  and (_08062_, _08061_, _08056_);
  and (_08063_, _07601_, _07624_);
  or (_08064_, _08063_, _08053_);
  or (_08065_, _08064_, _08062_);
  and (_08066_, _08065_, _08052_);
  or (_08067_, _08063_, _08061_);
  and (_08068_, _08067_, _08050_);
  or (_08069_, _08068_, _08051_);
  or (_08070_, _08069_, _08066_);
  and (_26842_[3], _08070_, _22762_);
  and (_08071_, _08043_, _23707_);
  and (_08072_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_00764_, _08072_, _08071_);
  and (_08073_, _07780_, _07762_);
  or (_08074_, _08073_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_08075_, _08074_, _08058_);
  or (_08076_, _08075_, _08057_);
  and (_08077_, _08076_, _08056_);
  and (_08078_, _08074_, _08050_);
  and (_08079_, _07790_, _07984_);
  and (_08080_, _07938_, _07648_);
  and (_08081_, _08080_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_08082_, _08081_, _08079_);
  or (_08083_, _08082_, _08078_);
  or (_08084_, _08083_, _08053_);
  or (_08085_, _08084_, _08077_);
  and (_26842_[4], _08085_, _22762_);
  and (_08087_, _02200_, _23824_);
  and (_08088_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_00828_, _08088_, _08087_);
  and (_08091_, _02321_, _23898_);
  and (_08093_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or (_27138_, _08093_, _08091_);
  or (_08095_, _07760_, _07946_);
  or (_08096_, _08095_, _08050_);
  not (_08097_, _07880_);
  or (_08098_, _08073_, _08057_);
  or (_08099_, _08098_, _08097_);
  and (_08101_, _08099_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08102_, _08053_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08104_, _07790_, _07762_);
  and (_08105_, _08051_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08106_, _08105_, _08104_);
  or (_08108_, _08106_, _08102_);
  or (_08109_, _08108_, _08101_);
  and (_08111_, _08109_, _08096_);
  or (_08112_, _08105_, _08053_);
  or (_08113_, _08112_, _08098_);
  or (_08114_, _08113_, _08111_);
  and (_26842_[5], _08114_, _22762_);
  and (_08116_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  and (_08117_, _05199_, _23824_);
  or (_00874_, _08117_, _08116_);
  and (_08119_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  and (_08120_, _05199_, _23649_);
  or (_00921_, _08120_, _08119_);
  nor (_08121_, _07880_, _08050_);
  and (_08122_, _07751_, _07762_);
  or (_08123_, _08122_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08124_, _08123_, _08121_);
  and (_08125_, _08098_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08126_, _08125_, _08104_);
  or (_08127_, _08126_, _08124_);
  and (_08128_, _08127_, _08095_);
  and (_08129_, _08123_, _08050_);
  and (_08130_, _08053_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08132_, _08051_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08133_, _08132_, _08057_);
  or (_08134_, _08133_, _08073_);
  or (_08135_, _08134_, _08130_);
  or (_08136_, _08135_, _08129_);
  or (_08137_, _08136_, _08128_);
  and (_26842_[6], _08137_, _22762_);
  not (_08138_, _07764_);
  and (_08139_, _08080_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_08140_, _07984_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_08141_, _08140_, _07782_);
  or (_08142_, _08141_, _08139_);
  or (_08143_, _08122_, _07577_);
  and (_08144_, _08143_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_08145_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_08146_, _07585_, _08145_);
  and (_08147_, _08146_, _07762_);
  or (_08148_, _08147_, _07763_);
  or (_08149_, _08148_, _08144_);
  or (_08150_, _08149_, _08142_);
  and (_08151_, _08150_, _08138_);
  and (_08152_, _08140_, _07570_);
  and (_08153_, _08053_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_08154_, _08147_, _08122_);
  or (_08155_, _08154_, _08153_);
  or (_08156_, _08155_, _08152_);
  or (_08157_, _08156_, _08151_);
  and (_08158_, _08157_, _08121_);
  and (_08159_, _08150_, _08050_);
  or (_08160_, _08139_, _08073_);
  or (_08163_, _08160_, _08104_);
  or (_08164_, _08163_, _08140_);
  or (_08165_, _08164_, _08159_);
  or (_08166_, _08165_, _08158_);
  and (_26842_[7], _08166_, _22762_);
  and (_08167_, _01809_, _24005_);
  and (_08168_, _08167_, _23946_);
  not (_08169_, _08167_);
  and (_08171_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or (_00995_, _08171_, _08168_);
  and (_08173_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  and (_08174_, _05199_, _23747_);
  or (_01020_, _08174_, _08173_);
  not (_08176_, _08058_);
  nor (_08177_, _07984_, _07951_);
  and (_08178_, _08177_, _07577_);
  or (_08180_, _08178_, _08176_);
  and (_08182_, _08180_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08184_, _07938_, _07577_);
  and (_08185_, _07762_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_08186_, _07764_, _07782_);
  and (_08187_, _08186_, _08185_);
  or (_08189_, _08104_, _07763_);
  or (_08191_, _08189_, _08187_);
  or (_08192_, _08191_, _08184_);
  or (_08193_, _08192_, _08122_);
  or (_08194_, _08193_, _08182_);
  and (_26842_[8], _08194_, _22762_);
  and (_08196_, _06602_, _23778_);
  and (_08197_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  or (_01104_, _08197_, _08196_);
  and (_08198_, _23903_, _23664_);
  and (_08199_, _08198_, _23898_);
  not (_08200_, _08198_);
  and (_08201_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_01130_, _08201_, _08199_);
  and (_08204_, _07880_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08206_, _07760_, _07940_);
  and (_08207_, _07992_, _07790_);
  nor (_08209_, _07880_, _07621_);
  or (_08211_, _08209_, _08207_);
  and (_08212_, _08211_, _08206_);
  or (_08213_, _08212_, _08184_);
  and (_08214_, _07608_, _07648_);
  and (_08216_, _08211_, _08050_);
  or (_08217_, _08216_, _08214_);
  or (_08218_, _08217_, _08213_);
  or (_08219_, _08218_, _08204_);
  and (_26842_[9], _08219_, _22762_);
  and (_08220_, _07947_, _07751_);
  not (_08222_, _07756_);
  and (_08223_, _08222_, _07655_);
  or (_08224_, _08223_, _08220_);
  not (_08225_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_08226_, _08040_, _08225_);
  and (_08227_, _07878_, _07648_);
  and (_08228_, _08227_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08229_, _08122_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08230_, _08229_, _07763_);
  or (_08231_, _08230_, _08228_);
  or (_08232_, _08231_, _08226_);
  or (_08233_, _08232_, _08207_);
  or (_08234_, _08233_, _08224_);
  or (_08235_, _08234_, _08184_);
  and (_26842_[10], _08235_, _22762_);
  and (_08236_, _08198_, _23778_);
  and (_08237_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or (_01277_, _08237_, _08236_);
  and (_08238_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and (_08239_, _05193_, _23898_);
  or (_01285_, _08239_, _08238_);
  and (_08241_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  and (_08242_, _05193_, _23778_);
  or (_01296_, _08242_, _08241_);
  nor (_08243_, _24628_, rst);
  and (_26888_, _08243_, _00289_);
  and (_08244_, _07947_, _07754_);
  and (_08245_, _08000_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08246_, _08245_, _08244_);
  and (_08247_, _07845_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08248_, _08080_, _07763_);
  and (_08249_, _08248_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08250_, _07812_, _07984_);
  and (_08251_, _08250_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08252_, _08251_, _08184_);
  or (_08253_, _08252_, _08249_);
  or (_08254_, _08253_, _08220_);
  or (_08255_, _08254_, _08247_);
  or (_08256_, _08255_, _08207_);
  or (_08257_, _08256_, _08246_);
  and (_26842_[11], _08257_, _22762_);
  and (_08259_, _02359_, _23707_);
  and (_08260_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  or (_01344_, _08260_, _08259_);
  and (_08261_, _08198_, _23649_);
  and (_08262_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_01348_, _08262_, _08261_);
  and (_08263_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  and (_08264_, _05193_, _23649_);
  or (_27228_, _08264_, _08263_);
  and (_08265_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and (_08266_, _04761_, _23898_);
  or (_01372_, _08266_, _08265_);
  and (_08267_, _08000_, _07782_);
  and (_08268_, _08267_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08269_, _07597_, _07648_);
  and (_08270_, _08269_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nand (_08271_, _08040_, _07940_);
  and (_08272_, _08271_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08273_, _07762_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_08274_, _08273_, _07992_);
  or (_08275_, _08274_, _08272_);
  or (_08276_, _08275_, _08270_);
  or (_08277_, _08276_, _08268_);
  and (_26842_[12], _08277_, _22762_);
  and (_08278_, _04333_, _24654_);
  nand (_08279_, _08278_, _23594_);
  or (_08280_, _08278_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_08281_, _08280_, _04339_);
  and (_08282_, _08281_, _08279_);
  nor (_08283_, _04339_, _23702_);
  or (_08284_, _08283_, _08282_);
  and (_01382_, _08284_, _22762_);
  or (_08285_, _04805_, _04725_);
  and (_08286_, _08285_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_08287_, _08286_, _04768_);
  and (_01384_, _08287_, _22762_);
  nor (_01386_, _06776_, rst);
  and (_08288_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  and (_08289_, _05193_, _23747_);
  or (_01393_, _08289_, _08288_);
  and (_08290_, _08198_, _23747_);
  and (_08291_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_01396_, _08291_, _08290_);
  and (_08292_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_08293_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_01407_, _08293_, _08292_);
  or (_08294_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_08295_, _08294_, _22762_);
  and (_08296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or (_08297_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_08298_, _08297_, rxd_i);
  or (_08299_, _08298_, _08296_);
  and (_08300_, _08299_, _04589_);
  and (_08301_, _04612_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_08302_, _08301_, _08300_);
  and (_08303_, _04602_, rxd_i);
  or (_08304_, _08303_, _04609_);
  or (_08305_, _08304_, _08302_);
  and (_01419_, _08305_, _08295_);
  or (_08306_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_08307_, _00273_, _24729_);
  or (_08308_, _08307_, _08306_);
  nand (_08309_, _05838_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_08310_, _08309_, _08307_);
  or (_08311_, _08310_, _05839_);
  and (_08312_, _08311_, _08308_);
  and (_08313_, _01975_, _24735_);
  or (_08314_, _08313_, _08312_);
  nand (_08315_, _08313_, _23702_);
  and (_08316_, _08315_, _22762_);
  and (_01438_, _08316_, _08314_);
  or (_08317_, _08053_, _07763_);
  or (_08318_, _08057_, _08122_);
  or (_08319_, _08318_, _08317_);
  or (_08320_, _08319_, _07879_);
  and (_08321_, _08320_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_08322_, _07597_, _07577_);
  or (_08323_, _08027_, _08322_);
  nor (_08324_, _08000_, _07572_);
  or (_08325_, _08324_, _08267_);
  and (_08326_, _08325_, _07586_);
  or (_08327_, _08326_, _08323_);
  or (_08328_, _08327_, _08321_);
  and (_26842_[13], _08328_, _22762_);
  and (_08329_, _04743_, _04582_);
  and (_08330_, _04727_, _08329_);
  nand (_08331_, _08330_, _04770_);
  or (_08332_, _08330_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_08333_, _08332_, _22762_);
  and (_01452_, _08333_, _08331_);
  or (_08334_, _06845_, rxd_i);
  nand (_08335_, _08334_, _04595_);
  or (_08336_, _04596_, _04578_);
  and (_08337_, _08336_, _08335_);
  or (_08338_, _04601_, _04579_);
  or (_08339_, _08338_, _04594_);
  or (_08340_, _08339_, _08337_);
  and (_01455_, _08340_, _02066_);
  or (_08341_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_08342_, _08341_, _22762_);
  nand (_08343_, _02034_, _23702_);
  and (_01457_, _08343_, _08342_);
  nand (_08344_, _04454_, _04449_);
  and (_08345_, _08344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_08346_, _08345_, _06799_);
  nor (_08347_, _04448_, _06800_);
  and (_08348_, _08347_, _08346_);
  or (_08349_, _08348_, _04569_);
  nand (_08350_, _08349_, _22762_);
  nor (_01466_, _08350_, _04462_);
  and (_08351_, _24201_, _24010_);
  not (_08352_, _08351_);
  and (_08353_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and (_08354_, _08351_, _23747_);
  or (_01495_, _08354_, _08353_);
  or (_08355_, _07860_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_26842_[14], _08355_, _22762_);
  and (_08356_, _23665_, _23649_);
  and (_08357_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  or (_01521_, _08357_, _08356_);
  and (_08358_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and (_08359_, _08351_, _23824_);
  or (_01524_, _08359_, _08358_);
  and (_08360_, _24005_, _23664_);
  and (_08361_, _08360_, _23747_);
  not (_08362_, _08360_);
  and (_08363_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  or (_01538_, _08363_, _08361_);
  and (_08364_, _08360_, _23824_);
  and (_08366_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  or (_01542_, _08366_, _08364_);
  and (_08367_, _23747_, _23665_);
  and (_08368_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  or (_27078_, _08368_, _08367_);
  and (_08369_, _05410_, _23824_);
  and (_08370_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  or (_01566_, _08370_, _08369_);
  and (_08371_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_08372_, _06896_, _24050_);
  or (_27022_, _08372_, _08371_);
  and (_08373_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_08374_, _06896_, _23707_);
  or (_01690_, _08374_, _08373_);
  and (_08375_, _24766_, _23911_);
  not (_08376_, _08375_);
  and (_08377_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and (_08378_, _08375_, _23898_);
  or (_01694_, _08378_, _08377_);
  and (_08379_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  and (_08381_, _08375_, _23747_);
  or (_01696_, _08381_, _08379_);
  and (_08382_, _02359_, _23898_);
  and (_08383_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  or (_01750_, _08383_, _08382_);
  and (_08384_, _02326_, _23898_);
  and (_08385_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_01761_, _08385_, _08384_);
  and (_08386_, _02326_, _23649_);
  and (_08387_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_01780_, _08387_, _08386_);
  and (_08388_, _02345_, _23946_);
  and (_08389_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_01784_, _08389_, _08388_);
  and (_08390_, _02359_, _23946_);
  and (_08391_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  or (_01789_, _08391_, _08390_);
  and (_08392_, _08010_, _08050_);
  not (_08393_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_08394_, _08015_, _07585_);
  nor (_08396_, _08394_, _08013_);
  and (_08397_, _08015_, _08058_);
  not (_08398_, _08397_);
  and (_08399_, _08398_, _08396_);
  and (_08400_, _08399_, _08015_);
  nor (_08401_, _08400_, _08393_);
  and (_08402_, _08015_, word_in[0]);
  and (_08403_, _08402_, _08399_);
  or (_08404_, _08403_, _08401_);
  or (_08405_, _08404_, _08392_);
  and (_08406_, _08000_, _07751_);
  and (_08407_, _08006_, _08406_);
  not (_08408_, _08407_);
  not (_08409_, _08392_);
  or (_08410_, _08409_, word_in[8]);
  and (_08411_, _08410_, _08408_);
  and (_08412_, _08411_, _08405_);
  and (_08413_, _07790_, _08000_);
  and (_08414_, _08028_, _08413_);
  and (_08415_, _08407_, word_in[16]);
  or (_08417_, _08415_, _08414_);
  or (_08418_, _08417_, _08412_);
  not (_08419_, _08414_);
  or (_08420_, _08419_, word_in[24]);
  and (_26843_[0], _08420_, _08418_);
  and (_08422_, _08006_, word_in[17]);
  and (_08423_, _08422_, _08406_);
  not (_08425_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_08426_, _08400_, _08425_);
  and (_08428_, _08015_, word_in[1]);
  and (_08430_, _08428_, _08399_);
  or (_08431_, _08430_, _08426_);
  and (_08433_, _08431_, _08409_);
  and (_08434_, _08392_, word_in[9]);
  or (_08436_, _08434_, _08433_);
  and (_08437_, _08436_, _08408_);
  or (_08438_, _08437_, _08423_);
  and (_08440_, _08438_, _08419_);
  and (_08441_, _08414_, word_in[25]);
  or (_26843_[1], _08441_, _08440_);
  and (_08443_, _02359_, _23747_);
  and (_08444_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  or (_01806_, _08444_, _08443_);
  and (_08445_, _08407_, word_in[18]);
  or (_08446_, _08409_, word_in[10]);
  and (_08447_, _08446_, _08408_);
  and (_08448_, _08400_, word_in[2]);
  not (_08450_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_08452_, _08400_, _08450_);
  or (_08453_, _08452_, _08448_);
  or (_08455_, _08453_, _08392_);
  and (_08456_, _08455_, _08447_);
  or (_08457_, _08456_, _08445_);
  and (_08459_, _08457_, _08419_);
  and (_08460_, _08414_, word_in[26]);
  or (_26843_[2], _08460_, _08459_);
  and (_08461_, _08028_, word_in[27]);
  and (_08462_, _08461_, _08413_);
  or (_08464_, _08409_, word_in[11]);
  and (_08465_, _08464_, _08408_);
  not (_08467_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_08468_, _08400_, _08467_);
  and (_08469_, _08400_, word_in[3]);
  or (_08470_, _08469_, _08468_);
  or (_08471_, _08470_, _08392_);
  and (_08472_, _08471_, _08465_);
  and (_08473_, _08407_, word_in[19]);
  or (_08474_, _08473_, _08472_);
  and (_08475_, _08474_, _08419_);
  or (_26843_[3], _08475_, _08462_);
  and (_08477_, _06506_, _23911_);
  not (_08478_, _08477_);
  and (_08479_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  and (_08480_, _08477_, _23707_);
  or (_26980_, _08480_, _08479_);
  and (_08481_, _08028_, word_in[28]);
  and (_08482_, _08481_, _08413_);
  or (_08483_, _08409_, word_in[12]);
  and (_08484_, _08483_, _08408_);
  not (_08485_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_08486_, _08400_, _08485_);
  and (_08488_, _08400_, word_in[4]);
  or (_08489_, _08488_, _08486_);
  or (_08490_, _08489_, _08392_);
  and (_08491_, _08490_, _08484_);
  and (_08492_, _08407_, word_in[20]);
  or (_08493_, _08492_, _08491_);
  and (_08494_, _08493_, _08419_);
  or (_26843_[4], _08494_, _08482_);
  and (_08495_, _08028_, word_in[29]);
  and (_08497_, _08495_, _08413_);
  and (_08498_, _08407_, word_in[21]);
  not (_08499_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_08500_, _08400_, _08499_);
  and (_08501_, _08015_, word_in[5]);
  and (_08502_, _08501_, _08400_);
  or (_08503_, _08502_, _08500_);
  or (_08504_, _08503_, _08392_);
  or (_08505_, _08409_, word_in[13]);
  and (_08506_, _08505_, _08408_);
  and (_08507_, _08506_, _08504_);
  or (_08508_, _08507_, _08498_);
  and (_08509_, _08508_, _08419_);
  or (_26843_[5], _08509_, _08497_);
  and (_08510_, _08028_, word_in[30]);
  and (_08511_, _08510_, _08413_);
  and (_08512_, _08407_, word_in[22]);
  or (_08513_, _08409_, word_in[14]);
  and (_08514_, _08513_, _08408_);
  not (_08515_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_08516_, _08400_, _08515_);
  and (_08517_, _08400_, word_in[6]);
  or (_08518_, _08517_, _08516_);
  or (_08519_, _08518_, _08392_);
  and (_08520_, _08519_, _08514_);
  or (_08521_, _08520_, _08512_);
  and (_08523_, _08521_, _08419_);
  or (_26843_[6], _08523_, _08511_);
  and (_08524_, _05410_, _23898_);
  and (_08525_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  or (_01820_, _08525_, _08524_);
  or (_08527_, _08409_, word_in[15]);
  and (_08528_, _08527_, _08408_);
  nor (_08529_, _08400_, _07837_);
  and (_08530_, _08400_, word_in[7]);
  or (_08531_, _08530_, _08529_);
  or (_08532_, _08531_, _08392_);
  and (_08533_, _08532_, _08528_);
  and (_08534_, _08407_, word_in[23]);
  or (_08535_, _08534_, _08533_);
  and (_08536_, _08535_, _08419_);
  and (_08537_, _08414_, word_in[31]);
  or (_26843_[7], _08537_, _08536_);
  and (_08539_, _06602_, _23747_);
  and (_08540_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  or (_01833_, _08540_, _08539_);
  and (_08541_, _06602_, _23707_);
  and (_08542_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  or (_01837_, _08542_, _08541_);
  and (_08543_, _06602_, _24050_);
  and (_08545_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  or (_27157_, _08545_, _08543_);
  and (_08546_, _05042_, _24050_);
  and (_08547_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_01860_, _08547_, _08546_);
  and (_08548_, _01809_, _24275_);
  and (_08549_, _08548_, _23747_);
  not (_08550_, _08548_);
  and (_08551_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or (_01866_, _08551_, _08549_);
  and (_08552_, _08028_, _08406_);
  and (_08553_, _08010_, _07780_);
  and (_08554_, _08553_, _07766_);
  not (_08555_, _08554_);
  not (_08556_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_08557_, _08013_, _07586_);
  and (_08558_, _08557_, _08398_);
  nor (_08559_, _08558_, _08556_);
  and (_08560_, _08558_, _08402_);
  or (_08561_, _08560_, _08559_);
  and (_08562_, _08561_, _08555_);
  and (_08563_, _08006_, _07754_);
  and (_08564_, _08563_, _07882_);
  and (_08565_, _08554_, word_in[8]);
  or (_08566_, _08565_, _08564_);
  or (_08567_, _08566_, _08562_);
  not (_08568_, _08564_);
  or (_08569_, _08568_, word_in[16]);
  and (_08570_, _08569_, _08567_);
  or (_08571_, _08570_, _08552_);
  not (_08573_, _08552_);
  or (_08574_, _08573_, word_in[24]);
  and (_26850_[0], _08574_, _08571_);
  not (_08575_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_08576_, _08558_, _08575_);
  and (_08577_, _08558_, _08428_);
  or (_08578_, _08577_, _08576_);
  and (_08579_, _08578_, _08555_);
  and (_08580_, _08554_, word_in[9]);
  or (_08581_, _08580_, _08564_);
  or (_08582_, _08581_, _08579_);
  or (_08583_, _08568_, word_in[17]);
  and (_08584_, _08583_, _08582_);
  or (_08585_, _08584_, _08552_);
  or (_08586_, _08573_, word_in[25]);
  and (_26850_[1], _08586_, _08585_);
  and (_08587_, _08548_, _23707_);
  and (_08588_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or (_01878_, _08588_, _08587_);
  not (_08589_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_08590_, _08558_, _08589_);
  and (_08591_, _08015_, word_in[2]);
  and (_08592_, _08558_, _08591_);
  or (_08593_, _08592_, _08590_);
  and (_08594_, _08593_, _08555_);
  and (_08595_, _08554_, word_in[10]);
  or (_08596_, _08595_, _08564_);
  or (_08597_, _08596_, _08594_);
  or (_08598_, _08568_, word_in[18]);
  and (_08599_, _08598_, _08597_);
  or (_08600_, _08599_, _08552_);
  or (_08601_, _08573_, word_in[26]);
  and (_26850_[2], _08601_, _08600_);
  not (_08602_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_08603_, _08558_, _08602_);
  and (_08604_, _08015_, word_in[3]);
  and (_08605_, _08558_, _08604_);
  or (_08606_, _08605_, _08603_);
  and (_08607_, _08606_, _08555_);
  and (_08608_, _08554_, word_in[11]);
  or (_08609_, _08608_, _08564_);
  or (_08610_, _08609_, _08607_);
  or (_08611_, _08568_, word_in[19]);
  and (_08612_, _08611_, _08610_);
  or (_08613_, _08612_, _08552_);
  or (_08614_, _08573_, word_in[27]);
  and (_26850_[3], _08614_, _08613_);
  and (_08615_, _08548_, _23946_);
  and (_08616_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or (_01881_, _08616_, _08615_);
  not (_08617_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_08618_, _08558_, _08617_);
  and (_08619_, _08015_, word_in[4]);
  and (_08620_, _08558_, _08619_);
  or (_08621_, _08620_, _08618_);
  and (_08622_, _08621_, _08555_);
  and (_08623_, _08554_, word_in[12]);
  or (_08624_, _08623_, _08564_);
  or (_08625_, _08624_, _08622_);
  or (_08626_, _08568_, word_in[20]);
  and (_08627_, _08626_, _08625_);
  or (_08628_, _08627_, _08552_);
  or (_08629_, _08573_, word_in[28]);
  and (_26850_[4], _08629_, _08628_);
  not (_08630_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_08631_, _08558_, _08630_);
  and (_08632_, _08558_, _08501_);
  or (_08633_, _08632_, _08631_);
  and (_08634_, _08633_, _08555_);
  and (_08635_, _08554_, word_in[13]);
  or (_08636_, _08635_, _08564_);
  or (_08637_, _08636_, _08634_);
  or (_08638_, _08568_, word_in[21]);
  and (_08639_, _08638_, _08637_);
  or (_08640_, _08639_, _08552_);
  or (_08641_, _08573_, word_in[29]);
  and (_26850_[5], _08641_, _08640_);
  and (_08642_, _02325_, _23784_);
  and (_08643_, _08642_, _23946_);
  not (_08644_, _08642_);
  and (_08645_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  or (_01885_, _08645_, _08643_);
  not (_08646_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_08647_, _08558_, _08646_);
  and (_08648_, _08015_, word_in[6]);
  and (_08649_, _08558_, _08648_);
  or (_08650_, _08649_, _08647_);
  and (_08651_, _08650_, _08555_);
  and (_08652_, _08554_, word_in[14]);
  or (_08653_, _08652_, _08564_);
  or (_08654_, _08653_, _08651_);
  or (_08655_, _08568_, word_in[22]);
  and (_08656_, _08655_, _08654_);
  or (_08657_, _08656_, _08552_);
  or (_08658_, _08573_, word_in[30]);
  and (_26850_[6], _08658_, _08657_);
  nor (_08659_, _08558_, _07675_);
  and (_08660_, _08558_, _08019_);
  or (_08661_, _08660_, _08659_);
  and (_08662_, _08661_, _08555_);
  and (_08663_, _08554_, word_in[15]);
  or (_08664_, _08663_, _08564_);
  or (_08665_, _08664_, _08662_);
  or (_08666_, _08568_, word_in[23]);
  and (_08667_, _08666_, _08665_);
  or (_08668_, _08667_, _08552_);
  or (_08669_, _08573_, word_in[31]);
  and (_26850_[7], _08669_, _08668_);
  and (_08670_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  and (_08671_, _08477_, _24050_);
  or (_01901_, _08671_, _08670_);
  and (_08673_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and (_08674_, _07513_, _23707_);
  or (_01928_, _08674_, _08673_);
  and (_08675_, _06544_, _23747_);
  and (_08676_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_01933_, _08676_, _08675_);
  and (_08677_, _08028_, _08050_);
  and (_08678_, _08006_, word_in[16]);
  and (_08679_, _08006_, _07780_);
  and (_08680_, _08679_, _07882_);
  not (_08681_, _08680_);
  or (_08682_, _08681_, _08678_);
  and (_08683_, _08010_, _07790_);
  and (_08684_, _08683_, _07766_);
  not (_08685_, _08684_);
  not (_08686_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  not (_08687_, _08013_);
  and (_08688_, _08394_, _08687_);
  and (_08689_, _08688_, _08176_);
  nor (_08690_, _08689_, _08686_);
  and (_08691_, _08689_, _08402_);
  or (_08692_, _08691_, _08690_);
  and (_08693_, _08692_, _08685_);
  and (_08694_, _08684_, word_in[8]);
  or (_08695_, _08694_, _08680_);
  or (_08696_, _08695_, _08693_);
  and (_08697_, _08696_, _08682_);
  or (_08698_, _08697_, _08677_);
  not (_08699_, _08677_);
  or (_08700_, _08699_, word_in[24]);
  and (_26851_[0], _08700_, _08698_);
  or (_08701_, _08681_, _08422_);
  not (_08702_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_08703_, _08689_, _08702_);
  and (_08704_, _08689_, _08428_);
  or (_08705_, _08704_, _08703_);
  and (_08706_, _08705_, _08685_);
  and (_08707_, _08684_, word_in[9]);
  or (_08708_, _08707_, _08680_);
  or (_08709_, _08708_, _08706_);
  and (_08710_, _08709_, _08701_);
  or (_08711_, _08710_, _08677_);
  or (_08712_, _08699_, word_in[25]);
  and (_26851_[1], _08712_, _08711_);
  and (_08713_, _06544_, _23707_);
  and (_08714_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_01943_, _08714_, _08713_);
  and (_08715_, _08006_, word_in[18]);
  or (_08716_, _08681_, _08715_);
  not (_08717_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_08718_, _08689_, _08717_);
  and (_08719_, _08689_, _08591_);
  or (_08720_, _08719_, _08718_);
  and (_08721_, _08720_, _08685_);
  and (_08722_, _08684_, word_in[10]);
  or (_08723_, _08722_, _08680_);
  or (_08724_, _08723_, _08721_);
  and (_08725_, _08724_, _08716_);
  or (_08726_, _08725_, _08677_);
  or (_08727_, _08699_, word_in[26]);
  and (_26851_[2], _08727_, _08726_);
  and (_08728_, _08006_, word_in[19]);
  or (_08729_, _08681_, _08728_);
  not (_08730_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_08731_, _08689_, _08730_);
  and (_08732_, _08689_, _08604_);
  or (_08733_, _08732_, _08731_);
  and (_08734_, _08733_, _08685_);
  and (_08735_, _08684_, word_in[11]);
  or (_08736_, _08735_, _08680_);
  or (_08737_, _08736_, _08734_);
  and (_08738_, _08737_, _08729_);
  or (_08739_, _08738_, _08677_);
  or (_08741_, _08699_, word_in[27]);
  and (_26851_[3], _08741_, _08739_);
  and (_08742_, _06530_, _23946_);
  and (_08743_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  or (_01946_, _08743_, _08742_);
  and (_08744_, _08006_, word_in[20]);
  or (_08745_, _08681_, _08744_);
  not (_08746_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_08747_, _08689_, _08746_);
  and (_08748_, _08689_, _08619_);
  or (_08750_, _08748_, _08747_);
  and (_08751_, _08750_, _08685_);
  and (_08752_, _08684_, word_in[12]);
  or (_08753_, _08752_, _08680_);
  or (_08754_, _08753_, _08751_);
  and (_08755_, _08754_, _08745_);
  or (_08756_, _08755_, _08677_);
  or (_08757_, _08699_, word_in[28]);
  and (_26851_[4], _08757_, _08756_);
  and (_08758_, _08006_, word_in[21]);
  or (_08759_, _08681_, _08758_);
  not (_08760_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_08761_, _08689_, _08760_);
  and (_08762_, _08689_, _08501_);
  or (_08763_, _08762_, _08761_);
  and (_08764_, _08763_, _08685_);
  and (_08766_, _08684_, word_in[13]);
  or (_08767_, _08766_, _08680_);
  or (_08768_, _08767_, _08764_);
  and (_08769_, _08768_, _08759_);
  or (_08770_, _08769_, _08677_);
  or (_08772_, _08699_, word_in[29]);
  and (_26851_[5], _08772_, _08770_);
  and (_08774_, _08006_, word_in[22]);
  or (_08775_, _08681_, _08774_);
  not (_08776_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_08778_, _08689_, _08776_);
  and (_08779_, _08689_, _08648_);
  or (_08780_, _08779_, _08778_);
  and (_08781_, _08780_, _08685_);
  and (_08782_, _08684_, word_in[14]);
  or (_08783_, _08782_, _08680_);
  or (_08784_, _08783_, _08781_);
  and (_08785_, _08784_, _08775_);
  or (_08786_, _08785_, _08677_);
  or (_08787_, _08699_, word_in[30]);
  and (_26851_[6], _08787_, _08786_);
  or (_08788_, _08681_, _08033_);
  nor (_08789_, _08689_, _07829_);
  and (_08790_, _08689_, _08019_);
  or (_08791_, _08790_, _08789_);
  and (_08792_, _08791_, _08685_);
  and (_08793_, _08684_, word_in[15]);
  or (_08794_, _08793_, _08680_);
  or (_08795_, _08794_, _08792_);
  and (_08796_, _08795_, _08788_);
  or (_08797_, _08796_, _08677_);
  or (_08798_, _08699_, word_in[31]);
  and (_26851_[7], _08798_, _08797_);
  and (_08799_, _25078_, _23664_);
  and (_08800_, _08799_, _23898_);
  not (_08801_, _08799_);
  and (_08802_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  or (_27077_, _08802_, _08800_);
  and (_08803_, _06517_, _23946_);
  and (_08804_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_01976_, _08804_, _08803_);
  and (_08805_, _06651_, _23649_);
  and (_08806_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  or (_01991_, _08806_, _08805_);
  and (_08807_, _08011_, _07766_);
  not (_08808_, _08807_);
  not (_08809_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_08810_, _08398_, _08014_);
  nor (_08811_, _08810_, _08809_);
  and (_08812_, _08810_, _08402_);
  or (_08813_, _08812_, _08811_);
  and (_08814_, _08813_, _08808_);
  and (_08815_, _08006_, _07790_);
  and (_08816_, _08815_, _07882_);
  and (_08817_, _08807_, word_in[8]);
  or (_08818_, _08817_, _08816_);
  or (_08819_, _08818_, _08814_);
  and (_08820_, _08028_, _08080_);
  not (_08821_, _08820_);
  not (_08822_, _08816_);
  or (_08823_, _08822_, _08678_);
  and (_08824_, _08823_, _08821_);
  and (_08825_, _08824_, _08819_);
  and (_08827_, _08820_, word_in[24]);
  or (_26852_[0], _08827_, _08825_);
  and (_08829_, _08820_, word_in[25]);
  not (_08830_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_08831_, _08810_, _08830_);
  and (_08832_, _08810_, _08428_);
  or (_08833_, _08832_, _08831_);
  and (_08834_, _08833_, _08808_);
  and (_08835_, _08807_, word_in[9]);
  or (_08836_, _08835_, _08816_);
  or (_08837_, _08836_, _08834_);
  or (_08838_, _08822_, word_in[17]);
  and (_08839_, _08838_, _08821_);
  and (_08840_, _08839_, _08837_);
  or (_26852_[1], _08840_, _08829_);
  and (_08841_, _06755_, _23946_);
  and (_08842_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_02003_, _08842_, _08841_);
  and (_08843_, _08820_, word_in[26]);
  not (_08844_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_08845_, _08810_, _08844_);
  and (_08846_, _08810_, _08591_);
  or (_08847_, _08846_, _08845_);
  and (_08848_, _08847_, _08808_);
  and (_08849_, _08807_, word_in[10]);
  or (_08850_, _08849_, _08816_);
  or (_08851_, _08850_, _08848_);
  or (_08853_, _08822_, word_in[18]);
  and (_08854_, _08853_, _08821_);
  and (_08855_, _08854_, _08851_);
  or (_26852_[2], _08855_, _08843_);
  and (_08856_, _08820_, word_in[27]);
  not (_08857_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_08858_, _08810_, _08857_);
  and (_08859_, _08810_, _08604_);
  or (_08860_, _08859_, _08858_);
  and (_08861_, _08860_, _08808_);
  and (_08862_, _08807_, word_in[11]);
  or (_08863_, _08862_, _08816_);
  or (_08864_, _08863_, _08861_);
  or (_08865_, _08822_, word_in[19]);
  and (_08866_, _08865_, _08821_);
  and (_08867_, _08866_, _08864_);
  or (_26852_[3], _08867_, _08856_);
  and (_08868_, _06755_, _23747_);
  and (_08869_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_02008_, _08869_, _08868_);
  not (_08870_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_08871_, _08810_, _08870_);
  and (_08872_, _08810_, _08619_);
  or (_08873_, _08872_, _08871_);
  and (_08874_, _08873_, _08808_);
  and (_08875_, _08807_, word_in[12]);
  or (_08876_, _08875_, _08816_);
  or (_08877_, _08876_, _08874_);
  or (_08878_, _08822_, word_in[20]);
  and (_08879_, _08878_, _08821_);
  and (_08880_, _08879_, _08877_);
  and (_08881_, _08820_, word_in[28]);
  or (_26852_[4], _08881_, _08880_);
  not (_08883_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_08884_, _08810_, _08883_);
  and (_08885_, _08810_, _08501_);
  or (_08886_, _08885_, _08884_);
  and (_08887_, _08886_, _08808_);
  and (_08888_, _08807_, word_in[13]);
  or (_08889_, _08888_, _08816_);
  or (_08890_, _08889_, _08887_);
  or (_08891_, _08822_, _08758_);
  and (_08892_, _08891_, _08821_);
  and (_08893_, _08892_, _08890_);
  and (_08894_, _08820_, word_in[29]);
  or (_26852_[5], _08894_, _08893_);
  and (_08895_, _06646_, _23824_);
  and (_08896_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_02013_, _08896_, _08895_);
  and (_08897_, _08820_, word_in[30]);
  not (_08898_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_08899_, _08810_, _08898_);
  and (_08900_, _08810_, _08648_);
  or (_08901_, _08900_, _08899_);
  and (_08902_, _08901_, _08808_);
  and (_08903_, _08807_, word_in[14]);
  or (_08904_, _08903_, _08816_);
  or (_08905_, _08904_, _08902_);
  or (_08906_, _08822_, word_in[22]);
  and (_08907_, _08906_, _08821_);
  and (_08910_, _08907_, _08905_);
  or (_26852_[6], _08910_, _08897_);
  nor (_08911_, _08810_, _07696_);
  and (_08912_, _08810_, _08019_);
  or (_08913_, _08912_, _08911_);
  and (_08914_, _08913_, _08808_);
  and (_08915_, _08807_, word_in[15]);
  or (_08916_, _08915_, _08816_);
  or (_08917_, _08916_, _08914_);
  or (_08918_, _08822_, word_in[23]);
  and (_08919_, _08918_, _08821_);
  and (_08920_, _08919_, _08917_);
  and (_08921_, _08820_, word_in[31]);
  or (_26852_[7], _08921_, _08920_);
  and (_08922_, _06646_, _23946_);
  and (_08923_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_02033_, _08923_, _08922_);
  and (_08924_, _05710_, _23898_);
  and (_08925_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  or (_02062_, _08925_, _08924_);
  and (_08927_, _06639_, _23824_);
  and (_08928_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_02068_, _08928_, _08927_);
  and (_08929_, _08028_, _07942_);
  and (_08930_, _08929_, _07948_);
  and (_08932_, _08930_, _07790_);
  and (_08933_, _08006_, _08053_);
  not (_08934_, _08933_);
  or (_08935_, _08934_, word_in[16]);
  and (_08936_, _08010_, _08057_);
  not (_08937_, _08936_);
  not (_08938_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_08940_, _08015_, _07762_);
  and (_08941_, _08940_, _08396_);
  nor (_08942_, _08941_, _08938_);
  and (_08944_, _08941_, _08402_);
  or (_08945_, _08944_, _08942_);
  and (_08946_, _08945_, _08937_);
  and (_08948_, _08936_, word_in[8]);
  or (_08949_, _08948_, _08933_);
  or (_08950_, _08949_, _08946_);
  and (_08952_, _08950_, _08935_);
  or (_08953_, _08952_, _08932_);
  and (_08954_, _08028_, word_in[24]);
  not (_08955_, _08932_);
  or (_08956_, _08955_, _08954_);
  and (_26853_[0], _08956_, _08953_);
  not (_08957_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_08958_, _08941_, _08957_);
  and (_08960_, _08941_, word_in[1]);
  or (_08961_, _08960_, _08958_);
  and (_08962_, _08961_, _08937_);
  and (_08964_, _08936_, word_in[9]);
  or (_08966_, _08964_, _08962_);
  or (_08967_, _08966_, _08933_);
  nor (_08968_, _08934_, _08422_);
  nor (_08970_, _08968_, _08932_);
  and (_08972_, _08970_, _08967_);
  and (_08973_, _08028_, word_in[25]);
  and (_08974_, _08932_, _08973_);
  or (_26853_[1], _08974_, _08972_);
  and (_08976_, _06639_, _23707_);
  and (_08978_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_02085_, _08978_, _08976_);
  not (_08979_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_08980_, _08941_, _08979_);
  and (_08982_, _08941_, word_in[2]);
  or (_08984_, _08982_, _08980_);
  and (_08985_, _08984_, _08937_);
  and (_08986_, _08936_, word_in[10]);
  or (_08987_, _08986_, _08985_);
  and (_08989_, _08987_, _08934_);
  and (_08990_, _08933_, word_in[18]);
  or (_08991_, _08990_, _08989_);
  and (_08992_, _08991_, _08955_);
  and (_08993_, _08028_, word_in[26]);
  and (_08994_, _08932_, _08993_);
  or (_26853_[2], _08994_, _08992_);
  not (_08996_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_08997_, _08941_, _08996_);
  and (_08998_, _08941_, word_in[3]);
  or (_08999_, _08998_, _08997_);
  and (_09000_, _08999_, _08937_);
  and (_09001_, _08936_, word_in[11]);
  or (_09003_, _09001_, _09000_);
  or (_09004_, _09003_, _08933_);
  nor (_09005_, _08934_, _08728_);
  nor (_09006_, _09005_, _08932_);
  and (_09007_, _09006_, _09004_);
  and (_09008_, _08932_, _08461_);
  or (_26853_[3], _09008_, _09007_);
  or (_09012_, _08934_, word_in[20]);
  not (_09013_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_09015_, _08941_, _09013_);
  and (_09016_, _08941_, _08619_);
  or (_09017_, _09016_, _09015_);
  or (_09019_, _09017_, _08936_);
  or (_09020_, _08937_, word_in[12]);
  and (_09021_, _09020_, _09019_);
  or (_09023_, _09021_, _08933_);
  and (_09024_, _09023_, _09012_);
  or (_09026_, _09024_, _08932_);
  or (_09027_, _08955_, _08481_);
  and (_26853_[4], _09027_, _09026_);
  or (_09028_, _08934_, word_in[21]);
  not (_09029_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_09030_, _08941_, _09029_);
  and (_09031_, _08941_, _08501_);
  or (_09032_, _09031_, _09030_);
  or (_09033_, _09032_, _08936_);
  or (_09034_, _08937_, word_in[13]);
  and (_09036_, _09034_, _09033_);
  or (_09037_, _09036_, _08933_);
  and (_09039_, _09037_, _09028_);
  or (_09040_, _09039_, _08932_);
  or (_09041_, _08955_, _08495_);
  and (_26853_[5], _09041_, _09040_);
  or (_09042_, _08934_, word_in[22]);
  not (_09043_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_09044_, _08941_, _09043_);
  and (_09045_, _08941_, _08648_);
  or (_09046_, _09045_, _09044_);
  or (_09048_, _09046_, _08936_);
  or (_09050_, _08937_, word_in[14]);
  and (_09051_, _09050_, _09048_);
  or (_09052_, _09051_, _08933_);
  and (_09053_, _09052_, _09042_);
  or (_09054_, _09053_, _08932_);
  or (_09055_, _08955_, _08510_);
  and (_26853_[6], _09055_, _09054_);
  and (_09057_, _25748_, _23649_);
  and (_09058_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_02098_, _09058_, _09057_);
  nor (_09060_, _08941_, _07852_);
  and (_09062_, _08941_, word_in[7]);
  or (_09063_, _09062_, _09060_);
  and (_09064_, _09063_, _08937_);
  and (_09065_, _08936_, word_in[15]);
  or (_09066_, _09065_, _09064_);
  and (_09067_, _09066_, _08934_);
  and (_09068_, _08933_, word_in[23]);
  or (_09069_, _09068_, _09067_);
  and (_09070_, _09069_, _08955_);
  and (_09072_, _08028_, word_in[31]);
  and (_09073_, _08932_, _09072_);
  or (_26853_[7], _09073_, _09070_);
  and (_09076_, _08563_, _08227_);
  not (_09077_, _09076_);
  and (_09078_, _08553_, _07845_);
  not (_09080_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_09082_, _08940_, _08557_);
  nor (_09083_, _09082_, _09080_);
  and (_09084_, _09082_, word_in[0]);
  nor (_09085_, _09084_, _09083_);
  nor (_09087_, _09085_, _09078_);
  and (_09088_, _09078_, word_in[8]);
  or (_09089_, _09088_, _09087_);
  and (_09090_, _09089_, _09077_);
  and (_09091_, _08930_, _07751_);
  and (_09092_, _09076_, _08678_);
  or (_09093_, _09092_, _09091_);
  or (_09095_, _09093_, _09090_);
  not (_09096_, _09091_);
  or (_09097_, _09096_, word_in[24]);
  and (_26854_[0], _09097_, _09095_);
  not (_09098_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_09099_, _09082_, _09098_);
  and (_09100_, _09082_, word_in[1]);
  nor (_09102_, _09100_, _09099_);
  nor (_09103_, _09102_, _09078_);
  and (_09104_, _09078_, word_in[9]);
  or (_09105_, _09104_, _09103_);
  and (_09106_, _09105_, _09077_);
  and (_09107_, _09076_, _08422_);
  or (_09108_, _09107_, _09091_);
  or (_09109_, _09108_, _09106_);
  or (_09111_, _09096_, word_in[25]);
  and (_26854_[1], _09111_, _09109_);
  not (_09113_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_09115_, _09082_, _09113_);
  and (_09116_, _09082_, word_in[2]);
  nor (_09117_, _09116_, _09115_);
  nor (_09119_, _09117_, _09078_);
  and (_09120_, _09078_, word_in[10]);
  or (_09121_, _09120_, _09119_);
  and (_09122_, _09121_, _09077_);
  and (_09123_, _09076_, _08715_);
  or (_09124_, _09123_, _09091_);
  or (_09125_, _09124_, _09122_);
  or (_09126_, _09096_, word_in[26]);
  and (_26854_[2], _09126_, _09125_);
  not (_09128_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_09129_, _09082_, _09128_);
  and (_09130_, _09082_, word_in[3]);
  nor (_09131_, _09130_, _09129_);
  nor (_09132_, _09131_, _09078_);
  and (_09133_, _09078_, word_in[11]);
  or (_09134_, _09133_, _09132_);
  and (_09135_, _09134_, _09077_);
  and (_09136_, _09076_, _08728_);
  or (_09137_, _09136_, _09091_);
  or (_09138_, _09137_, _09135_);
  or (_09139_, _09096_, word_in[27]);
  and (_26854_[3], _09139_, _09138_);
  not (_09141_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_09142_, _09082_, _09141_);
  and (_09143_, _09082_, word_in[4]);
  nor (_09144_, _09143_, _09142_);
  nor (_09145_, _09144_, _09078_);
  and (_09146_, _09078_, word_in[12]);
  or (_09147_, _09146_, _09145_);
  and (_09148_, _09147_, _09077_);
  and (_09149_, _09076_, _08744_);
  or (_09150_, _09149_, _09091_);
  or (_09151_, _09150_, _09148_);
  or (_09152_, _09096_, word_in[28]);
  and (_26854_[4], _09152_, _09151_);
  not (_09153_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_09154_, _09082_, _09153_);
  and (_09155_, _09082_, word_in[5]);
  nor (_09157_, _09155_, _09154_);
  nor (_09158_, _09157_, _09078_);
  and (_09159_, _09078_, word_in[13]);
  or (_09160_, _09159_, _09158_);
  and (_09161_, _09160_, _09077_);
  and (_09162_, _09076_, _08758_);
  or (_09163_, _09162_, _09091_);
  or (_09164_, _09163_, _09161_);
  or (_09165_, _09096_, word_in[29]);
  and (_26854_[5], _09165_, _09164_);
  not (_09166_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_09168_, _09082_, _09166_);
  and (_09169_, _09082_, word_in[6]);
  nor (_09170_, _09169_, _09168_);
  nor (_09171_, _09170_, _09078_);
  and (_09173_, _09078_, word_in[14]);
  or (_09175_, _09173_, _09171_);
  and (_09176_, _09175_, _09077_);
  and (_09177_, _09076_, _08774_);
  or (_09178_, _09177_, _09091_);
  or (_09180_, _09178_, _09176_);
  or (_09181_, _09096_, word_in[30]);
  and (_26854_[6], _09181_, _09180_);
  or (_09182_, _09077_, _08033_);
  nor (_09183_, _09082_, _07689_);
  and (_09185_, _09082_, word_in[7]);
  or (_09186_, _09185_, _09183_);
  or (_09187_, _09186_, _09078_);
  not (_09188_, word_in[15]);
  nand (_09189_, _09078_, _09188_);
  and (_09192_, _09189_, _09187_);
  or (_09193_, _09192_, _09076_);
  and (_09195_, _09193_, _09182_);
  or (_09196_, _09195_, _09091_);
  or (_09197_, _09096_, word_in[31]);
  and (_26854_[7], _09197_, _09196_);
  and (_09198_, _08930_, _07754_);
  and (_09199_, _08683_, _07845_);
  not (_09200_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_09201_, _08940_, _08688_);
  nor (_09203_, _09201_, _09200_);
  and (_09204_, _09201_, _08402_);
  or (_09205_, _09204_, _09203_);
  or (_09207_, _09205_, _09199_);
  not (_09208_, _09199_);
  or (_09209_, _09208_, word_in[8]);
  and (_09210_, _09209_, _09207_);
  and (_09211_, _08007_, _07915_);
  and (_09212_, _09211_, _07780_);
  or (_09213_, _09212_, _09210_);
  not (_09214_, _09212_);
  or (_09216_, _09214_, _08678_);
  and (_09217_, _09216_, _09213_);
  or (_09218_, _09217_, _09198_);
  not (_09220_, _09198_);
  or (_09221_, _09220_, word_in[24]);
  and (_26855_[0], _09221_, _09218_);
  not (_09222_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_09223_, _09201_, _09222_);
  and (_09224_, _09201_, _08428_);
  or (_09226_, _09224_, _09223_);
  and (_09227_, _09226_, _09208_);
  and (_09229_, _09199_, word_in[9]);
  or (_09230_, _09229_, _09227_);
  or (_09231_, _09230_, _09212_);
  or (_09232_, _09214_, _08422_);
  and (_09233_, _09232_, _09231_);
  or (_09234_, _09233_, _09198_);
  or (_09235_, _09220_, word_in[25]);
  and (_26855_[1], _09235_, _09234_);
  not (_09236_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_09237_, _09201_, _09236_);
  and (_09238_, _09201_, _08591_);
  or (_09239_, _09238_, _09237_);
  or (_09240_, _09239_, _09199_);
  or (_09241_, _09208_, word_in[10]);
  and (_09242_, _09241_, _09240_);
  or (_09243_, _09242_, _09212_);
  or (_09244_, _09214_, _08715_);
  and (_09245_, _09244_, _09243_);
  or (_09246_, _09245_, _09198_);
  or (_09247_, _09220_, word_in[26]);
  and (_26855_[2], _09247_, _09246_);
  not (_09248_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_09249_, _09201_, _09248_);
  and (_09250_, _09201_, _08604_);
  or (_09251_, _09250_, _09249_);
  and (_09252_, _09251_, _09208_);
  and (_09253_, _09199_, word_in[11]);
  or (_09255_, _09253_, _09252_);
  or (_09256_, _09255_, _09212_);
  or (_09257_, _09214_, _08728_);
  and (_09259_, _09257_, _09256_);
  or (_09260_, _09259_, _09198_);
  or (_09261_, _09220_, word_in[27]);
  and (_26855_[3], _09261_, _09260_);
  not (_09262_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_09263_, _09201_, _09262_);
  and (_09264_, _09201_, _08619_);
  or (_09265_, _09264_, _09263_);
  or (_09266_, _09265_, _09199_);
  or (_09267_, _09208_, word_in[12]);
  and (_09268_, _09267_, _09266_);
  or (_09269_, _09268_, _09212_);
  or (_09271_, _09214_, _08744_);
  and (_09272_, _09271_, _09269_);
  or (_09273_, _09272_, _09198_);
  or (_09275_, _09220_, word_in[28]);
  and (_26855_[4], _09275_, _09273_);
  and (_09276_, _02345_, _23707_);
  and (_09278_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_02210_, _09278_, _09276_);
  not (_09279_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_09280_, _09201_, _09279_);
  and (_09281_, _09201_, _08501_);
  or (_09283_, _09281_, _09280_);
  or (_09284_, _09283_, _09199_);
  or (_09285_, _09208_, word_in[13]);
  and (_09286_, _09285_, _09284_);
  or (_09287_, _09286_, _09212_);
  nor (_09288_, _09214_, _08758_);
  nor (_09289_, _09288_, _09198_);
  and (_09290_, _09289_, _09287_);
  and (_09292_, _09198_, word_in[29]);
  or (_26855_[5], _09292_, _09290_);
  not (_09293_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_09294_, _09201_, _09293_);
  and (_09295_, _09201_, _08648_);
  or (_09297_, _09295_, _09294_);
  and (_09298_, _09297_, _09208_);
  and (_09300_, _09199_, word_in[14]);
  or (_09301_, _09300_, _09298_);
  or (_09303_, _09301_, _09212_);
  nor (_09304_, _09214_, _08774_);
  nor (_09306_, _09304_, _09198_);
  and (_09307_, _09306_, _09303_);
  and (_09308_, _09198_, word_in[30]);
  or (_26855_[6], _09308_, _09307_);
  nor (_09310_, _09201_, _07846_);
  and (_09311_, _09201_, _08019_);
  or (_09313_, _09311_, _09310_);
  or (_09314_, _09313_, _09199_);
  nand (_09316_, _09199_, _09188_);
  and (_09318_, _09316_, _09314_);
  or (_09319_, _09318_, _09212_);
  nor (_09320_, _09214_, _08033_);
  nor (_09322_, _09320_, _09198_);
  and (_09323_, _09322_, _09319_);
  and (_09324_, _09198_, word_in[31]);
  or (_26855_[7], _09324_, _09323_);
  and (_09325_, _08028_, _08073_);
  not (_09326_, _09325_);
  and (_09328_, _08227_, _08815_);
  and (_09329_, _09328_, _08678_);
  not (_09330_, _09328_);
  and (_09332_, _08011_, _07845_);
  not (_09333_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_09335_, _08940_, _08014_);
  nor (_09336_, _09335_, _09333_);
  and (_09337_, _09335_, word_in[0]);
  nor (_09339_, _09337_, _09336_);
  nor (_09341_, _09339_, _09332_);
  and (_09342_, _09332_, word_in[8]);
  or (_09344_, _09342_, _09341_);
  and (_09345_, _09344_, _09330_);
  or (_09346_, _09345_, _09329_);
  and (_09348_, _09346_, _09326_);
  and (_09349_, _09325_, word_in[24]);
  or (_26856_[0], _09349_, _09348_);
  and (_09351_, _09325_, _08973_);
  not (_09352_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_09353_, _09335_, _09352_);
  and (_09355_, _09335_, word_in[1]);
  nor (_09356_, _09355_, _09353_);
  nor (_09358_, _09356_, _09332_);
  and (_09360_, _09332_, word_in[9]);
  or (_09361_, _09360_, _09358_);
  and (_09362_, _09361_, _09330_);
  and (_09363_, _09328_, _08422_);
  or (_09364_, _09363_, _09362_);
  and (_09367_, _09364_, _09326_);
  or (_26856_[1], _09367_, _09351_);
  and (_09369_, _09328_, _08715_);
  not (_09371_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_09372_, _09335_, _09371_);
  and (_09374_, _09335_, word_in[2]);
  nor (_09376_, _09374_, _09372_);
  nor (_09377_, _09376_, _09332_);
  and (_09378_, _09332_, word_in[10]);
  or (_09380_, _09378_, _09377_);
  and (_09381_, _09380_, _09330_);
  or (_09383_, _09381_, _09369_);
  and (_09385_, _09383_, _09326_);
  and (_09386_, _09325_, word_in[26]);
  or (_26856_[2], _09386_, _09385_);
  and (_09388_, _09328_, _08728_);
  not (_09389_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_09390_, _09335_, _09389_);
  and (_09391_, _09335_, word_in[3]);
  nor (_09392_, _09391_, _09390_);
  nor (_09394_, _09392_, _09332_);
  and (_09395_, _09332_, word_in[11]);
  or (_09396_, _09395_, _09394_);
  and (_09397_, _09396_, _09330_);
  or (_09398_, _09397_, _09388_);
  and (_09399_, _09398_, _09326_);
  and (_09400_, _09325_, word_in[27]);
  or (_26856_[3], _09400_, _09399_);
  and (_09401_, _09328_, _08744_);
  not (_09402_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_09403_, _09335_, _09402_);
  and (_09404_, _09335_, word_in[4]);
  nor (_09405_, _09404_, _09403_);
  nor (_09406_, _09405_, _09332_);
  and (_09407_, _09332_, word_in[12]);
  or (_09408_, _09407_, _09406_);
  and (_09409_, _09408_, _09330_);
  or (_09410_, _09409_, _09401_);
  and (_09411_, _09410_, _09326_);
  and (_09412_, _09325_, word_in[28]);
  or (_26856_[4], _09412_, _09411_);
  and (_09414_, _09325_, _08495_);
  not (_09415_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_09416_, _09335_, _09415_);
  and (_09417_, _09335_, word_in[5]);
  nor (_09418_, _09417_, _09416_);
  nor (_09419_, _09418_, _09332_);
  and (_09420_, _09332_, word_in[13]);
  or (_09422_, _09420_, _09419_);
  and (_09423_, _09422_, _09330_);
  and (_09424_, _09328_, _08758_);
  or (_09425_, _09424_, _09423_);
  and (_09426_, _09425_, _09326_);
  or (_26856_[5], _09426_, _09414_);
  and (_09427_, _09328_, _08774_);
  not (_09428_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_09429_, _09335_, _09428_);
  and (_09430_, _09335_, word_in[6]);
  nor (_09431_, _09430_, _09429_);
  nor (_09432_, _09431_, _09332_);
  and (_09434_, _09332_, word_in[14]);
  or (_09435_, _09434_, _09432_);
  and (_09436_, _09435_, _09330_);
  or (_09437_, _09436_, _09427_);
  and (_09438_, _09437_, _09326_);
  and (_09439_, _09325_, word_in[30]);
  or (_26856_[6], _09439_, _09438_);
  and (_09440_, _09328_, _08033_);
  nor (_09441_, _09335_, _07682_);
  and (_09442_, _09335_, word_in[7]);
  nor (_09443_, _09442_, _09441_);
  nor (_09444_, _09443_, _09332_);
  and (_09445_, _09332_, word_in[15]);
  or (_09446_, _09445_, _09444_);
  and (_09447_, _09446_, _09330_);
  or (_09448_, _09447_, _09440_);
  and (_09449_, _09448_, _09326_);
  and (_09450_, _09325_, word_in[31]);
  or (_26856_[7], _09450_, _09449_);
  and (_09451_, _08006_, _08122_);
  and (_09452_, _08010_, _07763_);
  not (_09453_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nand (_09454_, _07761_, _07577_);
  not (_09455_, _09454_);
  and (_09456_, _08015_, _09455_);
  and (_09457_, _09456_, _08396_);
  nor (_09458_, _09457_, _09453_);
  and (_09459_, _09457_, _08402_);
  or (_09460_, _09459_, _09458_);
  or (_09461_, _09460_, _09452_);
  not (_09462_, _09452_);
  or (_09463_, _09462_, word_in[8]);
  and (_09464_, _09463_, _09461_);
  or (_09465_, _09464_, _09451_);
  and (_09466_, _08028_, _07951_);
  and (_09467_, _09466_, _07790_);
  not (_09468_, _09451_);
  nor (_09469_, _09468_, word_in[16]);
  nor (_09470_, _09469_, _09467_);
  and (_09471_, _09470_, _09465_);
  and (_09472_, _09467_, word_in[24]);
  or (_26857_[0], _09472_, _09471_);
  or (_09473_, _09468_, word_in[17]);
  not (_09474_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_09475_, _09457_, _09474_);
  and (_09476_, _09457_, _08428_);
  or (_09477_, _09476_, _09475_);
  or (_09478_, _09477_, _09452_);
  or (_09479_, _09462_, word_in[9]);
  and (_09480_, _09479_, _09478_);
  or (_09481_, _09480_, _09451_);
  and (_09482_, _09481_, _09473_);
  or (_09483_, _09482_, _09467_);
  not (_09484_, _09467_);
  or (_09485_, _09484_, word_in[25]);
  and (_26857_[1], _09485_, _09483_);
  not (_09486_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_09487_, _09457_, _09486_);
  and (_09488_, _09457_, word_in[2]);
  or (_09489_, _09488_, _09487_);
  and (_09491_, _09489_, _09462_);
  and (_09492_, _09452_, word_in[10]);
  or (_09493_, _09492_, _09491_);
  and (_09494_, _09493_, _09468_);
  and (_09495_, _09451_, word_in[18]);
  or (_09496_, _09495_, _09494_);
  and (_09497_, _09496_, _09484_);
  and (_09498_, _09467_, word_in[26]);
  or (_26857_[2], _09498_, _09497_);
  not (_09499_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_09500_, _09457_, _09499_);
  and (_09501_, _09457_, _08604_);
  or (_09502_, _09501_, _09500_);
  or (_09503_, _09502_, _09452_);
  or (_09504_, _09462_, word_in[11]);
  and (_09505_, _09504_, _09468_);
  and (_09506_, _09505_, _09503_);
  and (_09507_, _09451_, word_in[19]);
  or (_09508_, _09507_, _09506_);
  or (_09509_, _09508_, _09467_);
  or (_09510_, _09484_, word_in[27]);
  and (_26857_[3], _09510_, _09509_);
  or (_09511_, _09468_, word_in[20]);
  not (_09512_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_09513_, _09457_, _09512_);
  and (_09514_, _09457_, _08619_);
  or (_09515_, _09514_, _09513_);
  or (_09516_, _09515_, _09452_);
  or (_09517_, _09462_, word_in[12]);
  and (_09518_, _09517_, _09516_);
  or (_09520_, _09518_, _09451_);
  and (_09521_, _09520_, _09511_);
  or (_09522_, _09521_, _09467_);
  or (_09524_, _09484_, word_in[28]);
  and (_26857_[4], _09524_, _09522_);
  not (_09525_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_09526_, _09457_, _09525_);
  and (_09527_, _09457_, _08501_);
  or (_09528_, _09527_, _09526_);
  or (_09529_, _09528_, _09452_);
  or (_09530_, _09462_, word_in[13]);
  and (_09531_, _09530_, _09529_);
  or (_09532_, _09531_, _09451_);
  or (_09533_, _09468_, word_in[21]);
  and (_09534_, _09533_, _09532_);
  or (_09535_, _09534_, _09467_);
  or (_09536_, _09484_, word_in[29]);
  and (_26857_[5], _09536_, _09535_);
  not (_09537_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_09538_, _09457_, _09537_);
  and (_09539_, _09457_, _08648_);
  or (_09540_, _09539_, _09538_);
  or (_09541_, _09540_, _09452_);
  or (_09542_, _09462_, word_in[14]);
  and (_09543_, _09542_, _09541_);
  or (_09544_, _09543_, _09451_);
  nor (_09545_, _09468_, word_in[22]);
  nor (_09546_, _09545_, _09467_);
  and (_09547_, _09546_, _09544_);
  and (_09548_, _09467_, word_in[30]);
  or (_26857_[6], _09548_, _09547_);
  nor (_09549_, _09457_, _07819_);
  and (_09550_, _09457_, word_in[7]);
  or (_09551_, _09550_, _09549_);
  and (_09552_, _09551_, _09462_);
  and (_09553_, _09452_, word_in[15]);
  or (_09554_, _09553_, _09552_);
  or (_09555_, _09554_, _09451_);
  nor (_09556_, _09468_, word_in[23]);
  nor (_09557_, _09556_, _09467_);
  and (_09558_, _09557_, _09555_);
  and (_09559_, _09467_, word_in[31]);
  or (_26857_[7], _09559_, _09558_);
  nor (_26860_[7], _24508_, rst);
  and (_09560_, _08799_, _23747_);
  and (_09561_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or (_02338_, _09561_, _09560_);
  and (_09562_, _24371_, _23898_);
  and (_09563_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_27197_, _09563_, _09562_);
  nor (_26887_[7], _26770_, rst);
  and (_09564_, _08799_, _23824_);
  and (_09565_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  or (_02348_, _09565_, _09564_);
  nor (_26860_[5], _24530_, rst);
  and (_09566_, _08043_, _23898_);
  and (_09567_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_02362_, _09567_, _09566_);
  and (_09568_, _08563_, _07887_);
  and (_09569_, _08553_, _07770_);
  not (_09570_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_09571_, _09456_, _08557_);
  nor (_09572_, _09571_, _09570_);
  and (_09573_, _09571_, _08402_);
  or (_09574_, _09573_, _09572_);
  or (_09575_, _09574_, _09569_);
  not (_09576_, _09569_);
  or (_09577_, _09576_, word_in[8]);
  and (_09578_, _09577_, _09575_);
  or (_09579_, _09578_, _09568_);
  and (_09580_, _09466_, _07751_);
  not (_09581_, _09568_);
  nor (_09582_, _09581_, _08678_);
  nor (_09583_, _09582_, _09580_);
  and (_09584_, _09583_, _09579_);
  and (_09585_, _09580_, word_in[24]);
  or (_26858_[0], _09585_, _09584_);
  not (_09586_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_09587_, _09571_, _09586_);
  and (_09588_, _09571_, _08428_);
  or (_09589_, _09588_, _09587_);
  or (_09590_, _09589_, _09569_);
  or (_09591_, _09576_, word_in[9]);
  and (_09592_, _09591_, _09590_);
  or (_09593_, _09592_, _09568_);
  nor (_09594_, _09581_, _08422_);
  nor (_09595_, _09594_, _09580_);
  and (_09596_, _09595_, _09593_);
  and (_09597_, _09580_, word_in[25]);
  or (_26858_[1], _09597_, _09596_);
  not (_09598_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_09599_, _09571_, _09598_);
  and (_09601_, _09571_, _08591_);
  or (_09602_, _09601_, _09599_);
  or (_09603_, _09602_, _09569_);
  or (_09604_, _09576_, word_in[10]);
  and (_09605_, _09604_, _09603_);
  or (_09606_, _09605_, _09568_);
  nor (_09607_, _09581_, _08715_);
  nor (_09608_, _09607_, _09580_);
  and (_09610_, _09608_, _09606_);
  and (_09611_, _09580_, word_in[26]);
  or (_26858_[2], _09611_, _09610_);
  not (_09613_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_09614_, _09571_, _09613_);
  and (_09615_, _09571_, _08604_);
  or (_09616_, _09615_, _09614_);
  or (_09617_, _09616_, _09569_);
  or (_09618_, _09576_, word_in[11]);
  and (_09619_, _09618_, _09617_);
  or (_09620_, _09619_, _09568_);
  nor (_09621_, _09581_, _08728_);
  nor (_09622_, _09621_, _09580_);
  and (_09623_, _09622_, _09620_);
  and (_09624_, _09580_, word_in[27]);
  or (_26858_[3], _09624_, _09623_);
  not (_09625_, _09580_);
  not (_09627_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_09628_, _09571_, _09627_);
  and (_09629_, _09571_, _08619_);
  nor (_09630_, _09629_, _09628_);
  nor (_09631_, _09630_, _09569_);
  and (_09632_, _09569_, word_in[12]);
  or (_09633_, _09632_, _09568_);
  or (_09634_, _09633_, _09631_);
  or (_09635_, _09581_, _08744_);
  and (_09636_, _09635_, _09634_);
  and (_09637_, _09636_, _09625_);
  and (_09639_, _09580_, word_in[28]);
  or (_26858_[4], _09639_, _09637_);
  or (_09640_, _09581_, _08758_);
  not (_09641_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_09642_, _09571_, _09641_);
  and (_09643_, _09571_, _08501_);
  nor (_09644_, _09643_, _09642_);
  nor (_09645_, _09644_, _09569_);
  and (_09646_, _09569_, word_in[13]);
  or (_09647_, _09646_, _09568_);
  or (_09648_, _09647_, _09645_);
  and (_09649_, _09648_, _09640_);
  and (_09651_, _09649_, _09625_);
  and (_09653_, _09580_, word_in[29]);
  or (_26858_[5], _09653_, _09651_);
  not (_09654_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_09655_, _09571_, _09654_);
  and (_09656_, _09571_, _08648_);
  or (_09657_, _09656_, _09655_);
  or (_09658_, _09657_, _09569_);
  or (_09659_, _09576_, word_in[14]);
  and (_09660_, _09659_, _09658_);
  or (_09661_, _09660_, _09568_);
  nor (_09662_, _09581_, _08774_);
  nor (_09663_, _09662_, _09580_);
  and (_09664_, _09663_, _09661_);
  and (_09665_, _09580_, word_in[30]);
  or (_26858_[6], _09665_, _09664_);
  nor (_09666_, _09571_, _07709_);
  and (_09667_, _09571_, _08019_);
  or (_09669_, _09667_, _09666_);
  or (_09670_, _09669_, _09569_);
  nand (_09671_, _09569_, _09188_);
  and (_09672_, _09671_, _09670_);
  or (_09673_, _09672_, _09568_);
  nor (_09674_, _09581_, _08033_);
  nor (_09675_, _09674_, _09580_);
  and (_09676_, _09675_, _09673_);
  and (_09677_, _09580_, word_in[31]);
  or (_26858_[7], _09677_, _09676_);
  and (_09678_, _24371_, _23778_);
  and (_09679_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_27196_, _09679_, _09678_);
  and (_09682_, _09466_, _07754_);
  and (_09683_, _08679_, _07887_);
  not (_09684_, _09683_);
  or (_09685_, _09684_, _08678_);
  not (_09686_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_09687_, _08688_, _09455_);
  nor (_09688_, _09687_, _09686_);
  and (_09689_, _09687_, _08402_);
  or (_09690_, _09689_, _09688_);
  and (_09691_, _08010_, _07770_);
  and (_09692_, _09691_, _08683_);
  not (_09693_, _09692_);
  and (_09694_, _09693_, _09690_);
  and (_09695_, _08683_, _07770_);
  and (_09696_, _09695_, word_in[8]);
  or (_09697_, _09696_, _09683_);
  or (_09698_, _09697_, _09694_);
  and (_09699_, _09698_, _09685_);
  or (_09700_, _09699_, _09682_);
  not (_09701_, _09682_);
  or (_09702_, _09701_, word_in[24]);
  and (_26844_[0], _09702_, _09700_);
  not (_09703_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_09704_, _09687_, _09703_);
  and (_09705_, _09687_, _08428_);
  or (_09706_, _09705_, _09704_);
  or (_09707_, _09706_, _09695_);
  not (_09708_, _09695_);
  or (_09709_, _09708_, word_in[9]);
  and (_09710_, _09709_, _09707_);
  or (_09711_, _09710_, _09683_);
  nor (_09712_, _09684_, _08422_);
  nor (_09713_, _09712_, _09682_);
  and (_09714_, _09713_, _09711_);
  and (_09715_, _09682_, word_in[25]);
  or (_26844_[1], _09715_, _09714_);
  not (_09716_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_09717_, _09687_, _09716_);
  and (_09718_, _09687_, _08591_);
  or (_09719_, _09718_, _09717_);
  or (_09720_, _09719_, _09695_);
  or (_09721_, _09708_, word_in[10]);
  and (_09722_, _09721_, _09720_);
  or (_09723_, _09722_, _09683_);
  nor (_09724_, _09684_, _08715_);
  nor (_09725_, _09724_, _09682_);
  and (_09726_, _09725_, _09723_);
  and (_09727_, _09682_, word_in[26]);
  or (_26844_[2], _09727_, _09726_);
  and (_09729_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and (_09730_, _08351_, _24050_);
  or (_02446_, _09730_, _09729_);
  not (_09732_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_09734_, _09687_, _09732_);
  and (_09735_, _09687_, _08604_);
  or (_09736_, _09735_, _09734_);
  or (_09738_, _09736_, _09695_);
  or (_09739_, _09708_, word_in[11]);
  and (_09740_, _09739_, _09738_);
  or (_09741_, _09740_, _09683_);
  nor (_09742_, _09684_, _08728_);
  nor (_09743_, _09742_, _09682_);
  and (_09744_, _09743_, _09741_);
  and (_09745_, _09682_, word_in[27]);
  or (_26844_[3], _09745_, _09744_);
  not (_09746_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_09747_, _09687_, _09746_);
  and (_09748_, _09687_, _08619_);
  or (_09749_, _09748_, _09747_);
  or (_09751_, _09749_, _09695_);
  or (_09752_, _09708_, word_in[12]);
  and (_09754_, _09752_, _09751_);
  or (_09755_, _09754_, _09683_);
  nor (_09756_, _09684_, _08744_);
  nor (_09757_, _09756_, _09682_);
  and (_09758_, _09757_, _09755_);
  and (_09759_, _09682_, word_in[28]);
  or (_26844_[4], _09759_, _09758_);
  not (_09760_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_09761_, _09687_, _09760_);
  and (_09762_, _09687_, _08501_);
  or (_09763_, _09762_, _09761_);
  or (_09764_, _09763_, _09695_);
  or (_09765_, _09708_, word_in[13]);
  and (_09766_, _09765_, _09764_);
  or (_09767_, _09766_, _09683_);
  nor (_09768_, _09684_, _08758_);
  nor (_09770_, _09768_, _09682_);
  and (_09771_, _09770_, _09767_);
  and (_09773_, _09682_, word_in[29]);
  or (_26844_[5], _09773_, _09771_);
  not (_09774_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_09775_, _09687_, _09774_);
  and (_09776_, _09687_, _08648_);
  or (_09777_, _09776_, _09775_);
  or (_09778_, _09777_, _09695_);
  or (_09779_, _09708_, word_in[14]);
  and (_09780_, _09779_, _09778_);
  or (_09781_, _09780_, _09683_);
  nor (_09782_, _09684_, _08774_);
  nor (_09783_, _09782_, _09682_);
  and (_09784_, _09783_, _09781_);
  and (_09785_, _09682_, word_in[30]);
  or (_26844_[6], _09785_, _09784_);
  or (_09786_, _09684_, _08033_);
  nor (_09787_, _09687_, _07813_);
  and (_09788_, _09687_, _08019_);
  or (_09789_, _09788_, _09787_);
  and (_09790_, _09789_, _09693_);
  and (_09792_, _09695_, word_in[15]);
  or (_09793_, _09792_, _09683_);
  or (_09794_, _09793_, _09790_);
  and (_09795_, _09794_, _09786_);
  or (_09796_, _09795_, _09682_);
  or (_09797_, _09701_, word_in[31]);
  and (_26844_[7], _09797_, _09796_);
  and (_09798_, _08043_, _23778_);
  and (_09799_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_27210_, _09799_, _09798_);
  and (_09800_, _09466_, _07780_);
  and (_09801_, _08011_, _07770_);
  not (_09802_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_09803_, _09456_, _08014_);
  nor (_09804_, _09803_, _09802_);
  and (_09805_, _09803_, _08402_);
  nor (_09806_, _09805_, _09804_);
  nor (_09807_, _09806_, _09801_);
  and (_09808_, _08815_, _07887_);
  and (_09809_, _09801_, word_in[8]);
  or (_09810_, _09809_, _09808_);
  or (_09811_, _09810_, _09807_);
  not (_09812_, _09808_);
  or (_09813_, _09812_, _08678_);
  and (_09814_, _09813_, _09811_);
  or (_09815_, _09814_, _09800_);
  not (_09816_, _09800_);
  or (_09817_, _09816_, word_in[24]);
  and (_26845_[0], _09817_, _09815_);
  not (_09819_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_09820_, _09803_, _09819_);
  and (_09822_, _09803_, _08428_);
  or (_09824_, _09822_, _09820_);
  or (_09825_, _09824_, _09801_);
  not (_09826_, _09801_);
  or (_09827_, _09826_, word_in[9]);
  and (_09828_, _09827_, _09825_);
  or (_09829_, _09828_, _09808_);
  nor (_09830_, _09812_, _08422_);
  nor (_09831_, _09830_, _09800_);
  and (_09832_, _09831_, _09829_);
  and (_09833_, _09800_, _08973_);
  or (_26845_[1], _09833_, _09832_);
  not (_09834_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_09835_, _09803_, _09834_);
  and (_09836_, _09803_, _08591_);
  nor (_09838_, _09836_, _09835_);
  nor (_09840_, _09838_, _09801_);
  and (_09841_, _09801_, word_in[10]);
  or (_09842_, _09841_, _09808_);
  or (_09844_, _09842_, _09840_);
  or (_09845_, _09812_, _08715_);
  and (_09846_, _09845_, _09844_);
  and (_09847_, _09846_, _09816_);
  and (_09848_, _09800_, word_in[26]);
  or (_26845_[2], _09848_, _09847_);
  not (_09849_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_09850_, _09803_, _09849_);
  and (_09851_, _09803_, _08604_);
  nor (_09852_, _09851_, _09850_);
  nor (_09853_, _09852_, _09801_);
  and (_09855_, _09801_, word_in[11]);
  or (_09856_, _09855_, _09808_);
  or (_09857_, _09856_, _09853_);
  or (_09858_, _09812_, _08728_);
  and (_09859_, _09858_, _09857_);
  and (_09861_, _09859_, _09816_);
  and (_09862_, _09800_, word_in[27]);
  or (_26845_[3], _09862_, _09861_);
  not (_09863_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_09864_, _09803_, _09863_);
  and (_09865_, _09803_, _08619_);
  nor (_09866_, _09865_, _09864_);
  nor (_09867_, _09866_, _09801_);
  and (_09868_, _09801_, word_in[12]);
  or (_09869_, _09868_, _09808_);
  or (_09870_, _09869_, _09867_);
  or (_09871_, _09812_, _08744_);
  and (_09872_, _09871_, _09870_);
  or (_09873_, _09872_, _09800_);
  or (_09874_, _09816_, word_in[28]);
  and (_26845_[4], _09874_, _09873_);
  not (_09875_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_09876_, _09803_, _09875_);
  and (_09877_, _09803_, _08501_);
  or (_09878_, _09877_, _09876_);
  or (_09879_, _09878_, _09801_);
  or (_09880_, _09826_, word_in[13]);
  and (_09881_, _09880_, _09879_);
  or (_09882_, _09881_, _09808_);
  nor (_09883_, _09812_, _08758_);
  nor (_09884_, _09883_, _09800_);
  and (_09885_, _09884_, _09882_);
  and (_09886_, _09800_, _08495_);
  or (_26845_[5], _09886_, _09885_);
  not (_09888_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_09889_, _09803_, _09888_);
  and (_09890_, _09803_, _08648_);
  nor (_09891_, _09890_, _09889_);
  nor (_09892_, _09891_, _09801_);
  and (_09893_, _09801_, word_in[14]);
  or (_09894_, _09893_, _09808_);
  or (_09895_, _09894_, _09892_);
  or (_09896_, _09812_, _08774_);
  and (_09897_, _09896_, _09895_);
  and (_09898_, _09897_, _09816_);
  and (_09899_, _09800_, word_in[30]);
  or (_26845_[6], _09899_, _09898_);
  nor (_09901_, _09803_, _07731_);
  and (_09902_, _09803_, _08019_);
  or (_09903_, _09902_, _09901_);
  or (_09904_, _09903_, _09801_);
  nand (_09905_, _09801_, _09188_);
  and (_09907_, _09905_, _09904_);
  or (_09908_, _09907_, _09808_);
  nor (_09909_, _09812_, _08033_);
  nor (_09910_, _09909_, _09800_);
  and (_09911_, _09910_, _09908_);
  and (_09912_, _09800_, _09072_);
  or (_26845_[7], _09912_, _09911_);
  and (_09913_, _24275_, _23754_);
  and (_09914_, _09913_, _23747_);
  not (_09915_, _09913_);
  and (_09916_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_02539_, _09916_, _09914_);
  and (_09917_, _26112_, _26110_);
  nor (_09918_, _09917_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_09920_, _09917_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_09921_, _09920_, _09918_);
  and (_09922_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_09924_, _09922_, _26118_);
  nor (_09925_, _09924_, _09921_);
  nor (_09926_, _09925_, _24299_);
  and (_09927_, _24299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_09928_, _09927_, _09926_);
  and (_09929_, _09928_, _24294_);
  and (_09930_, _24293_, _23816_);
  or (_09931_, _09930_, _09929_);
  and (_02555_, _09931_, _22762_);
  and (_09932_, _24371_, _23747_);
  and (_09933_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_02571_, _09933_, _09932_);
  not (_09934_, _07948_);
  and (_09935_, _08929_, _09934_);
  and (_09936_, _09935_, _07790_);
  not (_09937_, _09936_);
  and (_09938_, _08008_, _07751_);
  not (_09939_, _09938_);
  and (_09941_, _08010_, _08244_);
  not (_09942_, _09941_);
  and (_09943_, _08396_, _08016_);
  and (_09944_, _09943_, word_in[0]);
  not (_09946_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_09947_, _09943_, _09946_);
  or (_09948_, _09947_, _09944_);
  and (_09949_, _09948_, _09942_);
  and (_09951_, _09941_, word_in[8]);
  or (_09953_, _09951_, _09949_);
  and (_09955_, _09953_, _09939_);
  and (_09957_, _09938_, _08678_);
  or (_09959_, _09957_, _09955_);
  and (_09960_, _09959_, _09937_);
  and (_09961_, _09936_, _08954_);
  or (_26846_[0], _09961_, _09960_);
  or (_09962_, _09939_, _08422_);
  not (_09963_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_09965_, _09943_, _09963_);
  and (_09967_, _09943_, _08428_);
  or (_09968_, _09967_, _09965_);
  or (_09969_, _09968_, _09941_);
  or (_09970_, _09942_, word_in[9]);
  and (_09971_, _09970_, _09969_);
  or (_09972_, _09971_, _09938_);
  and (_09973_, _09972_, _09962_);
  or (_09975_, _09973_, _09936_);
  or (_09977_, _09937_, _08973_);
  and (_26846_[1], _09977_, _09975_);
  or (_09978_, _09939_, _08715_);
  not (_09979_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_09980_, _09943_, _09979_);
  and (_09982_, _09943_, _08591_);
  or (_09983_, _09982_, _09980_);
  or (_09984_, _09983_, _09941_);
  or (_09985_, _09942_, word_in[10]);
  and (_09986_, _09985_, _09984_);
  or (_09987_, _09986_, _09938_);
  and (_09989_, _09987_, _09978_);
  or (_09990_, _09989_, _09936_);
  or (_09992_, _09937_, _08993_);
  and (_26846_[2], _09992_, _09990_);
  or (_09993_, _09939_, _08728_);
  not (_09994_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_09995_, _09943_, _09994_);
  and (_09996_, _09943_, _08604_);
  or (_09997_, _09996_, _09995_);
  or (_09998_, _09997_, _09941_);
  or (_09999_, _09942_, word_in[11]);
  and (_10000_, _09999_, _09998_);
  or (_10001_, _10000_, _09938_);
  and (_10002_, _10001_, _09993_);
  or (_10003_, _10002_, _09936_);
  or (_10004_, _09937_, _08461_);
  and (_26846_[3], _10004_, _10003_);
  or (_10006_, _09939_, _08744_);
  not (_10008_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_10009_, _09943_, _10008_);
  and (_10010_, _09943_, _08619_);
  or (_10011_, _10010_, _10009_);
  or (_10012_, _10011_, _09941_);
  or (_10014_, _09942_, word_in[12]);
  and (_10016_, _10014_, _10012_);
  or (_10017_, _10016_, _09938_);
  and (_10018_, _10017_, _10006_);
  or (_10019_, _10018_, _09936_);
  or (_10020_, _09937_, _08481_);
  and (_26846_[4], _10020_, _10019_);
  or (_10022_, _09939_, _08758_);
  not (_10023_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_10024_, _09943_, _10023_);
  and (_10025_, _09943_, _08501_);
  or (_10026_, _10025_, _10024_);
  or (_10027_, _10026_, _09941_);
  or (_10028_, _09942_, word_in[13]);
  and (_10029_, _10028_, _10027_);
  or (_10030_, _10029_, _09938_);
  and (_10031_, _10030_, _10022_);
  or (_10032_, _10031_, _09936_);
  or (_10033_, _09937_, _08495_);
  and (_26846_[5], _10033_, _10032_);
  or (_10034_, _09939_, _08774_);
  not (_10035_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_10037_, _09943_, _10035_);
  and (_10038_, _09943_, _08648_);
  or (_10040_, _10038_, _10037_);
  or (_10041_, _10040_, _09941_);
  or (_10042_, _09942_, word_in[14]);
  and (_10043_, _10042_, _10041_);
  or (_10044_, _10043_, _09938_);
  and (_10045_, _10044_, _10034_);
  or (_10046_, _10045_, _09936_);
  or (_10047_, _09937_, _08510_);
  and (_26846_[6], _10047_, _10046_);
  or (_10049_, _09939_, _08033_);
  nor (_10051_, _09943_, _07866_);
  and (_10052_, _09943_, _08019_);
  or (_10053_, _10052_, _10051_);
  or (_10054_, _10053_, _09941_);
  nand (_10056_, _09941_, _09188_);
  and (_10057_, _10056_, _10054_);
  or (_10058_, _10057_, _09938_);
  and (_10059_, _10058_, _10049_);
  or (_10060_, _10059_, _09936_);
  or (_10061_, _09937_, _09072_);
  and (_26846_[7], _10061_, _10060_);
  and (_10062_, _05042_, _23824_);
  and (_10063_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_27135_, _10063_, _10062_);
  and (_10064_, _08008_, _07754_);
  not (_10065_, _10064_);
  and (_10066_, _08553_, _07860_);
  and (_10067_, _08557_, _08016_);
  and (_10068_, _10067_, word_in[0]);
  not (_10069_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_10070_, _10067_, _10069_);
  nor (_10071_, _10070_, _10068_);
  nor (_10072_, _10071_, _10066_);
  and (_10073_, _10066_, word_in[8]);
  or (_10075_, _10073_, _10072_);
  and (_10076_, _10075_, _10065_);
  and (_10077_, _09935_, _07751_);
  and (_10078_, _10064_, _08678_);
  or (_10079_, _10078_, _10077_);
  or (_10080_, _10079_, _10076_);
  not (_10081_, _10077_);
  or (_10082_, _10081_, word_in[24]);
  and (_26847_[0], _10082_, _10080_);
  not (_10084_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_10086_, _10067_, _10084_);
  and (_10087_, _10067_, word_in[1]);
  or (_10088_, _10087_, _10086_);
  or (_10090_, _10088_, _10066_);
  not (_10091_, _10066_);
  or (_10092_, _10091_, word_in[9]);
  and (_10093_, _10092_, _10090_);
  or (_10094_, _10093_, _10064_);
  or (_10095_, _10065_, _08422_);
  and (_10096_, _10095_, _10094_);
  and (_10098_, _10096_, _10081_);
  and (_10099_, _10077_, word_in[25]);
  or (_26847_[1], _10099_, _10098_);
  or (_10101_, _10065_, _08715_);
  not (_10102_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_10103_, _10067_, _10102_);
  and (_10105_, _10067_, word_in[2]);
  or (_10106_, _10105_, _10103_);
  or (_10107_, _10106_, _10066_);
  or (_10109_, _10091_, word_in[10]);
  and (_10111_, _10109_, _10107_);
  or (_10112_, _10111_, _10064_);
  and (_10113_, _10112_, _10101_);
  or (_10115_, _10113_, _10077_);
  or (_10116_, _10081_, word_in[26]);
  and (_26847_[2], _10116_, _10115_);
  or (_10117_, _10065_, _08728_);
  not (_10118_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_10119_, _10067_, _10118_);
  and (_10120_, _10067_, word_in[3]);
  or (_10121_, _10120_, _10119_);
  or (_10122_, _10121_, _10066_);
  or (_10123_, _10091_, word_in[11]);
  and (_10124_, _10123_, _10122_);
  or (_10126_, _10124_, _10064_);
  and (_10127_, _10126_, _10117_);
  and (_10129_, _10127_, _10081_);
  and (_10131_, _10077_, word_in[27]);
  or (_26847_[3], _10131_, _10129_);
  or (_10134_, _10065_, _08744_);
  not (_10135_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_10136_, _10067_, _10135_);
  and (_10137_, _10067_, word_in[4]);
  or (_10139_, _10137_, _10136_);
  or (_10140_, _10139_, _10066_);
  or (_10141_, _10091_, word_in[12]);
  and (_10142_, _10141_, _10140_);
  or (_10144_, _10142_, _10064_);
  and (_10145_, _10144_, _10134_);
  and (_10146_, _10145_, _10081_);
  and (_10148_, _10077_, word_in[28]);
  or (_26847_[4], _10148_, _10146_);
  and (_10149_, _10067_, word_in[5]);
  not (_10150_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_10151_, _10067_, _10150_);
  nor (_10152_, _10151_, _10149_);
  nor (_10153_, _10152_, _10066_);
  and (_10154_, _10066_, word_in[13]);
  or (_10155_, _10154_, _10153_);
  and (_10156_, _10155_, _10065_);
  and (_10158_, _10064_, _08758_);
  or (_10159_, _10158_, _10077_);
  or (_10160_, _10159_, _10156_);
  or (_10162_, _10081_, word_in[29]);
  and (_26847_[5], _10162_, _10160_);
  or (_10164_, _10091_, word_in[14]);
  not (_10166_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_10167_, _10067_, _10166_);
  and (_10168_, _10067_, word_in[6]);
  or (_10170_, _10168_, _10167_);
  or (_10171_, _10170_, _10066_);
  and (_10173_, _10171_, _10065_);
  and (_10174_, _10173_, _10164_);
  and (_10175_, _10064_, _08774_);
  or (_10176_, _10175_, _10077_);
  or (_10177_, _10176_, _10174_);
  or (_10178_, _10081_, word_in[30]);
  and (_26847_[6], _10178_, _10177_);
  or (_10180_, _10065_, _08033_);
  nor (_10181_, _10067_, _07717_);
  and (_10183_, _10067_, word_in[7]);
  or (_10184_, _10183_, _10181_);
  or (_10185_, _10184_, _10066_);
  nand (_10187_, _10066_, _09188_);
  and (_10189_, _10187_, _10185_);
  or (_10190_, _10189_, _10064_);
  and (_10191_, _10190_, _10180_);
  and (_10193_, _10191_, _10081_);
  and (_10195_, _10077_, word_in[31]);
  or (_26847_[7], _10195_, _10193_);
  and (_10198_, _02359_, _23778_);
  and (_10199_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  or (_27154_, _10199_, _10198_);
  and (_10200_, _09935_, _07754_);
  and (_10202_, _08008_, _07780_);
  not (_10203_, _10202_);
  or (_10204_, _10203_, _08678_);
  and (_10205_, _08683_, _07860_);
  not (_10207_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_10208_, _08688_, _08016_);
  nor (_10209_, _10208_, _10207_);
  and (_10210_, _10208_, _08402_);
  or (_10211_, _10210_, _10209_);
  or (_10213_, _10211_, _10205_);
  not (_10214_, _10205_);
  or (_10215_, _10214_, word_in[8]);
  and (_10216_, _10215_, _10213_);
  or (_10217_, _10216_, _10202_);
  and (_10218_, _10217_, _10204_);
  or (_10219_, _10218_, _10200_);
  not (_10220_, _10200_);
  or (_10222_, _10220_, word_in[24]);
  and (_26848_[0], _10222_, _10219_);
  not (_10223_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_10224_, _10208_, _10223_);
  and (_10226_, _10208_, _08428_);
  or (_10228_, _10226_, _10224_);
  or (_10229_, _10228_, _10205_);
  or (_10230_, _10214_, word_in[9]);
  and (_10232_, _10230_, _10229_);
  or (_10233_, _10232_, _10202_);
  or (_10234_, _10203_, _08422_);
  and (_10235_, _10234_, _10233_);
  or (_10237_, _10235_, _10200_);
  or (_10238_, _10220_, word_in[25]);
  and (_26848_[1], _10238_, _10237_);
  not (_10241_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_10242_, _10208_, _10241_);
  and (_10243_, _10208_, _08591_);
  or (_10244_, _10243_, _10242_);
  or (_10245_, _10244_, _10205_);
  or (_10246_, _10214_, word_in[10]);
  and (_10247_, _10246_, _10245_);
  or (_10248_, _10247_, _10202_);
  nor (_10249_, _10203_, _08715_);
  nor (_10250_, _10249_, _10200_);
  and (_10251_, _10250_, _10248_);
  and (_10252_, _10200_, word_in[26]);
  or (_26848_[2], _10252_, _10251_);
  or (_10254_, _10203_, _08728_);
  not (_10255_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_10256_, _10208_, _10255_);
  and (_10257_, _10208_, _08604_);
  or (_10259_, _10257_, _10256_);
  or (_10261_, _10259_, _10205_);
  or (_10262_, _10214_, word_in[11]);
  and (_10263_, _10262_, _10261_);
  or (_10264_, _10263_, _10202_);
  and (_10265_, _10264_, _10254_);
  and (_10266_, _10265_, _10220_);
  and (_10267_, _10200_, word_in[27]);
  or (_26848_[3], _10267_, _10266_);
  or (_10268_, _10203_, _08744_);
  not (_10269_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_10270_, _10208_, _10269_);
  and (_10271_, _10208_, _08619_);
  or (_10272_, _10271_, _10270_);
  or (_10273_, _10272_, _10205_);
  or (_10274_, _10214_, word_in[12]);
  and (_10275_, _10274_, _10273_);
  or (_10276_, _10275_, _10202_);
  and (_10277_, _10276_, _10268_);
  or (_10278_, _10277_, _10200_);
  or (_10279_, _10220_, word_in[28]);
  and (_26848_[4], _10279_, _10278_);
  or (_10281_, _10203_, _08758_);
  not (_10282_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_10283_, _10208_, _10282_);
  and (_10284_, _10208_, _08501_);
  or (_10285_, _10284_, _10283_);
  or (_10286_, _10285_, _10205_);
  or (_10288_, _10214_, word_in[13]);
  and (_10290_, _10288_, _10286_);
  or (_10292_, _10290_, _10202_);
  and (_10294_, _10292_, _10281_);
  or (_10295_, _10294_, _10200_);
  or (_10296_, _10220_, word_in[29]);
  and (_26848_[5], _10296_, _10295_);
  not (_10298_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_10299_, _10208_, _10298_);
  and (_10300_, _10208_, _08648_);
  or (_10302_, _10300_, _10299_);
  or (_10303_, _10302_, _10205_);
  or (_10305_, _10214_, word_in[14]);
  and (_10306_, _10305_, _10303_);
  or (_10307_, _10306_, _10202_);
  nor (_10309_, _10203_, _08774_);
  nor (_10311_, _10309_, _10200_);
  and (_10312_, _10311_, _10307_);
  and (_10313_, _10200_, word_in[30]);
  or (_26848_[6], _10313_, _10312_);
  nor (_10315_, _10208_, _07861_);
  and (_10316_, _10208_, _08019_);
  or (_10318_, _10316_, _10315_);
  or (_10319_, _10318_, _10205_);
  nand (_10320_, _10205_, _09188_);
  and (_10321_, _10320_, _10319_);
  or (_10322_, _10321_, _10202_);
  nor (_10323_, _10203_, _08033_);
  nor (_10324_, _10323_, _10200_);
  and (_10325_, _10324_, _10322_);
  and (_10326_, _10200_, word_in[31]);
  or (_26848_[7], _10326_, _10325_);
  and (_10327_, _05180_, _23946_);
  and (_10328_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_27132_, _10328_, _10327_);
  and (_10331_, _06506_, _24282_);
  not (_10332_, _10331_);
  and (_10333_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  and (_10334_, _10331_, _23778_);
  or (_26981_, _10334_, _10333_);
  and (_10335_, _05180_, _23778_);
  and (_10337_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_27130_, _10337_, _10335_);
  and (_10339_, _08167_, _24050_);
  and (_10340_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or (_27129_, _10340_, _10339_);
  and (_10343_, _08167_, _23898_);
  and (_10344_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  or (_27128_, _10344_, _10343_);
  and (_10347_, _01809_, _23986_);
  and (_10348_, _10347_, _23946_);
  not (_10350_, _10347_);
  and (_10351_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  or (_27127_, _10351_, _10348_);
  and (_10352_, _10347_, _23747_);
  and (_10354_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or (_27126_, _10354_, _10352_);
  and (_10356_, _04797_, _24050_);
  and (_10357_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_27124_, _10357_, _10356_);
  and (_10358_, _04797_, _23649_);
  and (_10359_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_27123_, _10359_, _10358_);
  and (_10361_, _01810_, _24050_);
  and (_10362_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_27122_, _10362_, _10361_);
  and (_10363_, _01810_, _23649_);
  and (_10365_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_27121_, _10365_, _10363_);
  and (_10366_, _08954_, _08029_);
  and (_10367_, _08017_, word_in[0]);
  not (_10369_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_10371_, _08017_, _10369_);
  nor (_10372_, _10371_, _10367_);
  nor (_10373_, _10372_, _08012_);
  and (_10374_, _08012_, word_in[8]);
  or (_10376_, _10374_, _10373_);
  and (_10378_, _10376_, _08031_);
  and (_10380_, _08678_, _08009_);
  or (_10381_, _10380_, _10378_);
  and (_10383_, _10381_, _08030_);
  or (_26849_[0], _10383_, _10366_);
  and (_10385_, _01810_, _23778_);
  and (_10386_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_27120_, _10386_, _10385_);
  and (_10387_, _08017_, word_in[1]);
  not (_10388_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_10389_, _08017_, _10388_);
  nor (_10391_, _10389_, _10387_);
  nor (_10392_, _10391_, _08012_);
  and (_10393_, _08012_, word_in[9]);
  or (_10394_, _10393_, _10392_);
  and (_10396_, _10394_, _08031_);
  and (_10398_, _08422_, _08009_);
  or (_10400_, _10398_, _10396_);
  and (_10402_, _10400_, _08030_);
  and (_10404_, _08029_, word_in[25]);
  or (_26849_[1], _10404_, _10402_);
  and (_10405_, _02284_, _23707_);
  and (_10407_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or (_27119_, _10407_, _10405_);
  and (_10408_, _08017_, word_in[2]);
  not (_10410_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_10411_, _08017_, _10410_);
  nor (_10412_, _10411_, _10408_);
  nor (_10414_, _10412_, _08012_);
  and (_10415_, _08012_, word_in[10]);
  or (_10417_, _10415_, _10414_);
  and (_10418_, _10417_, _08031_);
  and (_10419_, _08715_, _08009_);
  or (_10420_, _10419_, _10418_);
  and (_10421_, _10420_, _08030_);
  and (_10422_, _08993_, _08029_);
  or (_26849_[2], _10422_, _10421_);
  and (_10423_, _02284_, _23946_);
  and (_10424_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or (_27118_, _10424_, _10423_);
  and (_10425_, _08017_, word_in[3]);
  not (_10426_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_10427_, _08017_, _10426_);
  nor (_10428_, _10427_, _10425_);
  nor (_10429_, _10428_, _08012_);
  and (_10430_, _08012_, word_in[11]);
  or (_10432_, _10430_, _10429_);
  and (_10433_, _10432_, _08031_);
  and (_10434_, _08728_, _08009_);
  or (_10435_, _10434_, _10433_);
  and (_10437_, _10435_, _08030_);
  and (_10438_, _08029_, word_in[27]);
  or (_26849_[3], _10438_, _10437_);
  and (_10439_, _08481_, _08029_);
  and (_10440_, _08017_, word_in[4]);
  not (_10441_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_10442_, _08017_, _10441_);
  nor (_10443_, _10442_, _10440_);
  nor (_10444_, _10443_, _08012_);
  and (_10445_, _08012_, word_in[12]);
  or (_10446_, _10445_, _10444_);
  and (_10447_, _10446_, _08031_);
  and (_10448_, _08744_, _08009_);
  or (_10449_, _10448_, _10447_);
  and (_10450_, _10449_, _08030_);
  or (_26849_[4], _10450_, _10439_);
  and (_10451_, _08017_, word_in[5]);
  not (_10453_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_10455_, _08017_, _10453_);
  nor (_10456_, _10455_, _10451_);
  nor (_10457_, _10456_, _08012_);
  and (_10458_, _08012_, word_in[13]);
  or (_10459_, _10458_, _10457_);
  and (_10460_, _10459_, _08031_);
  and (_10461_, _08758_, _08009_);
  or (_10462_, _10461_, _10460_);
  and (_10463_, _10462_, _08030_);
  and (_10464_, _08029_, word_in[29]);
  or (_26849_[5], _10464_, _10463_);
  and (_10465_, _08510_, _08029_);
  and (_10466_, _08017_, word_in[6]);
  not (_10467_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_10468_, _08017_, _10467_);
  nor (_10469_, _10468_, _10466_);
  nor (_10470_, _10469_, _08012_);
  and (_10472_, _08012_, word_in[14]);
  or (_10473_, _10472_, _10470_);
  and (_10474_, _10473_, _08031_);
  and (_10475_, _08774_, _08009_);
  or (_10476_, _10475_, _10474_);
  and (_10477_, _10476_, _08030_);
  or (_26849_[6], _10477_, _10465_);
  and (_10478_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and (_10479_, _08351_, _23946_);
  or (_02826_, _10479_, _10478_);
  and (_10480_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and (_10481_, _08375_, _23946_);
  or (_02844_, _10481_, _10480_);
  and (_10482_, _02302_, _23649_);
  and (_10483_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_02874_, _10483_, _10482_);
  and (_10484_, _02302_, _23778_);
  and (_10485_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_02876_, _10485_, _10484_);
  and (_10486_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  and (_10487_, _08375_, _24050_);
  or (_02880_, _10487_, _10486_);
  and (_10488_, _02374_, _23946_);
  and (_10489_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or (_02882_, _10489_, _10488_);
  and (_10490_, _03339_, _23747_);
  and (_10491_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_27113_, _10491_, _10490_);
  and (_10492_, _03339_, _23898_);
  and (_10493_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_27111_, _10493_, _10492_);
  and (_10494_, _24766_, _24282_);
  not (_10495_, _10494_);
  and (_10496_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and (_10497_, _10494_, _23778_);
  or (_02893_, _10497_, _10496_);
  and (_10498_, _04917_, _23649_);
  and (_10499_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_27109_, _10499_, _10498_);
  and (_10501_, _04917_, _23824_);
  and (_10502_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_02906_, _10502_, _10501_);
  and (_10503_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  and (_10504_, _10494_, _23898_);
  or (_02908_, _10504_, _10503_);
  and (_10505_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  and (_10506_, _10494_, _23747_);
  or (_02911_, _10506_, _10505_);
  and (_10507_, _07471_, _24050_);
  and (_10508_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or (_02923_, _10508_, _10507_);
  and (_10509_, _07673_, word_in[0]);
  nand (_10510_, _07570_, _08556_);
  or (_10512_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_10513_, _10512_, _10510_);
  and (_10514_, _10513_, _07624_);
  or (_10515_, _10514_, _07577_);
  nand (_10517_, _07570_, _09080_);
  or (_10518_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_10519_, _10518_, _10517_);
  and (_10520_, _10519_, _07591_);
  nand (_10521_, _07570_, _09333_);
  or (_10522_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_10523_, _10522_, _10521_);
  and (_10524_, _10523_, _07608_);
  nand (_10525_, _07570_, _08809_);
  or (_10526_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_10527_, _10526_, _10525_);
  and (_10528_, _10527_, _07597_);
  or (_10529_, _10528_, _10524_);
  or (_10530_, _10529_, _10520_);
  or (_10531_, _10530_, _10515_);
  nand (_10532_, _07570_, _09570_);
  or (_10533_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_10534_, _10533_, _10532_);
  and (_10535_, _10534_, _07624_);
  or (_10536_, _10535_, _07648_);
  nand (_10537_, _07570_, _10069_);
  or (_10538_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_10539_, _10538_, _10537_);
  and (_10541_, _10539_, _07591_);
  nand (_10542_, _07570_, _10369_);
  or (_10543_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_10544_, _10543_, _10542_);
  and (_10545_, _10544_, _07608_);
  nand (_10546_, _07570_, _09802_);
  or (_10547_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_10548_, _10547_, _10546_);
  and (_10549_, _10548_, _07597_);
  or (_10551_, _10549_, _10545_);
  or (_10552_, _10551_, _10541_);
  or (_10553_, _10552_, _10536_);
  and (_10554_, _10553_, _10531_);
  and (_10555_, _10554_, _07672_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _10555_, _10509_);
  and (_10556_, _07673_, word_in[1]);
  nand (_10557_, _07570_, _08575_);
  or (_10558_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_10560_, _10558_, _10557_);
  and (_10561_, _10560_, _07624_);
  or (_10562_, _10561_, _07577_);
  nand (_10563_, _07570_, _09098_);
  or (_10564_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_10565_, _10564_, _10563_);
  and (_10566_, _10565_, _07591_);
  nand (_10567_, _07570_, _09352_);
  or (_10568_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_10570_, _10568_, _10567_);
  and (_10571_, _10570_, _07608_);
  nand (_10572_, _07570_, _08830_);
  or (_10573_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_10575_, _10573_, _10572_);
  and (_10576_, _10575_, _07597_);
  or (_10577_, _10576_, _10571_);
  or (_10578_, _10577_, _10566_);
  or (_10579_, _10578_, _10562_);
  nand (_10580_, _07570_, _09586_);
  or (_10581_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_10582_, _10581_, _10580_);
  and (_10583_, _10582_, _07624_);
  or (_10584_, _10583_, _07648_);
  nand (_10585_, _07570_, _10084_);
  or (_10586_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_10587_, _10586_, _10585_);
  and (_10588_, _10587_, _07591_);
  nand (_10589_, _07570_, _10388_);
  or (_10590_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_10591_, _10590_, _10589_);
  and (_10592_, _10591_, _07608_);
  nand (_10593_, _07570_, _09819_);
  or (_10594_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_10595_, _10594_, _10593_);
  and (_10596_, _10595_, _07597_);
  or (_10597_, _10596_, _10592_);
  or (_10598_, _10597_, _10588_);
  or (_10600_, _10598_, _10584_);
  and (_10601_, _10600_, _10579_);
  and (_10602_, _10601_, _07672_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _10602_, _10556_);
  and (_10603_, _07673_, word_in[2]);
  nand (_10605_, _07570_, _08844_);
  or (_10607_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_10608_, _10607_, _10605_);
  and (_10609_, _10608_, _07597_);
  or (_10610_, _10609_, _07577_);
  nand (_10611_, _07570_, _09113_);
  or (_10612_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_10613_, _10612_, _10611_);
  and (_10614_, _10613_, _07591_);
  nand (_10615_, _07570_, _09371_);
  or (_10616_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_10617_, _10616_, _10615_);
  and (_10618_, _10617_, _07608_);
  nand (_10619_, _07570_, _08589_);
  or (_10620_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_10621_, _10620_, _10619_);
  and (_10622_, _10621_, _07624_);
  or (_10624_, _10622_, _10618_);
  or (_10626_, _10624_, _10614_);
  or (_10627_, _10626_, _10610_);
  nand (_10629_, _07570_, _09834_);
  or (_10630_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_10631_, _10630_, _10629_);
  and (_10632_, _10631_, _07597_);
  or (_10633_, _10632_, _07648_);
  nand (_10634_, _07570_, _10410_);
  or (_10635_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_10636_, _10635_, _10634_);
  and (_10637_, _10636_, _07608_);
  nand (_10638_, _07570_, _10102_);
  or (_10639_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_10640_, _10639_, _10638_);
  and (_10642_, _10640_, _07591_);
  or (_10643_, _10642_, _10637_);
  nand (_10644_, _07570_, _09598_);
  or (_10645_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_10647_, _10645_, _10644_);
  and (_10648_, _10647_, _07624_);
  or (_10649_, _10648_, _10643_);
  or (_10651_, _10649_, _10633_);
  and (_10653_, _10651_, _10627_);
  and (_10654_, _10653_, _07672_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _10654_, _10603_);
  and (_10655_, _07673_, word_in[3]);
  nand (_10656_, _07570_, _08857_);
  or (_10658_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_10659_, _10658_, _10656_);
  and (_10661_, _10659_, _07597_);
  or (_10662_, _10661_, _07577_);
  nand (_10663_, _07570_, _09128_);
  or (_10664_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_10665_, _10664_, _10663_);
  and (_10666_, _10665_, _07591_);
  nand (_10667_, _07570_, _09389_);
  or (_10668_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_10669_, _10668_, _10667_);
  and (_10670_, _10669_, _07608_);
  nand (_10671_, _07570_, _08602_);
  or (_10672_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_10673_, _10672_, _10671_);
  and (_10674_, _10673_, _07624_);
  or (_10675_, _10674_, _10670_);
  or (_10676_, _10675_, _10666_);
  or (_10678_, _10676_, _10662_);
  nand (_10680_, _07570_, _09849_);
  or (_10681_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_10682_, _10681_, _10680_);
  and (_10683_, _10682_, _07597_);
  or (_10684_, _10683_, _07648_);
  nand (_10685_, _07570_, _10426_);
  or (_10686_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_10687_, _10686_, _10685_);
  and (_10688_, _10687_, _07608_);
  nand (_10689_, _07570_, _10118_);
  or (_10690_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_10691_, _10690_, _10689_);
  and (_10692_, _10691_, _07591_);
  or (_10693_, _10692_, _10688_);
  nand (_10694_, _07570_, _09613_);
  or (_10695_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_10696_, _10695_, _10694_);
  and (_10697_, _10696_, _07624_);
  or (_10698_, _10697_, _10693_);
  or (_10699_, _10698_, _10684_);
  and (_10700_, _10699_, _10678_);
  and (_10702_, _10700_, _07672_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _10702_, _10655_);
  and (_10703_, _07673_, word_in[4]);
  nand (_10704_, _07570_, _08617_);
  or (_10705_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_10707_, _10705_, _10704_);
  and (_10708_, _10707_, _07624_);
  or (_10709_, _10708_, _07577_);
  nand (_10711_, _07570_, _09141_);
  or (_10712_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_10713_, _10712_, _10711_);
  and (_10714_, _10713_, _07591_);
  nand (_10715_, _07570_, _09402_);
  or (_10716_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_10717_, _10716_, _10715_);
  and (_10719_, _10717_, _07608_);
  nand (_10720_, _07570_, _08870_);
  or (_10721_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_10722_, _10721_, _10720_);
  and (_10723_, _10722_, _07597_);
  or (_10724_, _10723_, _10719_);
  or (_10725_, _10724_, _10714_);
  or (_10726_, _10725_, _10709_);
  nand (_10727_, _07570_, _09627_);
  or (_10728_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_10729_, _10728_, _10727_);
  and (_10730_, _10729_, _07624_);
  or (_10732_, _10730_, _07648_);
  nand (_10733_, _07570_, _10135_);
  or (_10734_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_10736_, _10734_, _10733_);
  and (_10738_, _10736_, _07591_);
  nand (_10739_, _07570_, _10441_);
  or (_10740_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_10741_, _10740_, _10739_);
  and (_10743_, _10741_, _07608_);
  nand (_10744_, _07570_, _09863_);
  or (_10746_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_10747_, _10746_, _10744_);
  and (_10749_, _10747_, _07597_);
  or (_10751_, _10749_, _10743_);
  or (_10752_, _10751_, _10738_);
  or (_10753_, _10752_, _10732_);
  and (_10754_, _10753_, _10726_);
  and (_10756_, _10754_, _07672_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _10756_, _10703_);
  and (_10758_, _07673_, word_in[5]);
  nand (_10759_, _07570_, _08630_);
  or (_10760_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_10761_, _10760_, _10759_);
  and (_10762_, _10761_, _07624_);
  or (_10763_, _10762_, _07577_);
  nand (_10764_, _07570_, _09153_);
  or (_10765_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_10766_, _10765_, _10764_);
  and (_10767_, _10766_, _07591_);
  nand (_10768_, _07570_, _09415_);
  or (_10769_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_10771_, _10769_, _10768_);
  and (_10772_, _10771_, _07608_);
  nand (_10773_, _07570_, _08883_);
  or (_10774_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_10776_, _10774_, _10773_);
  and (_10777_, _10776_, _07597_);
  or (_10778_, _10777_, _10772_);
  or (_10781_, _10778_, _10767_);
  or (_10782_, _10781_, _10763_);
  nand (_10783_, _07570_, _09641_);
  or (_10785_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_10786_, _10785_, _10783_);
  and (_10787_, _10786_, _07624_);
  or (_10789_, _10787_, _07648_);
  nand (_10790_, _07570_, _10150_);
  or (_10792_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_10793_, _10792_, _10790_);
  and (_10794_, _10793_, _07591_);
  nand (_10795_, _07570_, _10453_);
  or (_10796_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_10798_, _10796_, _10795_);
  and (_10800_, _10798_, _07608_);
  nand (_10801_, _07570_, _09875_);
  or (_10802_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_10803_, _10802_, _10801_);
  and (_10804_, _10803_, _07597_);
  or (_10805_, _10804_, _10800_);
  or (_10807_, _10805_, _10794_);
  or (_10808_, _10807_, _10789_);
  and (_10809_, _10808_, _10782_);
  and (_10811_, _10809_, _07672_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _10811_, _10758_);
  and (_10812_, _07673_, word_in[6]);
  nand (_10814_, _07570_, _08898_);
  or (_10815_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_10816_, _10815_, _10814_);
  and (_10817_, _10816_, _07597_);
  or (_10818_, _10817_, _07577_);
  nand (_10819_, _07570_, _09166_);
  or (_10820_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_10821_, _10820_, _10819_);
  and (_10822_, _10821_, _07591_);
  nand (_10823_, _07570_, _09428_);
  or (_10824_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_10825_, _10824_, _10823_);
  and (_10827_, _10825_, _07608_);
  nand (_10828_, _07570_, _08646_);
  or (_10831_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_10833_, _10831_, _10828_);
  and (_10835_, _10833_, _07624_);
  or (_10836_, _10835_, _10827_);
  or (_10837_, _10836_, _10822_);
  or (_10839_, _10837_, _10818_);
  nand (_10840_, _07570_, _09888_);
  or (_10841_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_10842_, _10841_, _10840_);
  and (_10843_, _10842_, _07597_);
  or (_10845_, _10843_, _07648_);
  nand (_10846_, _07570_, _10467_);
  or (_10847_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_10848_, _10847_, _10846_);
  and (_10849_, _10848_, _07608_);
  nand (_10850_, _07570_, _10166_);
  or (_10851_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_10852_, _10851_, _10850_);
  and (_10853_, _10852_, _07591_);
  or (_10854_, _10853_, _10849_);
  nand (_10857_, _07570_, _09654_);
  or (_10858_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_10859_, _10858_, _10857_);
  and (_10860_, _10859_, _07624_);
  or (_10861_, _10860_, _10854_);
  or (_10862_, _10861_, _10845_);
  and (_10863_, _10862_, _10839_);
  and (_10865_, _10863_, _07672_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _10865_, _10812_);
  and (_10866_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  and (_10867_, _10494_, _23649_);
  or (_27024_, _10867_, _10866_);
  and (_10868_, _07810_, word_in[8]);
  nand (_10869_, _07570_, _08686_);
  or (_10870_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_10871_, _10870_, _10869_);
  and (_10872_, _10871_, _07812_);
  nand (_10874_, _07570_, _08393_);
  or (_10875_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_10877_, _10875_, _10874_);
  and (_10878_, _10877_, _07811_);
  or (_10879_, _10878_, _10872_);
  and (_10881_, _10879_, _07766_);
  nand (_10882_, _07570_, _09686_);
  or (_10883_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_10884_, _10883_, _10882_);
  and (_10885_, _10884_, _07812_);
  nand (_10887_, _07570_, _09453_);
  or (_10889_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_10890_, _10889_, _10887_);
  and (_10893_, _10890_, _07811_);
  or (_10894_, _10893_, _10885_);
  and (_10896_, _10894_, _07770_);
  nand (_10898_, _07570_, _09200_);
  or (_10899_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_10900_, _10899_, _10898_);
  and (_10901_, _10900_, _07812_);
  nand (_10903_, _07570_, _08938_);
  or (_10904_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_10905_, _10904_, _10903_);
  and (_10906_, _10905_, _07811_);
  or (_10907_, _10906_, _10901_);
  and (_10908_, _10907_, _07845_);
  nand (_10909_, _07570_, _10207_);
  or (_10910_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_10911_, _10910_, _10909_);
  and (_10912_, _10911_, _07812_);
  nand (_10913_, _07570_, _09946_);
  or (_10914_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_10916_, _10914_, _10913_);
  and (_10917_, _10916_, _07811_);
  or (_10918_, _10917_, _10912_);
  and (_10919_, _10918_, _07860_);
  or (_10921_, _10919_, _10908_);
  or (_10922_, _10921_, _10896_);
  nor (_10923_, _10922_, _10881_);
  nor (_10924_, _10923_, _07810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _10924_, _10868_);
  and (_10925_, _07810_, word_in[9]);
  nand (_10926_, _07570_, _08702_);
  or (_10927_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_10929_, _10927_, _10926_);
  and (_10931_, _10929_, _07812_);
  nand (_10932_, _07570_, _08425_);
  or (_10933_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_10934_, _10933_, _10932_);
  and (_10935_, _10934_, _07811_);
  or (_10936_, _10935_, _10931_);
  and (_10937_, _10936_, _07766_);
  nand (_10939_, _07570_, _09703_);
  or (_10941_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_10942_, _10941_, _10939_);
  and (_10943_, _10942_, _07812_);
  nand (_10944_, _07570_, _09474_);
  or (_10946_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_10948_, _10946_, _10944_);
  and (_10949_, _10948_, _07811_);
  or (_10950_, _10949_, _10943_);
  and (_10951_, _10950_, _07770_);
  nand (_10953_, _07570_, _09222_);
  or (_10954_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_10956_, _10954_, _10953_);
  and (_10957_, _10956_, _07812_);
  nand (_10959_, _07570_, _08957_);
  or (_10961_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_10962_, _10961_, _10959_);
  and (_10963_, _10962_, _07811_);
  or (_10964_, _10963_, _10957_);
  and (_10965_, _10964_, _07845_);
  nand (_10967_, _07570_, _10223_);
  or (_10969_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_10970_, _10969_, _10967_);
  and (_10971_, _10970_, _07812_);
  nand (_10972_, _07570_, _09963_);
  or (_10974_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_10976_, _10974_, _10972_);
  and (_10977_, _10976_, _07811_);
  or (_10978_, _10977_, _10971_);
  and (_10979_, _10978_, _07860_);
  or (_10981_, _10979_, _10965_);
  or (_10983_, _10981_, _10951_);
  nor (_10984_, _10983_, _10937_);
  nor (_10985_, _10984_, _07810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _10985_, _10925_);
  and (_10986_, _07810_, word_in[10]);
  nand (_10987_, _07570_, _08717_);
  or (_10988_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_10989_, _10988_, _10987_);
  and (_10990_, _10989_, _07812_);
  nand (_10991_, _07570_, _08450_);
  or (_10992_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_10993_, _10992_, _10991_);
  and (_10994_, _10993_, _07811_);
  or (_10995_, _10994_, _10990_);
  and (_10996_, _10995_, _07766_);
  nand (_10997_, _07570_, _09716_);
  or (_10998_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_10999_, _10998_, _10997_);
  and (_11000_, _10999_, _07812_);
  nand (_11001_, _07570_, _09486_);
  or (_11002_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_11003_, _11002_, _11001_);
  and (_11004_, _11003_, _07811_);
  or (_11005_, _11004_, _11000_);
  and (_11006_, _11005_, _07770_);
  nand (_11007_, _07570_, _09236_);
  or (_11008_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_11009_, _11008_, _11007_);
  and (_11010_, _11009_, _07812_);
  nand (_11011_, _07570_, _08979_);
  or (_11012_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_11013_, _11012_, _11011_);
  and (_11014_, _11013_, _07811_);
  or (_11015_, _11014_, _11010_);
  and (_11016_, _11015_, _07845_);
  nand (_11017_, _07570_, _10241_);
  or (_11018_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_11019_, _11018_, _11017_);
  and (_11020_, _11019_, _07812_);
  nand (_11021_, _07570_, _09979_);
  or (_11022_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_11023_, _11022_, _11021_);
  and (_11024_, _11023_, _07811_);
  or (_11025_, _11024_, _11020_);
  and (_11026_, _11025_, _07860_);
  or (_11027_, _11026_, _11016_);
  or (_11028_, _11027_, _11006_);
  nor (_11029_, _11028_, _10996_);
  nor (_11030_, _11029_, _07810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _11030_, _10986_);
  and (_11031_, _07810_, word_in[11]);
  nand (_11032_, _07570_, _08730_);
  or (_11033_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_11034_, _11033_, _11032_);
  and (_11035_, _11034_, _07812_);
  nand (_11036_, _07570_, _08467_);
  or (_11037_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_11038_, _11037_, _11036_);
  and (_11039_, _11038_, _07811_);
  or (_11040_, _11039_, _11035_);
  and (_11041_, _11040_, _07766_);
  nand (_11042_, _07570_, _09732_);
  or (_11043_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_11044_, _11043_, _11042_);
  and (_11045_, _11044_, _07812_);
  nand (_11046_, _07570_, _09499_);
  or (_11047_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_11048_, _11047_, _11046_);
  and (_11049_, _11048_, _07811_);
  or (_11050_, _11049_, _11045_);
  and (_11052_, _11050_, _07770_);
  nand (_11054_, _07570_, _09248_);
  or (_11055_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_11056_, _11055_, _11054_);
  and (_11058_, _11056_, _07812_);
  nand (_11059_, _07570_, _08996_);
  or (_11060_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_11061_, _11060_, _11059_);
  and (_11063_, _11061_, _07811_);
  or (_11064_, _11063_, _11058_);
  and (_11065_, _11064_, _07845_);
  nand (_11066_, _07570_, _10255_);
  or (_11067_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_11068_, _11067_, _11066_);
  and (_11069_, _11068_, _07812_);
  nand (_11070_, _07570_, _09994_);
  or (_11072_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_11073_, _11072_, _11070_);
  and (_11075_, _11073_, _07811_);
  or (_11076_, _11075_, _11069_);
  and (_11078_, _11076_, _07860_);
  or (_11079_, _11078_, _11065_);
  or (_11081_, _11079_, _11052_);
  nor (_11082_, _11081_, _11041_);
  nor (_11084_, _11082_, _07810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _11084_, _11031_);
  and (_11087_, _07810_, word_in[12]);
  nand (_11088_, _07570_, _08746_);
  or (_11089_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_11090_, _11089_, _11088_);
  and (_11093_, _11090_, _07812_);
  nand (_11095_, _07570_, _08485_);
  or (_11096_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_11097_, _11096_, _11095_);
  and (_11098_, _11097_, _07811_);
  or (_11099_, _11098_, _11093_);
  and (_11101_, _11099_, _07766_);
  nand (_11103_, _07570_, _09746_);
  or (_11105_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_11107_, _11105_, _11103_);
  and (_11108_, _11107_, _07812_);
  nand (_11110_, _07570_, _09512_);
  or (_11112_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_11113_, _11112_, _11110_);
  and (_11114_, _11113_, _07811_);
  or (_11115_, _11114_, _11108_);
  and (_11116_, _11115_, _07770_);
  nand (_11118_, _07570_, _09262_);
  or (_11120_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_11121_, _11120_, _11118_);
  and (_11122_, _11121_, _07812_);
  nand (_11123_, _07570_, _09013_);
  or (_11125_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_11126_, _11125_, _11123_);
  and (_11128_, _11126_, _07811_);
  or (_11129_, _11128_, _11122_);
  and (_11130_, _11129_, _07845_);
  nand (_11131_, _07570_, _10269_);
  or (_11133_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_11135_, _11133_, _11131_);
  and (_11137_, _11135_, _07812_);
  nand (_11138_, _07570_, _10008_);
  or (_11140_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_11142_, _11140_, _11138_);
  and (_11143_, _11142_, _07811_);
  or (_11144_, _11143_, _11137_);
  and (_11145_, _11144_, _07860_);
  or (_11146_, _11145_, _11130_);
  or (_11148_, _11146_, _11116_);
  nor (_11150_, _11148_, _11101_);
  nor (_11151_, _11150_, _07810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _11151_, _11087_);
  and (_11152_, _07810_, word_in[13]);
  nand (_11154_, _07570_, _08760_);
  or (_11155_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_11157_, _11155_, _11154_);
  and (_11158_, _11157_, _07812_);
  nand (_11160_, _07570_, _08499_);
  or (_11162_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_11163_, _11162_, _11160_);
  and (_11165_, _11163_, _07811_);
  or (_11166_, _11165_, _11158_);
  and (_11167_, _11166_, _07766_);
  nand (_11168_, _07570_, _09760_);
  or (_11169_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_11170_, _11169_, _11168_);
  and (_11171_, _11170_, _07812_);
  nand (_11172_, _07570_, _09525_);
  or (_11173_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_11174_, _11173_, _11172_);
  and (_11176_, _11174_, _07811_);
  or (_11177_, _11176_, _11171_);
  and (_11178_, _11177_, _07770_);
  nand (_11179_, _07570_, _09279_);
  or (_11180_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_11181_, _11180_, _11179_);
  and (_11182_, _11181_, _07812_);
  nand (_11184_, _07570_, _09029_);
  or (_11185_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_11186_, _11185_, _11184_);
  and (_11187_, _11186_, _07811_);
  or (_11188_, _11187_, _11182_);
  and (_11190_, _11188_, _07845_);
  nand (_11191_, _07570_, _10282_);
  or (_11192_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_11194_, _11192_, _11191_);
  and (_11196_, _11194_, _07812_);
  nand (_11197_, _07570_, _10023_);
  or (_11198_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_11199_, _11198_, _11197_);
  and (_11201_, _11199_, _07811_);
  or (_11202_, _11201_, _11196_);
  and (_11204_, _11202_, _07860_);
  or (_11205_, _11204_, _11190_);
  or (_11206_, _11205_, _11178_);
  nor (_11208_, _11206_, _11167_);
  nor (_11209_, _11208_, _07810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _11209_, _11152_);
  and (_11210_, _07810_, word_in[14]);
  nand (_11211_, _07570_, _08776_);
  or (_11212_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_11213_, _11212_, _11211_);
  and (_11214_, _11213_, _07812_);
  nand (_11215_, _07570_, _08515_);
  or (_11217_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_11218_, _11217_, _11215_);
  and (_11219_, _11218_, _07811_);
  or (_11220_, _11219_, _11214_);
  and (_11221_, _11220_, _07766_);
  nand (_11223_, _07570_, _09774_);
  or (_11224_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_11225_, _11224_, _11223_);
  and (_11226_, _11225_, _07812_);
  nand (_11227_, _07570_, _09537_);
  or (_11229_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_11231_, _11229_, _11227_);
  and (_11232_, _11231_, _07811_);
  or (_11233_, _11232_, _11226_);
  and (_11234_, _11233_, _07770_);
  nand (_11235_, _07570_, _09293_);
  or (_11237_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_11238_, _11237_, _11235_);
  and (_11239_, _11238_, _07812_);
  nand (_11240_, _07570_, _09043_);
  or (_11241_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_11243_, _11241_, _11240_);
  and (_11245_, _11243_, _07811_);
  or (_11247_, _11245_, _11239_);
  and (_11248_, _11247_, _07845_);
  nand (_11249_, _07570_, _10298_);
  or (_11250_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_11251_, _11250_, _11249_);
  and (_11253_, _11251_, _07812_);
  nand (_11254_, _07570_, _10035_);
  or (_11256_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_11257_, _11256_, _11254_);
  and (_11259_, _11257_, _07811_);
  or (_11260_, _11259_, _11253_);
  and (_11261_, _11260_, _07860_);
  or (_11263_, _11261_, _11248_);
  or (_11264_, _11263_, _11234_);
  nor (_11266_, _11264_, _11221_);
  nor (_11268_, _11266_, _07810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _11268_, _11210_);
  and (_11269_, _07471_, _23898_);
  and (_11271_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or (_02972_, _11271_, _11269_);
  and (_11272_, _07914_, word_in[16]);
  and (_11274_, _10523_, _07591_);
  and (_11275_, _10527_, _07624_);
  or (_11276_, _11275_, _11274_);
  and (_11277_, _10519_, _07597_);
  and (_11278_, _10513_, _07608_);
  or (_11279_, _11278_, _11277_);
  or (_11281_, _11279_, _11276_);
  or (_11282_, _11281_, _07881_);
  and (_11283_, _10548_, _07624_);
  and (_11284_, _10534_, _07608_);
  or (_11285_, _11284_, _11283_);
  and (_11287_, _10544_, _07591_);
  and (_11288_, _10539_, _07597_);
  or (_11290_, _11288_, _11287_);
  or (_11291_, _11290_, _11285_);
  or (_11292_, _11291_, _07915_);
  nand (_11293_, _11292_, _11282_);
  nor (_11294_, _11293_, _07914_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _11294_, _11272_);
  and (_11295_, _07914_, word_in[17]);
  and (_11297_, _10575_, _07624_);
  and (_11298_, _10565_, _07597_);
  or (_11300_, _11298_, _11297_);
  and (_11301_, _10570_, _07591_);
  and (_11302_, _10560_, _07608_);
  or (_11303_, _11302_, _11301_);
  or (_11304_, _11303_, _11300_);
  or (_11305_, _11304_, _07881_);
  and (_11306_, _10591_, _07591_);
  and (_11308_, _10587_, _07597_);
  or (_11309_, _11308_, _11306_);
  and (_11310_, _10595_, _07624_);
  and (_11311_, _10582_, _07608_);
  or (_11313_, _11311_, _11310_);
  or (_11314_, _11313_, _11309_);
  or (_11316_, _11314_, _07915_);
  nand (_11318_, _11316_, _11305_);
  nor (_11320_, _11318_, _07914_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _11320_, _11295_);
  and (_11321_, _07914_, word_in[18]);
  and (_11323_, _10617_, _07591_);
  and (_11324_, _10608_, _07624_);
  or (_11325_, _11324_, _11323_);
  and (_11326_, _10613_, _07597_);
  and (_11327_, _10621_, _07608_);
  or (_11328_, _11327_, _11326_);
  or (_11330_, _11328_, _11325_);
  or (_11332_, _11330_, _07881_);
  and (_11333_, _10631_, _07624_);
  and (_11334_, _10640_, _07597_);
  or (_11336_, _11334_, _11333_);
  and (_11337_, _10636_, _07591_);
  and (_11338_, _10647_, _07608_);
  or (_11339_, _11338_, _11337_);
  or (_11340_, _11339_, _11336_);
  or (_11342_, _11340_, _07915_);
  nand (_11343_, _11342_, _11332_);
  nor (_11344_, _11343_, _07914_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _11344_, _11321_);
  and (_11345_, _07914_, word_in[19]);
  and (_11347_, _10659_, _07624_);
  and (_11348_, _10665_, _07597_);
  or (_11350_, _11348_, _11347_);
  and (_11351_, _10669_, _07591_);
  and (_11352_, _10673_, _07608_);
  or (_11354_, _11352_, _11351_);
  or (_11355_, _11354_, _11350_);
  or (_11357_, _11355_, _07881_);
  and (_11359_, _10682_, _07624_);
  and (_11360_, _10691_, _07597_);
  or (_11361_, _11360_, _11359_);
  and (_11362_, _10687_, _07591_);
  and (_11363_, _10696_, _07608_);
  or (_11365_, _11363_, _11362_);
  or (_11366_, _11365_, _11361_);
  or (_11367_, _11366_, _07915_);
  nand (_11369_, _11367_, _11357_);
  nor (_11370_, _11369_, _07914_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _11370_, _11345_);
  and (_11371_, _07914_, word_in[20]);
  and (_11372_, _10722_, _07624_);
  and (_11373_, _10713_, _07597_);
  or (_11375_, _11373_, _11372_);
  and (_11377_, _10717_, _07591_);
  and (_11378_, _10707_, _07608_);
  or (_11379_, _11378_, _11377_);
  or (_11380_, _11379_, _11375_);
  or (_11381_, _11380_, _07881_);
  and (_11382_, _10741_, _07591_);
  and (_11383_, _10747_, _07624_);
  or (_11384_, _11383_, _11382_);
  and (_11385_, _10736_, _07597_);
  and (_11386_, _10729_, _07608_);
  or (_11387_, _11386_, _11385_);
  or (_11389_, _11387_, _11384_);
  or (_11390_, _11389_, _07915_);
  nand (_11391_, _11390_, _11381_);
  nor (_11392_, _11391_, _07914_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _11392_, _11371_);
  and (_11393_, _07914_, word_in[21]);
  and (_11395_, _10766_, _07597_);
  and (_11397_, _10761_, _07608_);
  or (_11398_, _11397_, _11395_);
  and (_11399_, _10771_, _07591_);
  and (_11401_, _10776_, _07624_);
  or (_11402_, _11401_, _11399_);
  or (_11403_, _11402_, _11398_);
  or (_11405_, _11403_, _07881_);
  and (_11407_, _10793_, _07597_);
  and (_11409_, _10786_, _07608_);
  or (_11411_, _11409_, _11407_);
  and (_11412_, _10798_, _07591_);
  and (_11415_, _10803_, _07624_);
  or (_11416_, _11415_, _11412_);
  or (_11417_, _11416_, _11411_);
  or (_11419_, _11417_, _07915_);
  nand (_11420_, _11419_, _11405_);
  nor (_11421_, _11420_, _07914_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _11421_, _11393_);
  and (_11422_, _07914_, word_in[22]);
  and (_11423_, _10825_, _07591_);
  and (_11424_, _10816_, _07624_);
  or (_11426_, _11424_, _11423_);
  and (_11427_, _10821_, _07597_);
  and (_11428_, _10833_, _07608_);
  or (_11429_, _11428_, _11427_);
  or (_11430_, _11429_, _11426_);
  or (_11431_, _11430_, _07881_);
  and (_11432_, _10848_, _07591_);
  and (_11433_, _10842_, _07624_);
  or (_11434_, _11433_, _11432_);
  and (_11435_, _10852_, _07597_);
  and (_11436_, _10859_, _07608_);
  or (_11437_, _11436_, _11435_);
  or (_11438_, _11437_, _11434_);
  or (_11439_, _11438_, _07915_);
  nand (_11440_, _11439_, _11431_);
  nor (_11441_, _11440_, _07914_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _11441_, _11422_);
  and (_11442_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  and (_11443_, _10494_, _23707_);
  or (_02996_, _11443_, _11442_);
  and (_11444_, _07975_, word_in[24]);
  and (_11445_, _10877_, _07812_);
  and (_11446_, _10871_, _07811_);
  or (_11447_, _11446_, _11445_);
  and (_11448_, _11447_, _07949_);
  and (_11449_, _10890_, _07812_);
  and (_11450_, _10884_, _07811_);
  or (_11451_, _11450_, _11449_);
  and (_11452_, _11451_, _07951_);
  and (_11453_, _10905_, _07812_);
  and (_11455_, _10900_, _07811_);
  or (_11457_, _11455_, _11453_);
  and (_11459_, _11457_, _07984_);
  and (_11461_, _10916_, _07812_);
  and (_11462_, _10911_, _07811_);
  or (_11464_, _11462_, _11461_);
  and (_11465_, _11464_, _07992_);
  or (_11466_, _11465_, _11459_);
  or (_11467_, _11466_, _11452_);
  nor (_11469_, _11467_, _11448_);
  nor (_11470_, _11469_, _07975_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _11470_, _11444_);
  and (_11472_, _07975_, word_in[25]);
  and (_11474_, _10934_, _07812_);
  and (_11475_, _10929_, _07811_);
  or (_11476_, _11475_, _11474_);
  and (_11477_, _11476_, _07949_);
  and (_11479_, _10948_, _07812_);
  and (_11480_, _10942_, _07811_);
  or (_11481_, _11480_, _11479_);
  and (_11484_, _11481_, _07951_);
  and (_11486_, _10962_, _07812_);
  and (_11488_, _10956_, _07811_);
  or (_11490_, _11488_, _11486_);
  and (_11492_, _11490_, _07984_);
  and (_11494_, _10976_, _07812_);
  and (_11495_, _10970_, _07811_);
  or (_11496_, _11495_, _11494_);
  and (_11498_, _11496_, _07992_);
  or (_11500_, _11498_, _11492_);
  or (_11501_, _11500_, _11484_);
  nor (_11503_, _11501_, _11477_);
  nor (_11504_, _11503_, _07975_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _11504_, _11472_);
  and (_11507_, _07975_, word_in[26]);
  and (_11508_, _10993_, _07812_);
  and (_11509_, _10989_, _07811_);
  or (_11511_, _11509_, _11508_);
  and (_11513_, _11511_, _07949_);
  and (_11514_, _11003_, _07812_);
  and (_11516_, _10999_, _07811_);
  or (_11517_, _11516_, _11514_);
  and (_11518_, _11517_, _07951_);
  and (_11520_, _11013_, _07812_);
  and (_11521_, _11009_, _07811_);
  or (_11523_, _11521_, _11520_);
  and (_11525_, _11523_, _07984_);
  and (_11527_, _11023_, _07812_);
  and (_11529_, _11019_, _07811_);
  or (_11530_, _11529_, _11527_);
  and (_11531_, _11530_, _07992_);
  or (_11533_, _11531_, _11525_);
  or (_11535_, _11533_, _11518_);
  nor (_11536_, _11535_, _11513_);
  nor (_11537_, _11536_, _07975_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _11537_, _11507_);
  and (_11540_, _07975_, word_in[27]);
  and (_11542_, _11038_, _07812_);
  and (_11544_, _11034_, _07811_);
  or (_11546_, _11544_, _11542_);
  and (_11547_, _11546_, _07949_);
  and (_11549_, _11048_, _07812_);
  and (_11550_, _11044_, _07811_);
  or (_11551_, _11550_, _11549_);
  and (_11552_, _11551_, _07951_);
  and (_11553_, _11061_, _07812_);
  and (_11554_, _11056_, _07811_);
  or (_11555_, _11554_, _11553_);
  and (_11556_, _11555_, _07984_);
  and (_11557_, _11073_, _07812_);
  and (_11559_, _11068_, _07811_);
  or (_11560_, _11559_, _11557_);
  and (_11561_, _11560_, _07992_);
  or (_11563_, _11561_, _11556_);
  or (_11564_, _11563_, _11552_);
  nor (_11566_, _11564_, _11547_);
  nor (_11567_, _11566_, _07975_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _11567_, _11540_);
  and (_11570_, _07975_, word_in[28]);
  and (_11571_, _11097_, _07812_);
  and (_11572_, _11090_, _07811_);
  or (_11573_, _11572_, _11571_);
  and (_11574_, _11573_, _07949_);
  and (_11575_, _11113_, _07812_);
  and (_11576_, _11107_, _07811_);
  or (_11578_, _11576_, _11575_);
  and (_11579_, _11578_, _07951_);
  and (_11580_, _11126_, _07812_);
  and (_11581_, _11121_, _07811_);
  or (_11582_, _11581_, _11580_);
  and (_11584_, _11582_, _07984_);
  and (_11585_, _11142_, _07812_);
  and (_11586_, _11135_, _07811_);
  or (_11587_, _11586_, _11585_);
  and (_11588_, _11587_, _07992_);
  or (_11589_, _11588_, _11584_);
  or (_11590_, _11589_, _11579_);
  nor (_11592_, _11590_, _11574_);
  nor (_11593_, _11592_, _07975_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _11593_, _11570_);
  and (_11594_, _07975_, word_in[29]);
  and (_11596_, _11163_, _07812_);
  and (_11597_, _11157_, _07811_);
  or (_11598_, _11597_, _11596_);
  and (_11599_, _11598_, _07949_);
  and (_11600_, _11174_, _07812_);
  and (_11601_, _11170_, _07811_);
  or (_11602_, _11601_, _11600_);
  and (_11603_, _11602_, _07951_);
  and (_11605_, _11186_, _07812_);
  and (_11606_, _11181_, _07811_);
  or (_11607_, _11606_, _11605_);
  and (_11608_, _11607_, _07984_);
  and (_11610_, _11199_, _07812_);
  and (_11611_, _11194_, _07811_);
  or (_11612_, _11611_, _11610_);
  and (_11614_, _11612_, _07992_);
  or (_11616_, _11614_, _11608_);
  or (_11618_, _11616_, _11603_);
  nor (_11619_, _11618_, _11599_);
  nor (_11620_, _11619_, _07975_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _11620_, _11594_);
  and (_11623_, _07975_, word_in[30]);
  and (_11624_, _11231_, _07812_);
  and (_11626_, _11225_, _07811_);
  or (_11627_, _11626_, _11624_);
  and (_11629_, _11627_, _07951_);
  and (_11630_, _11218_, _07812_);
  and (_11631_, _11213_, _07811_);
  or (_11632_, _11631_, _11630_);
  and (_11633_, _11632_, _07949_);
  and (_11634_, _11243_, _07812_);
  and (_11635_, _11238_, _07811_);
  or (_11636_, _11635_, _11634_);
  and (_11638_, _11636_, _07984_);
  and (_11639_, _11257_, _07812_);
  and (_11640_, _11251_, _07811_);
  or (_11641_, _11640_, _11639_);
  and (_11642_, _11641_, _07992_);
  or (_11644_, _11642_, _11638_);
  or (_11646_, _11644_, _11633_);
  nor (_11647_, _11646_, _11629_);
  nor (_11648_, _11647_, _07975_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _11648_, _11623_);
  and (_11649_, _05445_, _23707_);
  and (_11650_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  or (_03046_, _11650_, _11649_);
  and (_11652_, _25078_, _24766_);
  not (_11653_, _11652_);
  and (_11654_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_11655_, _11652_, _23778_);
  or (_03052_, _11655_, _11654_);
  and (_11657_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_11658_, _11652_, _23824_);
  or (_03069_, _11658_, _11657_);
  and (_11660_, _05445_, _23824_);
  and (_11661_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  or (_03108_, _11661_, _11660_);
  and (_11664_, _02374_, _23778_);
  and (_11666_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  or (_03114_, _11666_, _11664_);
  and (_11667_, _24086_, _23898_);
  and (_11668_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_03117_, _11668_, _11667_);
  and (_11669_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_11670_, _11652_, _23747_);
  or (_03123_, _11670_, _11669_);
  and (_11671_, _07536_, _23946_);
  and (_11672_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or (_03125_, _11672_, _11671_);
  and (_11673_, _07536_, _23898_);
  and (_11674_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  or (_03129_, _11674_, _11673_);
  and (_11675_, _07536_, _23747_);
  and (_11676_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or (_03139_, _11676_, _11675_);
  and (_11678_, _02345_, _23824_);
  and (_11679_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_27191_, _11679_, _11678_);
  and (_11680_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_11682_, _11652_, _24050_);
  or (_03144_, _11682_, _11680_);
  nor (_26887_[1], _00094_, rst);
  and (_11685_, _05180_, _23824_);
  and (_11686_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_03160_, _11686_, _11685_);
  and (_11688_, _08167_, _23747_);
  and (_11689_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  or (_03164_, _11689_, _11688_);
  and (_11691_, _10347_, _23707_);
  and (_11692_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  or (_03168_, _11692_, _11691_);
  and (_11693_, _24766_, _23656_);
  not (_11695_, _11693_);
  and (_11697_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_11699_, _11693_, _23898_);
  or (_03175_, _11699_, _11697_);
  and (_11700_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_11701_, _11693_, _23747_);
  or (_03177_, _11701_, _11700_);
  and (_11702_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_11703_, _11693_, _23946_);
  or (_03194_, _11703_, _11702_);
  and (_11705_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_11706_, _11693_, _23707_);
  or (_03199_, _11706_, _11705_);
  and (_11708_, _02284_, _23898_);
  and (_11709_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  or (_27116_, _11709_, _11708_);
  and (_11712_, _04811_, _23898_);
  and (_11713_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or (_03209_, _11713_, _11712_);
  and (_11714_, _02302_, _24050_);
  and (_11716_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_03211_, _11716_, _11714_);
  and (_11717_, _02302_, _23824_);
  and (_11719_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_03222_, _11719_, _11717_);
  and (_11720_, _02374_, _23707_);
  and (_11722_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  or (_03225_, _11722_, _11720_);
  and (_11725_, _03339_, _23946_);
  and (_11727_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_03227_, _11727_, _11725_);
  and (_11729_, _24766_, _23752_);
  not (_11730_, _11729_);
  and (_11731_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and (_11732_, _11729_, _23778_);
  or (_03231_, _11732_, _11731_);
  and (_11735_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  and (_11736_, _11729_, _23824_);
  or (_03233_, _11736_, _11735_);
  and (_11737_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  and (_11739_, _11729_, _23946_);
  or (_03244_, _11739_, _11737_);
  and (_11740_, _04917_, _24050_);
  and (_11741_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_27110_, _11741_, _11740_);
  and (_11742_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and (_11743_, _11729_, _24050_);
  or (_27026_, _11743_, _11742_);
  and (_11744_, _07471_, _23747_);
  and (_11745_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  or (_03270_, _11745_, _11744_);
  and (_11746_, _24766_, _24329_);
  not (_11747_, _11746_);
  and (_11748_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_11749_, _11746_, _23778_);
  or (_03282_, _11749_, _11748_);
  and (_11750_, _05445_, _23649_);
  and (_11751_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  or (_03287_, _11751_, _11750_);
  and (_11752_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_11753_, _11746_, _23898_);
  or (_03289_, _11753_, _11752_);
  and (_11756_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_11757_, _11746_, _23649_);
  or (_03291_, _11757_, _11756_);
  and (_11760_, _02374_, _23824_);
  and (_11761_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or (_03294_, _11761_, _11760_);
  and (_11763_, _09913_, _23946_);
  and (_11764_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_03304_, _11764_, _11763_);
  and (_11765_, _07536_, _23707_);
  and (_11766_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or (_03310_, _11766_, _11765_);
  and (_11767_, _05180_, _24050_);
  and (_11768_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_27133_, _11768_, _11767_);
  and (_11769_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_11770_, _11746_, _23946_);
  or (_03326_, _11770_, _11769_);
  and (_11771_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_11772_, _11746_, _23707_);
  or (_27030_, _11772_, _11771_);
  and (_11773_, _08167_, _23707_);
  and (_11774_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or (_03333_, _11774_, _11773_);
  and (_11775_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  and (_11776_, _04748_, _23778_);
  or (_03341_, _11776_, _11775_);
  and (_11777_, _10347_, _23778_);
  and (_11778_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  or (_03346_, _11778_, _11777_);
  and (_11779_, _04797_, _23778_);
  and (_11780_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_03357_, _11780_, _11779_);
  and (_11781_, _01810_, _23898_);
  and (_11782_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_03362_, _11782_, _11781_);
  and (_11784_, _24371_, _23649_);
  and (_11785_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_03365_, _11785_, _11784_);
  and (_11786_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  and (_11788_, _06888_, _23707_);
  or (_03371_, _11788_, _11786_);
  and (_11789_, _07471_, _23707_);
  and (_11790_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or (_03391_, _11790_, _11789_);
  and (_11794_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  and (_11796_, _06888_, _24050_);
  or (_03398_, _11796_, _11794_);
  and (_11798_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_11799_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or (_11800_, _11799_, _11798_);
  and (_11801_, _11800_, _02445_);
  and (_11802_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_11804_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or (_11805_, _11804_, _11802_);
  and (_11806_, _11805_, _02393_);
  or (_11807_, _11806_, _11801_);
  or (_11808_, _11807_, _02459_);
  and (_11809_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_11810_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or (_11811_, _11810_, _11809_);
  and (_11812_, _11811_, _02445_);
  and (_11813_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_11814_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or (_11815_, _11814_, _11813_);
  and (_11816_, _11815_, _02393_);
  or (_11818_, _11816_, _11812_);
  or (_11819_, _11818_, _02421_);
  and (_11820_, _11819_, _02458_);
  and (_11821_, _11820_, _11808_);
  or (_11822_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or (_11823_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_11824_, _11823_, _02393_);
  and (_11825_, _11824_, _11822_);
  or (_11826_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or (_11827_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_11829_, _11827_, _02445_);
  and (_11831_, _11829_, _11826_);
  or (_11832_, _11831_, _11825_);
  or (_11833_, _11832_, _02459_);
  or (_11835_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or (_11836_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_11837_, _11836_, _02393_);
  and (_11838_, _11837_, _11835_);
  or (_11839_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or (_11840_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_11841_, _11840_, _02445_);
  and (_11842_, _11841_, _11839_);
  or (_11843_, _11842_, _11838_);
  or (_11844_, _11843_, _02421_);
  and (_11845_, _11844_, _02414_);
  and (_11846_, _11845_, _11833_);
  or (_11847_, _11846_, _11821_);
  or (_11848_, _11847_, _02398_);
  and (_11850_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and (_11851_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_11852_, _11851_, _02393_);
  or (_11854_, _11852_, _11850_);
  and (_11856_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and (_11858_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_11860_, _11858_, _02445_);
  or (_11861_, _11860_, _11856_);
  and (_11862_, _11861_, _11854_);
  or (_11864_, _11862_, _02459_);
  and (_11865_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and (_11866_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_11868_, _11866_, _02393_);
  or (_11869_, _11868_, _11865_);
  and (_11870_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and (_11871_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_11873_, _11871_, _02445_);
  or (_11874_, _11873_, _11870_);
  and (_11875_, _11874_, _11869_);
  or (_11876_, _11875_, _02421_);
  and (_11877_, _11876_, _02458_);
  and (_11879_, _11877_, _11864_);
  or (_11880_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_11881_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and (_11883_, _11881_, _11880_);
  or (_11885_, _11883_, _02445_);
  or (_11886_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_11887_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and (_11888_, _11887_, _11886_);
  or (_11889_, _11888_, _02393_);
  and (_11890_, _11889_, _11885_);
  or (_11892_, _11890_, _02459_);
  or (_11893_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_11894_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and (_11895_, _11894_, _11893_);
  or (_11896_, _11895_, _02445_);
  or (_11897_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_11898_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and (_11899_, _11898_, _11897_);
  or (_11900_, _11899_, _02393_);
  and (_11901_, _11900_, _11896_);
  or (_11902_, _11901_, _02421_);
  and (_11903_, _11902_, _02414_);
  and (_11904_, _11903_, _11892_);
  or (_11905_, _11904_, _11879_);
  or (_11906_, _11905_, _02496_);
  and (_11907_, _11906_, _02546_);
  and (_11908_, _11907_, _11848_);
  and (_11909_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_11910_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_11912_, _11910_, _11909_);
  and (_11913_, _11912_, _02393_);
  and (_11914_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and (_11915_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or (_11916_, _11915_, _11914_);
  and (_11917_, _11916_, _02445_);
  or (_11918_, _11917_, _11913_);
  and (_11919_, _11918_, _02421_);
  and (_11920_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_11921_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or (_11922_, _11921_, _11920_);
  and (_11923_, _11922_, _02393_);
  and (_11925_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_11926_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_11927_, _11926_, _11925_);
  and (_11928_, _11927_, _02445_);
  or (_11929_, _11928_, _11923_);
  and (_11930_, _11929_, _02459_);
  or (_11931_, _11930_, _11919_);
  and (_11932_, _11931_, _02458_);
  or (_11933_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_11934_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and (_11935_, _11934_, _11933_);
  and (_11936_, _11935_, _02393_);
  or (_11937_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or (_11938_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_11939_, _11938_, _11937_);
  and (_11940_, _11939_, _02445_);
  or (_11941_, _11940_, _11936_);
  and (_11942_, _11941_, _02421_);
  or (_11943_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_11944_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and (_11945_, _11944_, _11943_);
  and (_11946_, _11945_, _02393_);
  or (_11947_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_11948_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_11949_, _11948_, _11947_);
  and (_11950_, _11949_, _02445_);
  or (_11951_, _11950_, _11946_);
  and (_11952_, _11951_, _02459_);
  or (_11953_, _11952_, _11942_);
  and (_11955_, _11953_, _02414_);
  or (_11956_, _11955_, _11932_);
  and (_11957_, _11956_, _02398_);
  and (_11958_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  and (_11959_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  or (_11960_, _11959_, _11958_);
  and (_11961_, _11960_, _02393_);
  and (_11963_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  and (_11965_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  or (_11966_, _11965_, _11963_);
  and (_11967_, _11966_, _02445_);
  or (_11968_, _11967_, _11961_);
  and (_11969_, _11968_, _02421_);
  and (_11970_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  and (_11971_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  or (_11972_, _11971_, _11970_);
  and (_11973_, _11972_, _02393_);
  and (_11974_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  and (_11975_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  or (_11976_, _11975_, _11974_);
  and (_11977_, _11976_, _02445_);
  or (_11978_, _11977_, _11973_);
  and (_11979_, _11978_, _02459_);
  or (_11980_, _11979_, _11969_);
  and (_11981_, _11980_, _02458_);
  or (_11982_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  or (_11983_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  and (_11984_, _11983_, _11982_);
  and (_11985_, _11984_, _02393_);
  or (_11986_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  or (_11988_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  and (_11989_, _11988_, _11986_);
  and (_11990_, _11989_, _02445_);
  or (_11991_, _11990_, _11985_);
  and (_11992_, _11991_, _02421_);
  or (_11993_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  or (_11994_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  and (_11995_, _11994_, _11993_);
  and (_11996_, _11995_, _02393_);
  or (_11997_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  or (_11999_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  and (_12000_, _11999_, _11997_);
  and (_12001_, _12000_, _02445_);
  or (_12003_, _12001_, _11996_);
  and (_12004_, _12003_, _02459_);
  or (_12005_, _12004_, _11992_);
  and (_12006_, _12005_, _02414_);
  or (_12007_, _12006_, _11981_);
  and (_12008_, _12007_, _02496_);
  or (_12010_, _12008_, _11957_);
  and (_12011_, _12010_, _02400_);
  or (_12012_, _12011_, _11908_);
  and (_12013_, _12012_, _02646_);
  or (_12014_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_12015_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and (_12016_, _12015_, _02445_);
  and (_12017_, _12016_, _12014_);
  or (_12018_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_12019_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and (_12020_, _12019_, _02393_);
  and (_12021_, _12020_, _12018_);
  or (_12023_, _12021_, _12017_);
  and (_12025_, _12023_, _02459_);
  or (_12027_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_12029_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and (_12030_, _12029_, _02445_);
  and (_12031_, _12030_, _12027_);
  or (_12032_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_12033_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and (_12034_, _12033_, _02393_);
  and (_12036_, _12034_, _12032_);
  or (_12038_, _12036_, _12031_);
  and (_12039_, _12038_, _02421_);
  or (_12041_, _12039_, _12025_);
  and (_12043_, _12041_, _02414_);
  and (_12045_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and (_12046_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_12047_, _12046_, _12045_);
  and (_12049_, _12047_, _02393_);
  and (_12051_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and (_12053_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_12055_, _12053_, _12051_);
  and (_12057_, _12055_, _02445_);
  or (_12058_, _12057_, _12049_);
  and (_12059_, _12058_, _02459_);
  and (_12061_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and (_12062_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_12064_, _12062_, _12061_);
  and (_12065_, _12064_, _02393_);
  and (_12067_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and (_12069_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_12071_, _12069_, _12067_);
  and (_12073_, _12071_, _02445_);
  or (_12074_, _12073_, _12065_);
  and (_12075_, _12074_, _02421_);
  or (_12076_, _12075_, _12059_);
  and (_12077_, _12076_, _02458_);
  or (_12078_, _12077_, _12043_);
  and (_12079_, _12078_, _02496_);
  or (_12080_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_12081_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_12082_, _12081_, _12080_);
  and (_12083_, _12082_, _02393_);
  or (_12084_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_12085_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and (_12087_, _12085_, _12084_);
  and (_12088_, _12087_, _02445_);
  or (_12089_, _12088_, _12083_);
  and (_12090_, _12089_, _02459_);
  or (_12091_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or (_12092_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and (_12093_, _12092_, _12091_);
  and (_12094_, _12093_, _02393_);
  or (_12095_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or (_12096_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_12097_, _12096_, _12095_);
  and (_12098_, _12097_, _02445_);
  or (_12099_, _12098_, _12094_);
  and (_12100_, _12099_, _02421_);
  or (_12102_, _12100_, _12090_);
  and (_12103_, _12102_, _02414_);
  and (_12104_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_12106_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or (_12108_, _12106_, _12104_);
  and (_12110_, _12108_, _02393_);
  and (_12112_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_12114_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_12115_, _12114_, _12112_);
  and (_12117_, _12115_, _02445_);
  or (_12118_, _12117_, _12110_);
  and (_12119_, _12118_, _02459_);
  and (_12120_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_12121_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or (_12122_, _12121_, _12120_);
  and (_12123_, _12122_, _02393_);
  and (_12124_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and (_12125_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_12126_, _12125_, _12124_);
  and (_12127_, _12126_, _02445_);
  or (_12128_, _12127_, _12123_);
  and (_12129_, _12128_, _02421_);
  or (_12130_, _12129_, _12119_);
  and (_12131_, _12130_, _02458_);
  or (_12132_, _12131_, _12103_);
  and (_12133_, _12132_, _02398_);
  or (_12134_, _12133_, _12079_);
  and (_12135_, _12134_, _02400_);
  and (_12136_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_12137_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_12138_, _12137_, _12136_);
  and (_12140_, _12138_, _02393_);
  and (_12141_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and (_12142_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_12143_, _12142_, _12141_);
  and (_12144_, _12143_, _02445_);
  or (_12145_, _12144_, _12140_);
  or (_12146_, _12145_, _02459_);
  and (_12147_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and (_12148_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_12149_, _12148_, _12147_);
  and (_12150_, _12149_, _02393_);
  and (_12151_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and (_12152_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_12153_, _12152_, _12151_);
  and (_12154_, _12153_, _02445_);
  or (_12155_, _12154_, _12150_);
  or (_12156_, _12155_, _02421_);
  and (_12157_, _12156_, _02458_);
  and (_12158_, _12157_, _12146_);
  or (_12159_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_12160_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_12161_, _12160_, _12159_);
  and (_12162_, _12161_, _02393_);
  or (_12163_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_12164_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and (_12165_, _12164_, _12163_);
  and (_12166_, _12165_, _02445_);
  or (_12167_, _12166_, _12162_);
  or (_12168_, _12167_, _02459_);
  or (_12169_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_12171_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_12172_, _12171_, _12169_);
  and (_12173_, _12172_, _02393_);
  or (_12174_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_12175_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and (_12176_, _12175_, _12174_);
  and (_12177_, _12176_, _02445_);
  or (_12178_, _12177_, _12173_);
  or (_12179_, _12178_, _02421_);
  and (_12180_, _12179_, _02414_);
  and (_12181_, _12180_, _12168_);
  or (_12182_, _12181_, _12158_);
  and (_12183_, _12182_, _02398_);
  and (_12184_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and (_12186_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_12187_, _12186_, _12184_);
  and (_12188_, _12187_, _02393_);
  and (_12189_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and (_12190_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_12191_, _12190_, _12189_);
  and (_12193_, _12191_, _02445_);
  or (_12194_, _12193_, _12188_);
  or (_12195_, _12194_, _02459_);
  and (_12196_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and (_12197_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_12198_, _12197_, _12196_);
  and (_12199_, _12198_, _02393_);
  and (_12200_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and (_12201_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_12202_, _12201_, _12200_);
  and (_12203_, _12202_, _02445_);
  or (_12204_, _12203_, _12199_);
  or (_12205_, _12204_, _02421_);
  and (_12206_, _12205_, _02458_);
  and (_12207_, _12206_, _12195_);
  or (_12208_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_12209_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and (_12210_, _12209_, _02445_);
  and (_12211_, _12210_, _12208_);
  or (_12212_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_12213_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and (_12214_, _12213_, _02393_);
  and (_12215_, _12214_, _12212_);
  or (_12216_, _12215_, _12211_);
  or (_12217_, _12216_, _02459_);
  or (_12218_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_12219_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and (_12220_, _12219_, _02445_);
  and (_12221_, _12220_, _12218_);
  or (_12222_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_12225_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and (_12227_, _12225_, _02393_);
  and (_12229_, _12227_, _12222_);
  or (_12231_, _12229_, _12221_);
  or (_12233_, _12231_, _02421_);
  and (_12235_, _12233_, _02414_);
  and (_12236_, _12235_, _12217_);
  or (_12238_, _12236_, _12207_);
  and (_12240_, _12238_, _02496_);
  or (_12242_, _12240_, _12183_);
  and (_12244_, _12242_, _02546_);
  or (_12246_, _12244_, _12135_);
  and (_12248_, _12246_, _02405_);
  or (_12250_, _12248_, _12013_);
  and (_12251_, _12250_, _26777_);
  and (_12253_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and (_12255_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_12257_, _12255_, _12253_);
  and (_12259_, _12257_, _02393_);
  and (_12261_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and (_12262_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_12263_, _12262_, _12261_);
  and (_12265_, _12263_, _02445_);
  or (_12267_, _12265_, _12259_);
  and (_12269_, _12267_, _02421_);
  and (_12270_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and (_12271_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_12272_, _12271_, _12270_);
  and (_12274_, _12272_, _02393_);
  and (_12275_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and (_12276_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_12278_, _12276_, _12275_);
  and (_12279_, _12278_, _02445_);
  or (_12281_, _12279_, _12274_);
  and (_12283_, _12281_, _02459_);
  or (_12285_, _12283_, _12269_);
  and (_12286_, _12285_, _02458_);
  or (_12287_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_12289_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and (_12291_, _12289_, _12287_);
  and (_12293_, _12291_, _02393_);
  or (_12295_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_12296_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and (_12297_, _12296_, _12295_);
  and (_12298_, _12297_, _02445_);
  or (_12299_, _12298_, _12293_);
  and (_12300_, _12299_, _02421_);
  or (_12301_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_12302_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and (_12303_, _12302_, _12301_);
  and (_12304_, _12303_, _02393_);
  or (_12305_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_12306_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and (_12307_, _12306_, _12305_);
  and (_12308_, _12307_, _02445_);
  or (_12309_, _12308_, _12304_);
  and (_12310_, _12309_, _02459_);
  or (_12311_, _12310_, _12300_);
  and (_12312_, _12311_, _02414_);
  or (_12313_, _12312_, _12286_);
  and (_12314_, _12313_, _02398_);
  and (_12315_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_12316_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_12317_, _12316_, _12315_);
  and (_12318_, _12317_, _02393_);
  and (_12319_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_12320_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_12321_, _12320_, _12319_);
  and (_12322_, _12321_, _02445_);
  or (_12323_, _12322_, _12318_);
  and (_12324_, _12323_, _02421_);
  and (_12325_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_12326_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_12327_, _12326_, _12325_);
  and (_12328_, _12327_, _02393_);
  and (_12329_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_12330_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_12331_, _12330_, _12329_);
  and (_12332_, _12331_, _02445_);
  or (_12333_, _12332_, _12328_);
  and (_12334_, _12333_, _02459_);
  or (_12335_, _12334_, _12324_);
  and (_12336_, _12335_, _02458_);
  or (_12337_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_12338_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_12339_, _12338_, _02445_);
  and (_12340_, _12339_, _12337_);
  or (_12341_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_12342_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_12343_, _12342_, _02393_);
  and (_12345_, _12343_, _12341_);
  or (_12346_, _12345_, _12340_);
  and (_12347_, _12346_, _02421_);
  or (_12348_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_12349_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_12350_, _12349_, _02445_);
  and (_12351_, _12350_, _12348_);
  or (_12352_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_12353_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_12354_, _12353_, _02393_);
  and (_12355_, _12354_, _12352_);
  or (_12356_, _12355_, _12351_);
  and (_12357_, _12356_, _02459_);
  or (_12358_, _12357_, _12347_);
  and (_12359_, _12358_, _02414_);
  or (_12360_, _12359_, _12336_);
  and (_12361_, _12360_, _02496_);
  or (_12362_, _12361_, _12314_);
  and (_12363_, _12362_, _02400_);
  and (_12364_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and (_12365_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_12366_, _12365_, _12364_);
  and (_12367_, _12366_, _02393_);
  and (_12368_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and (_12369_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_12370_, _12369_, _12368_);
  and (_12371_, _12370_, _02445_);
  or (_12372_, _12371_, _12367_);
  or (_12373_, _12372_, _02459_);
  and (_12374_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and (_12375_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_12376_, _12375_, _12374_);
  and (_12377_, _12376_, _02393_);
  and (_12378_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and (_12379_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_12380_, _12379_, _12378_);
  and (_12381_, _12380_, _02445_);
  or (_12382_, _12381_, _12377_);
  or (_12383_, _12382_, _02421_);
  and (_12384_, _12383_, _02458_);
  and (_12385_, _12384_, _12373_);
  or (_12386_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_12387_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and (_12388_, _12387_, _02445_);
  and (_12389_, _12388_, _12386_);
  or (_12390_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_12391_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and (_12392_, _12391_, _02393_);
  and (_12393_, _12392_, _12390_);
  or (_12394_, _12393_, _12389_);
  or (_12396_, _12394_, _02459_);
  or (_12397_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_12398_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and (_12399_, _12398_, _02445_);
  and (_12400_, _12399_, _12397_);
  or (_12401_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_12402_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and (_12403_, _12402_, _02393_);
  and (_12404_, _12403_, _12401_);
  or (_12405_, _12404_, _12400_);
  or (_12406_, _12405_, _02421_);
  and (_12407_, _12406_, _02414_);
  and (_12408_, _12407_, _12396_);
  or (_12409_, _12408_, _12385_);
  and (_12410_, _12409_, _02496_);
  and (_12411_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and (_12412_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_12413_, _12412_, _12411_);
  and (_12414_, _12413_, _02393_);
  and (_12415_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and (_12416_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_12417_, _12416_, _12415_);
  and (_12418_, _12417_, _02445_);
  or (_12419_, _12418_, _12414_);
  or (_12420_, _12419_, _02459_);
  and (_12421_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and (_12422_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_12423_, _12422_, _12421_);
  and (_12424_, _12423_, _02393_);
  and (_12425_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and (_12426_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_12427_, _12426_, _12425_);
  and (_12428_, _12427_, _02445_);
  or (_12429_, _12428_, _12424_);
  or (_12430_, _12429_, _02421_);
  and (_12431_, _12430_, _02458_);
  and (_12432_, _12431_, _12420_);
  or (_12433_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_12434_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and (_12435_, _12434_, _12433_);
  and (_12436_, _12435_, _02393_);
  or (_12437_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_12438_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and (_12439_, _12438_, _12437_);
  and (_12440_, _12439_, _02445_);
  or (_12441_, _12440_, _12436_);
  or (_12442_, _12441_, _02459_);
  or (_12443_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_12444_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and (_12445_, _12444_, _12443_);
  and (_12446_, _12445_, _02393_);
  or (_12447_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_12448_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and (_12449_, _12448_, _12447_);
  and (_12450_, _12449_, _02445_);
  or (_12451_, _12450_, _12446_);
  or (_12452_, _12451_, _02421_);
  and (_12453_, _12452_, _02414_);
  and (_12454_, _12453_, _12442_);
  or (_12455_, _12454_, _12432_);
  and (_12456_, _12455_, _02398_);
  or (_12457_, _12456_, _12410_);
  and (_12458_, _12457_, _02546_);
  or (_12459_, _12458_, _12363_);
  and (_12460_, _12459_, _02646_);
  or (_12461_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_12462_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and (_12463_, _12462_, _02445_);
  and (_12464_, _12463_, _12461_);
  or (_12465_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or (_12466_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and (_12467_, _12466_, _02393_);
  and (_12468_, _12467_, _12465_);
  or (_12469_, _12468_, _12464_);
  and (_12470_, _12469_, _02459_);
  or (_12471_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_12472_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and (_12473_, _12472_, _02445_);
  and (_12474_, _12473_, _12471_);
  or (_12475_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or (_12476_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and (_12478_, _12476_, _02393_);
  and (_12479_, _12478_, _12475_);
  or (_12480_, _12479_, _12474_);
  and (_12481_, _12480_, _02421_);
  or (_12482_, _12481_, _12470_);
  and (_12483_, _12482_, _02414_);
  and (_12484_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and (_12485_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or (_12486_, _12485_, _12484_);
  and (_12487_, _12486_, _02393_);
  and (_12488_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and (_12489_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or (_12490_, _12489_, _12488_);
  and (_12491_, _12490_, _02445_);
  or (_12492_, _12491_, _12487_);
  and (_12493_, _12492_, _02459_);
  and (_12494_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and (_12495_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or (_12496_, _12495_, _12494_);
  and (_12497_, _12496_, _02393_);
  and (_12498_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and (_12499_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_12500_, _12499_, _12498_);
  and (_12501_, _12500_, _02445_);
  or (_12502_, _12501_, _12497_);
  and (_12503_, _12502_, _02421_);
  or (_12504_, _12503_, _12493_);
  and (_12505_, _12504_, _02458_);
  or (_12506_, _12505_, _12483_);
  and (_12508_, _12506_, _02496_);
  or (_12510_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_12511_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and (_12512_, _12511_, _12510_);
  and (_12513_, _12512_, _02393_);
  or (_12514_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_12515_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and (_12516_, _12515_, _12514_);
  and (_12517_, _12516_, _02445_);
  or (_12518_, _12517_, _12513_);
  and (_12519_, _12518_, _02459_);
  or (_12520_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_12521_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and (_12522_, _12521_, _12520_);
  and (_12523_, _12522_, _02393_);
  or (_12524_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_12525_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and (_12526_, _12525_, _12524_);
  and (_12527_, _12526_, _02445_);
  or (_12528_, _12527_, _12523_);
  and (_12530_, _12528_, _02421_);
  or (_12531_, _12530_, _12519_);
  and (_12532_, _12531_, _02414_);
  and (_12533_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and (_12534_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_12535_, _12534_, _12533_);
  and (_12536_, _12535_, _02393_);
  and (_12537_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and (_12538_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_12539_, _12538_, _12537_);
  and (_12541_, _12539_, _02445_);
  or (_12542_, _12541_, _12536_);
  and (_12544_, _12542_, _02459_);
  and (_12546_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and (_12547_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_12548_, _12547_, _12546_);
  and (_12549_, _12548_, _02393_);
  and (_12550_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and (_12551_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_12552_, _12551_, _12550_);
  and (_12553_, _12552_, _02445_);
  or (_12554_, _12553_, _12549_);
  and (_12555_, _12554_, _02421_);
  or (_12556_, _12555_, _12544_);
  and (_12557_, _12556_, _02458_);
  or (_12558_, _12557_, _12532_);
  and (_12559_, _12558_, _02398_);
  or (_12560_, _12559_, _12508_);
  and (_12561_, _12560_, _02400_);
  and (_12562_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and (_12563_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_12564_, _12563_, _12562_);
  and (_12566_, _12564_, _02393_);
  and (_12567_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and (_12568_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_12570_, _12568_, _12567_);
  and (_12571_, _12570_, _02445_);
  or (_12572_, _12571_, _12566_);
  or (_12573_, _12572_, _02459_);
  and (_12574_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and (_12575_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_12576_, _12575_, _12574_);
  and (_12577_, _12576_, _02393_);
  and (_12578_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and (_12579_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_12580_, _12579_, _12578_);
  and (_12581_, _12580_, _02445_);
  or (_12582_, _12581_, _12577_);
  or (_12583_, _12582_, _02421_);
  and (_12584_, _12583_, _02458_);
  and (_12585_, _12584_, _12573_);
  or (_12587_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_12588_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and (_12589_, _12588_, _12587_);
  and (_12590_, _12589_, _02393_);
  or (_12591_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_12592_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and (_12593_, _12592_, _12591_);
  and (_12594_, _12593_, _02445_);
  or (_12595_, _12594_, _12590_);
  or (_12596_, _12595_, _02459_);
  or (_12597_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_12598_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and (_12599_, _12598_, _12597_);
  and (_12600_, _12599_, _02393_);
  or (_12601_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_12602_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and (_12603_, _12602_, _12601_);
  and (_12604_, _12603_, _02445_);
  or (_12605_, _12604_, _12600_);
  or (_12606_, _12605_, _02421_);
  and (_12607_, _12606_, _02414_);
  and (_12608_, _12607_, _12596_);
  or (_12609_, _12608_, _12585_);
  and (_12610_, _12609_, _02398_);
  and (_12611_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and (_12612_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_12614_, _12612_, _12611_);
  and (_12616_, _12614_, _02393_);
  and (_12618_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and (_12619_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_12620_, _12619_, _12618_);
  and (_12621_, _12620_, _02445_);
  or (_12622_, _12621_, _12616_);
  or (_12623_, _12622_, _02459_);
  and (_12624_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and (_12625_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_12626_, _12625_, _12624_);
  and (_12627_, _12626_, _02393_);
  and (_12628_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and (_12629_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_12630_, _12629_, _12628_);
  and (_12631_, _12630_, _02445_);
  or (_12633_, _12631_, _12627_);
  or (_12634_, _12633_, _02421_);
  and (_12635_, _12634_, _02458_);
  and (_12636_, _12635_, _12623_);
  or (_12637_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_12638_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and (_12639_, _12638_, _02445_);
  and (_12640_, _12639_, _12637_);
  or (_12641_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_12642_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and (_12643_, _12642_, _02393_);
  and (_12644_, _12643_, _12641_);
  or (_12645_, _12644_, _12640_);
  or (_12646_, _12645_, _02459_);
  or (_12647_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_12648_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and (_12649_, _12648_, _02445_);
  and (_12650_, _12649_, _12647_);
  or (_12651_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_12652_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and (_12653_, _12652_, _02393_);
  and (_12654_, _12653_, _12651_);
  or (_12655_, _12654_, _12650_);
  or (_12656_, _12655_, _02421_);
  and (_12657_, _12656_, _02414_);
  and (_12658_, _12657_, _12646_);
  or (_12659_, _12658_, _12636_);
  and (_12660_, _12659_, _02496_);
  or (_12661_, _12660_, _12610_);
  and (_12662_, _12661_, _02546_);
  or (_12663_, _12662_, _12561_);
  and (_12664_, _12663_, _02405_);
  or (_12665_, _12664_, _12460_);
  and (_12666_, _12665_, _02444_);
  or (_12667_, _12666_, _12251_);
  or (_12668_, _12667_, _02443_);
  or (_12669_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_12670_, _12669_, _22762_);
  and (_03400_, _12670_, _12668_);
  not (_12671_, _02077_);
  or (_12673_, _12671_, _23892_);
  not (_12675_, _02073_);
  and (_12676_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_12677_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_12678_, _12677_, _12676_);
  or (_12680_, _12678_, _02077_);
  and (_12682_, _12680_, _12675_);
  and (_12683_, _12682_, _12673_);
  and (_12684_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_12685_, _12684_, _12683_);
  and (_03406_, _12685_, _22762_);
  or (_12686_, _12675_, _23642_);
  not (_12687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_12688_, _02078_, _12687_);
  and (_12689_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_12690_, _12689_, _12688_);
  or (_12691_, _12690_, _02073_);
  and (_12692_, _12691_, _22762_);
  and (_03409_, _12692_, _12686_);
  and (_12693_, _02284_, _23824_);
  and (_12694_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  or (_27117_, _12694_, _12693_);
  and (_12695_, _03339_, _24050_);
  and (_12696_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_03418_, _12696_, _12695_);
  and (_12697_, _02374_, _23747_);
  and (_12698_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  or (_03433_, _12698_, _12697_);
  and (_12699_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  and (_12700_, _06888_, _23778_);
  or (_03436_, _12700_, _12699_);
  and (_12701_, _05180_, _23707_);
  and (_12702_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_03439_, _12702_, _12701_);
  and (_12703_, _04797_, _23898_);
  and (_12705_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_03441_, _12705_, _12703_);
  or (_12707_, _02009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_12708_, _02009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_12709_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_12710_, _12709_, _01996_);
  nand (_12712_, _12710_, _12708_);
  and (_12713_, _12712_, _12707_);
  or (_12714_, _12713_, _02001_);
  or (_12715_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_12716_, _12715_, _01979_);
  and (_12718_, _12716_, _12714_);
  and (_12719_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_12721_, _01977_, _24685_);
  or (_12722_, _12721_, _12719_);
  or (_12723_, _12722_, _12718_);
  and (_03444_, _12723_, _22762_);
  and (_12724_, _08360_, _24050_);
  and (_12725_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or (_03448_, _12725_, _12724_);
  and (_12726_, _08198_, _23946_);
  and (_12727_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_03453_, _12727_, _12726_);
  and (_12728_, _06886_, _23986_);
  not (_12729_, _12728_);
  and (_12730_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  and (_12732_, _12728_, _23707_);
  or (_03463_, _12732_, _12730_);
  and (_12733_, _23986_, _23664_);
  and (_12734_, _12733_, _23649_);
  not (_12735_, _12733_);
  and (_12737_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  or (_27085_, _12737_, _12734_);
  and (_12738_, _01977_, _23642_);
  and (_12739_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_12740_, _12739_, _02041_);
  nand (_12742_, _02009_, _01983_);
  nor (_12743_, _12742_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_12744_, _12742_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_12745_, _12744_, _02001_);
  or (_12746_, _12745_, _12743_);
  or (_12747_, _12746_, _12740_);
  or (_12748_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_12749_, _12748_, _01979_);
  and (_12750_, _12749_, _12747_);
  and (_12751_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_12752_, _12751_, _12750_);
  or (_12753_, _12752_, _12738_);
  and (_03477_, _12753_, _22762_);
  not (_12754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_12755_, _02025_, _12754_);
  nand (_12756_, _12755_, _02041_);
  not (_12757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand (_12758_, _02009_, _01989_);
  and (_12759_, _12758_, _12757_);
  nor (_12760_, _12758_, _12757_);
  or (_12761_, _12760_, _12759_);
  and (_12762_, _12761_, _02002_);
  nand (_12763_, _12762_, _12756_);
  not (_12764_, _01979_);
  and (_12765_, _02001_, _12754_);
  nor (_12766_, _12765_, _12764_);
  and (_12767_, _12766_, _12763_);
  and (_12768_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_12769_, _12768_, _12767_);
  and (_12770_, _01978_, _23816_);
  or (_12771_, _12770_, _12769_);
  and (_03486_, _12771_, _22762_);
  and (_12772_, _08307_, _24291_);
  nand (_12773_, _12772_, _23594_);
  not (_12774_, _08313_);
  or (_12775_, _12772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_12776_, _12775_, _12774_);
  and (_12777_, _12776_, _12773_);
  and (_12778_, _08313_, _23816_);
  or (_12779_, _12778_, _12777_);
  and (_03500_, _12779_, _22762_);
  and (_12780_, _08799_, _23778_);
  and (_12781_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or (_03505_, _12781_, _12780_);
  and (_12782_, _24282_, _23664_);
  and (_12783_, _12782_, _23824_);
  not (_12784_, _12782_);
  and (_12785_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_03509_, _12785_, _12783_);
  and (_12786_, _24010_, _23664_);
  and (_12787_, _12786_, _23707_);
  not (_12788_, _12786_);
  and (_12789_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or (_03518_, _12789_, _12787_);
  and (_12790_, _08360_, _23946_);
  and (_12791_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or (_03524_, _12791_, _12790_);
  and (_12792_, _05350_, _23898_);
  and (_12793_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  or (_03539_, _12793_, _12792_);
  and (_12794_, _09913_, _23898_);
  and (_12795_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_03557_, _12795_, _12794_);
  and (_12796_, _25739_, _23747_);
  and (_12797_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or (_03574_, _12797_, _12796_);
  and (_12798_, _02370_, _23946_);
  and (_12799_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_03577_, _12799_, _12798_);
  and (_12800_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  and (_12801_, _06888_, _23824_);
  or (_27013_, _12801_, _12800_);
  and (_12802_, _04811_, _23778_);
  and (_12803_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or (_27066_, _12803_, _12802_);
  and (_12804_, _03300_, _23778_);
  and (_12806_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or (_03605_, _12806_, _12804_);
  and (_12807_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  and (_12808_, _06888_, _23898_);
  or (_03608_, _12808_, _12807_);
  and (_12809_, _23755_, _23707_);
  and (_12810_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or (_03613_, _12810_, _12809_);
  and (_12811_, _26110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_12812_, _12811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_12813_, _12812_, _09917_);
  and (_12814_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_12815_, _12814_, _26118_);
  nor (_12816_, _12815_, _12813_);
  nor (_12817_, _12816_, _24299_);
  and (_12818_, _24299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_12819_, _12818_, _12817_);
  and (_12820_, _12819_, _24294_);
  and (_12821_, _24293_, _23892_);
  or (_12822_, _12821_, _12820_);
  and (_03628_, _12822_, _22762_);
  and (_12823_, _24226_, _23946_);
  and (_12824_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or (_03638_, _12824_, _12823_);
  and (_12825_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and (_12826_, _25252_, _23778_);
  or (_03656_, _12826_, _12825_);
  and (_12827_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  and (_12828_, _25542_, _23747_);
  or (_03664_, _12828_, _12827_);
  and (_12829_, _24201_, _24085_);
  not (_12830_, _12829_);
  and (_12831_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and (_12832_, _12829_, _24050_);
  or (_03676_, _12832_, _12831_);
  and (_12833_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and (_12834_, _02245_, _23898_);
  or (_27035_, _12834_, _12833_);
  and (_12835_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  and (_12836_, _12728_, _23824_);
  or (_03680_, _12836_, _12835_);
  and (_12837_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  and (_12838_, _12728_, _23898_);
  or (_03683_, _12838_, _12837_);
  and (_12839_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  and (_12840_, _04748_, _24050_);
  or (_27032_, _12840_, _12839_);
  and (_12841_, _05008_, _23649_);
  and (_12842_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_03701_, _12842_, _12841_);
  and (_12843_, _05008_, _23898_);
  and (_12844_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_03703_, _12844_, _12843_);
  and (_12845_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  and (_12846_, _12728_, _23778_);
  or (_03710_, _12846_, _12845_);
  and (_12847_, _05288_, _23946_);
  and (_12848_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or (_03713_, _12848_, _12847_);
  and (_12849_, _05701_, _23747_);
  and (_12850_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_03724_, _12850_, _12849_);
  and (_12851_, _01971_, _23649_);
  and (_12852_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  or (_03742_, _12852_, _12851_);
  and (_12853_, _24050_, _23665_);
  and (_12854_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  or (_03748_, _12854_, _12853_);
  and (_12855_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and (_12856_, _06918_, _23649_);
  or (_03751_, _12856_, _12855_);
  or (_12857_, _04945_, _24591_);
  and (_12858_, _24604_, _26582_);
  and (_12859_, _26625_, _24599_);
  or (_12860_, _12859_, _12858_);
  or (_12861_, _12860_, _12857_);
  and (_12862_, _25638_, _26582_);
  and (_12863_, _24604_, _24445_);
  or (_12864_, _12863_, _12862_);
  or (_12865_, _04958_, _04982_);
  or (_12866_, _12865_, _12864_);
  or (_12867_, _12866_, _12861_);
  and (_12868_, _24556_, _24541_);
  or (_12869_, _05016_, _12868_);
  or (_12870_, _12869_, _12867_);
  or (_12871_, _04974_, _04970_);
  or (_12872_, _12871_, _04943_);
  or (_12873_, _24605_, _24586_);
  or (_12874_, _12873_, _24600_);
  or (_12875_, _02269_, _24537_);
  or (_12876_, _12875_, _12874_);
  or (_12877_, _12876_, _12872_);
  or (_12878_, _12877_, _12870_);
  and (_12879_, _12878_, _22768_);
  and (_12880_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_12881_, _12880_, _05003_);
  or (_12882_, _12881_, _12879_);
  and (_26866_[0], _12882_, _22762_);
  and (_12883_, _25748_, _24050_);
  and (_12884_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_03763_, _12884_, _12883_);
  and (_12885_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  and (_12886_, _12728_, _23946_);
  or (_03765_, _12886_, _12885_);
  and (_12887_, _05281_, _23946_);
  and (_12888_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_03768_, _12888_, _12887_);
  and (_12889_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  and (_12890_, _12728_, _23649_);
  or (_03775_, _12890_, _12889_);
  and (_12891_, _24331_, _23649_);
  and (_12892_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_03792_, _12892_, _12891_);
  and (_12893_, _24081_, _23707_);
  and (_12894_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_03802_, _12894_, _12893_);
  and (_12895_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  and (_12896_, _25252_, _23946_);
  or (_03809_, _12896_, _12895_);
  and (_12897_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_12898_, _25763_, _23649_);
  or (_27041_, _12898_, _12897_);
  not (_12899_, _25644_);
  and (_12900_, _24598_, _24567_);
  nor (_12901_, _12900_, _04981_);
  or (_26862_[1], _12901_, _12899_);
  and (_12902_, _12786_, _23778_);
  and (_12903_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or (_03846_, _12903_, _12902_);
  and (_12904_, _09913_, _23824_);
  and (_12905_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_03849_, _12905_, _12904_);
  and (_12906_, _06886_, _23069_);
  not (_12907_, _12906_);
  and (_12908_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_12909_, _12906_, _23649_);
  or (_03865_, _12909_, _12908_);
  and (_12910_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  and (_12911_, _25542_, _23649_);
  or (_03871_, _12911_, _12910_);
  or (_12912_, _04663_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_12913_, _04682_, _04666_);
  or (_12914_, _12913_, _12912_);
  and (_12915_, _12914_, _04694_);
  nor (_12916_, _04693_, _24564_);
  or (_12917_, _12916_, rst);
  or (_26863_[0], _12917_, _12915_);
  and (_12918_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and (_12919_, _12906_, _23747_);
  or (_03878_, _12919_, _12918_);
  and (_12921_, _23833_, _23778_);
  and (_12922_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_03880_, _12922_, _12921_);
  and (_12923_, _05125_, _23824_);
  and (_12924_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  or (_03883_, _12924_, _12923_);
  and (_12925_, _08799_, _23707_);
  and (_12926_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or (_03894_, _12926_, _12925_);
  and (_12927_, _05336_, _23991_);
  not (_12928_, _12927_);
  and (_12929_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_12930_, _12927_, _23747_);
  or (_03936_, _12930_, _12929_);
  and (_12931_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_12932_, _12927_, _23778_);
  or (_27103_, _12932_, _12931_);
  and (_12933_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and (_12934_, _12829_, _23946_);
  or (_03969_, _12934_, _12933_);
  and (_12935_, _05336_, _23903_);
  not (_12936_, _12935_);
  and (_12937_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_12938_, _12935_, _23649_);
  or (_27102_, _12938_, _12937_);
  and (_12939_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_12940_, _12906_, _23707_);
  or (_03980_, _12940_, _12939_);
  and (_12941_, _05336_, _24005_);
  not (_12942_, _12941_);
  and (_12943_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  and (_12944_, _12941_, _24050_);
  or (_03984_, _12944_, _12943_);
  and (_12945_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  and (_12946_, _12941_, _23649_);
  or (_03987_, _12946_, _12945_);
  and (_12947_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and (_12948_, _12829_, _23649_);
  or (_03995_, _12948_, _12947_);
  or (_12949_, _24171_, _24043_);
  and (_12951_, _24151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_12952_, _12951_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_12953_, _12951_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_12954_, _12953_, _12952_);
  nor (_12955_, _24184_, _24132_);
  nor (_12956_, _12955_, _24127_);
  and (_12957_, _12956_, _12954_);
  not (_12958_, _12956_);
  and (_12959_, _12958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_12960_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_12961_, _12960_, _24127_);
  or (_12962_, _12961_, _12959_);
  or (_12963_, _12962_, _12957_);
  or (_12964_, _12963_, _24120_);
  and (_12965_, _12964_, _22762_);
  and (_03997_, _12965_, _12949_);
  and (_12966_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_12967_, _12906_, _24050_);
  or (_04003_, _12967_, _12966_);
  and (_12968_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_12969_, _12906_, _23946_);
  or (_04007_, _12969_, _12968_);
  and (_12970_, _05336_, _23986_);
  not (_12971_, _12970_);
  and (_12972_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  and (_12973_, _12970_, _23898_);
  or (_27098_, _12973_, _12972_);
  and (_12974_, _05336_, _23069_);
  not (_12975_, _12974_);
  and (_12976_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_12977_, _12974_, _23649_);
  or (_27096_, _12977_, _12976_);
  and (_12978_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_12979_, _06918_, _23898_);
  or (_04025_, _12979_, _12978_);
  and (_12980_, _05336_, _01808_);
  not (_12981_, _12980_);
  and (_12982_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and (_12983_, _12980_, _23649_);
  or (_04031_, _12983_, _12982_);
  and (_12984_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_12985_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_12986_, _12985_, _12984_);
  and (_12987_, _12986_, _02393_);
  and (_12988_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_12989_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or (_12990_, _12989_, _12988_);
  and (_12991_, _12990_, _02445_);
  or (_12992_, _12991_, _12987_);
  and (_12993_, _12992_, _02421_);
  and (_12994_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and (_12995_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or (_12996_, _12995_, _12994_);
  and (_12997_, _12996_, _02393_);
  and (_12998_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_12999_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_13000_, _12999_, _12998_);
  and (_13001_, _13000_, _02445_);
  or (_13002_, _13001_, _12997_);
  and (_13003_, _13002_, _02459_);
  or (_13004_, _13003_, _12993_);
  and (_13005_, _13004_, _02458_);
  or (_13006_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_13007_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_13008_, _13007_, _13006_);
  and (_13009_, _13008_, _02393_);
  or (_13010_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_13011_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_13012_, _13011_, _13010_);
  and (_13013_, _13012_, _02445_);
  or (_13014_, _13013_, _13009_);
  and (_13015_, _13014_, _02421_);
  or (_13016_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_13017_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_13018_, _13017_, _13016_);
  and (_13019_, _13018_, _02393_);
  or (_13020_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or (_13021_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_13022_, _13021_, _13020_);
  and (_13023_, _13022_, _02445_);
  or (_13024_, _13023_, _13019_);
  and (_13025_, _13024_, _02459_);
  or (_13026_, _13025_, _13015_);
  and (_13027_, _13026_, _02414_);
  or (_13028_, _13027_, _13005_);
  and (_13029_, _13028_, _02398_);
  and (_13030_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and (_13031_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_13032_, _13031_, _13030_);
  and (_13033_, _13032_, _02393_);
  and (_13034_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and (_13035_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_13036_, _13035_, _13034_);
  and (_13037_, _13036_, _02445_);
  or (_13038_, _13037_, _13033_);
  and (_13039_, _13038_, _02421_);
  and (_13040_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and (_13041_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_13042_, _13041_, _13040_);
  and (_13043_, _13042_, _02393_);
  and (_13044_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_13045_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_13046_, _13045_, _13044_);
  and (_13047_, _13046_, _02445_);
  or (_13048_, _13047_, _13043_);
  and (_13049_, _13048_, _02459_);
  or (_13050_, _13049_, _13039_);
  and (_13051_, _13050_, _02458_);
  or (_13052_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_13053_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and (_13054_, _13053_, _02445_);
  and (_13055_, _13054_, _13052_);
  or (_13056_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_13057_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and (_13058_, _13057_, _02393_);
  and (_13059_, _13058_, _13056_);
  or (_13060_, _13059_, _13055_);
  and (_13061_, _13060_, _02421_);
  or (_13062_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_13063_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_13064_, _13063_, _02445_);
  and (_13065_, _13064_, _13062_);
  or (_13066_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_13067_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_13068_, _13067_, _02393_);
  and (_13069_, _13068_, _13066_);
  or (_13070_, _13069_, _13065_);
  and (_13071_, _13070_, _02459_);
  or (_13072_, _13071_, _13061_);
  and (_13073_, _13072_, _02414_);
  or (_13074_, _13073_, _13051_);
  and (_13075_, _13074_, _02496_);
  or (_13076_, _13075_, _13029_);
  and (_13077_, _13076_, _02400_);
  and (_13078_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_13079_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or (_13080_, _13079_, _13078_);
  and (_13081_, _13080_, _02393_);
  and (_13082_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_13083_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or (_13084_, _13083_, _13082_);
  and (_13085_, _13084_, _02445_);
  or (_13086_, _13085_, _13081_);
  or (_13087_, _13086_, _02459_);
  and (_13088_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_13089_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or (_13090_, _13089_, _13088_);
  and (_13091_, _13090_, _02393_);
  and (_13092_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_13093_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or (_13094_, _13093_, _13092_);
  and (_13095_, _13094_, _02445_);
  or (_13096_, _13095_, _13091_);
  or (_13097_, _13096_, _02421_);
  and (_13098_, _13097_, _02458_);
  and (_13099_, _13098_, _13087_);
  or (_13100_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or (_13101_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_13102_, _13101_, _02445_);
  and (_13103_, _13102_, _13100_);
  or (_13104_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or (_13105_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_13106_, _13105_, _02393_);
  and (_13107_, _13106_, _13104_);
  or (_13108_, _13107_, _13103_);
  or (_13109_, _13108_, _02459_);
  or (_13110_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or (_13111_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_13112_, _13111_, _02445_);
  and (_13113_, _13112_, _13110_);
  or (_13114_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or (_13115_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_13116_, _13115_, _02393_);
  and (_13117_, _13116_, _13114_);
  or (_13118_, _13117_, _13113_);
  or (_13119_, _13118_, _02421_);
  and (_13120_, _13119_, _02414_);
  and (_13121_, _13120_, _13109_);
  or (_13122_, _13121_, _13099_);
  and (_13123_, _13122_, _02496_);
  and (_13124_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and (_13125_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_13126_, _13125_, _13124_);
  and (_13127_, _13126_, _02393_);
  and (_13128_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and (_13129_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_13130_, _13129_, _13128_);
  and (_13131_, _13130_, _02445_);
  or (_13132_, _13131_, _13127_);
  or (_13133_, _13132_, _02459_);
  and (_13134_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and (_13135_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_13136_, _13135_, _13134_);
  and (_13137_, _13136_, _02393_);
  and (_13138_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and (_13139_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_13140_, _13139_, _13138_);
  and (_13141_, _13140_, _02445_);
  or (_13142_, _13141_, _13137_);
  or (_13143_, _13142_, _02421_);
  and (_13144_, _13143_, _02458_);
  and (_13145_, _13144_, _13133_);
  or (_13146_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_13147_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and (_13148_, _13147_, _13146_);
  and (_13149_, _13148_, _02393_);
  or (_13150_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_13151_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and (_13152_, _13151_, _13150_);
  and (_13153_, _13152_, _02445_);
  or (_13154_, _13153_, _13149_);
  or (_13155_, _13154_, _02459_);
  or (_13156_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_13157_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and (_13158_, _13157_, _13156_);
  and (_13159_, _13158_, _02393_);
  or (_13160_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_13161_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and (_13162_, _13161_, _13160_);
  and (_13163_, _13162_, _02445_);
  or (_13164_, _13163_, _13159_);
  or (_13165_, _13164_, _02421_);
  and (_13166_, _13165_, _02414_);
  and (_13167_, _13166_, _13155_);
  or (_13168_, _13167_, _13145_);
  and (_13169_, _13168_, _02398_);
  or (_13170_, _13169_, _13123_);
  and (_13171_, _13170_, _02546_);
  or (_13172_, _13171_, _13077_);
  and (_13173_, _13172_, _02646_);
  or (_13174_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_13175_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and (_13176_, _13175_, _02445_);
  and (_13177_, _13176_, _13174_);
  or (_13178_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_13179_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and (_13180_, _13179_, _02393_);
  and (_13181_, _13180_, _13178_);
  or (_13182_, _13181_, _13177_);
  and (_13183_, _13182_, _02459_);
  or (_13184_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_13185_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and (_13186_, _13185_, _02445_);
  and (_13187_, _13186_, _13184_);
  or (_13188_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or (_13189_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and (_13190_, _13189_, _02393_);
  and (_13191_, _13190_, _13188_);
  or (_13192_, _13191_, _13187_);
  and (_13193_, _13192_, _02421_);
  or (_13194_, _13193_, _13183_);
  and (_13195_, _13194_, _02414_);
  and (_13196_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and (_13197_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_13198_, _13197_, _13196_);
  and (_13199_, _13198_, _02393_);
  and (_13200_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and (_13201_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_13202_, _13201_, _13200_);
  and (_13203_, _13202_, _02445_);
  or (_13204_, _13203_, _13199_);
  and (_13205_, _13204_, _02459_);
  and (_13206_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and (_13207_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_13208_, _13207_, _13206_);
  and (_13209_, _13208_, _02393_);
  and (_13210_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and (_13211_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_13212_, _13211_, _13210_);
  and (_13213_, _13212_, _02445_);
  or (_13214_, _13213_, _13209_);
  and (_13215_, _13214_, _02421_);
  or (_13216_, _13215_, _13205_);
  and (_13217_, _13216_, _02458_);
  or (_13218_, _13217_, _13195_);
  and (_13219_, _13218_, _02496_);
  or (_13220_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or (_13221_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and (_13222_, _13221_, _13220_);
  and (_13223_, _13222_, _02393_);
  or (_13224_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_13225_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_13226_, _13225_, _13224_);
  and (_13227_, _13226_, _02445_);
  or (_13228_, _13227_, _13223_);
  and (_13229_, _13228_, _02459_);
  or (_13230_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_13231_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and (_13232_, _13231_, _13230_);
  and (_13233_, _13232_, _02393_);
  or (_13234_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_13235_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_13236_, _13235_, _13234_);
  and (_13237_, _13236_, _02445_);
  or (_13238_, _13237_, _13233_);
  and (_13239_, _13238_, _02421_);
  or (_13240_, _13239_, _13229_);
  and (_13241_, _13240_, _02414_);
  and (_13242_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and (_13243_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_13244_, _13243_, _13242_);
  and (_13245_, _13244_, _02393_);
  and (_13246_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_13247_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_13248_, _13247_, _13246_);
  and (_13249_, _13248_, _02445_);
  or (_13250_, _13249_, _13245_);
  and (_13251_, _13250_, _02459_);
  and (_13252_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_13253_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_13254_, _13253_, _13252_);
  and (_13255_, _13254_, _02393_);
  and (_13256_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_13257_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or (_13258_, _13257_, _13256_);
  and (_13259_, _13258_, _02445_);
  or (_13260_, _13259_, _13255_);
  and (_13261_, _13260_, _02421_);
  or (_13262_, _13261_, _13251_);
  and (_13263_, _13262_, _02458_);
  or (_13264_, _13263_, _13241_);
  and (_13265_, _13264_, _02398_);
  or (_13266_, _13265_, _13219_);
  and (_13267_, _13266_, _02400_);
  and (_13268_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and (_13269_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_13270_, _13269_, _13268_);
  and (_13271_, _13270_, _02393_);
  and (_13272_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and (_13273_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_13274_, _13273_, _13272_);
  and (_13275_, _13274_, _02445_);
  or (_13276_, _13275_, _13271_);
  or (_13277_, _13276_, _02459_);
  and (_13278_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and (_13279_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_13280_, _13279_, _13278_);
  and (_13281_, _13280_, _02393_);
  and (_13282_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_13283_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_13284_, _13283_, _13282_);
  and (_13285_, _13284_, _02445_);
  or (_13286_, _13285_, _13281_);
  or (_13287_, _13286_, _02421_);
  and (_13288_, _13287_, _02458_);
  and (_13289_, _13288_, _13277_);
  or (_13290_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_13291_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and (_13292_, _13291_, _13290_);
  and (_13293_, _13292_, _02393_);
  or (_13294_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_13295_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and (_13296_, _13295_, _13294_);
  and (_13297_, _13296_, _02445_);
  or (_13298_, _13297_, _13293_);
  or (_13299_, _13298_, _02459_);
  or (_13300_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_13301_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_13302_, _13301_, _13300_);
  and (_13303_, _13302_, _02393_);
  or (_13304_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_13305_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and (_13306_, _13305_, _13304_);
  and (_13307_, _13306_, _02445_);
  or (_13308_, _13307_, _13303_);
  or (_13309_, _13308_, _02421_);
  and (_13310_, _13309_, _02414_);
  and (_13311_, _13310_, _13299_);
  or (_13312_, _13311_, _13289_);
  and (_13313_, _13312_, _02398_);
  and (_13314_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and (_13315_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_13316_, _13315_, _13314_);
  and (_13317_, _13316_, _02393_);
  and (_13318_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and (_13319_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_13320_, _13319_, _13318_);
  and (_13321_, _13320_, _02445_);
  or (_13322_, _13321_, _13317_);
  or (_13323_, _13322_, _02459_);
  and (_13324_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and (_13325_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_13326_, _13325_, _13324_);
  and (_13327_, _13326_, _02393_);
  and (_13328_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and (_13329_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_13330_, _13329_, _13328_);
  and (_13331_, _13330_, _02445_);
  or (_13332_, _13331_, _13327_);
  or (_13333_, _13332_, _02421_);
  and (_13334_, _13333_, _02458_);
  and (_13335_, _13334_, _13323_);
  or (_13336_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_13337_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and (_13338_, _13337_, _02445_);
  and (_13339_, _13338_, _13336_);
  or (_13340_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_13341_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and (_13342_, _13341_, _02393_);
  and (_13343_, _13342_, _13340_);
  or (_13344_, _13343_, _13339_);
  or (_13345_, _13344_, _02459_);
  or (_13346_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_13347_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and (_13348_, _13347_, _02445_);
  and (_13349_, _13348_, _13346_);
  or (_13350_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_13351_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and (_13352_, _13351_, _02393_);
  and (_13353_, _13352_, _13350_);
  or (_13354_, _13353_, _13349_);
  or (_13355_, _13354_, _02421_);
  and (_13356_, _13355_, _02414_);
  and (_13357_, _13356_, _13345_);
  or (_13358_, _13357_, _13335_);
  and (_13359_, _13358_, _02496_);
  or (_13360_, _13359_, _13313_);
  and (_13361_, _13360_, _02546_);
  or (_13362_, _13361_, _13267_);
  and (_13363_, _13362_, _02405_);
  or (_13364_, _13363_, _13173_);
  and (_13365_, _13364_, _26777_);
  and (_13366_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and (_13367_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_13368_, _13367_, _13366_);
  and (_13369_, _13368_, _02393_);
  and (_13370_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and (_13371_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_13372_, _13371_, _13370_);
  and (_13373_, _13372_, _02445_);
  or (_13374_, _13373_, _13369_);
  and (_13375_, _13374_, _02421_);
  and (_13376_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and (_13377_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_13378_, _13377_, _13376_);
  and (_13379_, _13378_, _02393_);
  and (_13380_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and (_13381_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_13382_, _13381_, _13380_);
  and (_13383_, _13382_, _02445_);
  or (_13384_, _13383_, _13379_);
  and (_13385_, _13384_, _02459_);
  or (_13386_, _13385_, _02414_);
  or (_13387_, _13386_, _13375_);
  or (_13388_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_13389_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and (_13390_, _13389_, _13388_);
  and (_13391_, _13390_, _02393_);
  or (_13392_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_13393_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and (_13394_, _13393_, _13392_);
  and (_13395_, _13394_, _02445_);
  or (_13396_, _13395_, _13391_);
  and (_13397_, _13396_, _02421_);
  or (_13398_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_13399_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and (_13400_, _13399_, _13398_);
  and (_13401_, _13400_, _02393_);
  or (_13402_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_13403_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and (_13404_, _13403_, _13402_);
  and (_13405_, _13404_, _02445_);
  or (_13406_, _13405_, _13401_);
  and (_13407_, _13406_, _02459_);
  or (_13408_, _13407_, _02458_);
  or (_13409_, _13408_, _13397_);
  and (_13410_, _13409_, _13387_);
  or (_13411_, _13410_, _02496_);
  and (_13412_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_13413_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_13414_, _13413_, _13412_);
  and (_13415_, _13414_, _02393_);
  and (_13416_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_13417_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_13418_, _13417_, _13416_);
  and (_13419_, _13418_, _02445_);
  or (_13420_, _13419_, _13415_);
  and (_13421_, _13420_, _02421_);
  and (_13422_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_13423_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_13424_, _13423_, _13422_);
  and (_13425_, _13424_, _02393_);
  and (_13426_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_13427_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_13428_, _13427_, _13426_);
  and (_13429_, _13428_, _02445_);
  or (_13430_, _13429_, _13425_);
  and (_13431_, _13430_, _02459_);
  or (_13432_, _13431_, _02414_);
  or (_13433_, _13432_, _13421_);
  or (_13434_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_13435_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_13436_, _13435_, _02445_);
  and (_13437_, _13436_, _13434_);
  or (_13438_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_13439_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_13440_, _13439_, _02393_);
  and (_13441_, _13440_, _13438_);
  or (_13442_, _13441_, _13437_);
  and (_13443_, _13442_, _02421_);
  or (_13444_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_13445_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_13446_, _13445_, _02445_);
  and (_13447_, _13446_, _13444_);
  or (_13448_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_13449_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_13450_, _13449_, _02393_);
  and (_13451_, _13450_, _13448_);
  or (_13452_, _13451_, _13447_);
  and (_13453_, _13452_, _02459_);
  or (_13454_, _13453_, _02458_);
  or (_13455_, _13454_, _13443_);
  and (_13456_, _13455_, _13433_);
  or (_13457_, _13456_, _02398_);
  and (_13458_, _13457_, _13411_);
  and (_13459_, _13458_, _02400_);
  and (_13460_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and (_13461_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_13462_, _13461_, _13460_);
  and (_13463_, _13462_, _02393_);
  and (_13464_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and (_13465_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_13466_, _13465_, _13464_);
  and (_13467_, _13466_, _02445_);
  or (_13468_, _13467_, _13463_);
  or (_13469_, _13468_, _02459_);
  and (_13470_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and (_13471_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_13472_, _13471_, _13470_);
  and (_13473_, _13472_, _02393_);
  and (_13474_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and (_13475_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_13476_, _13475_, _13474_);
  and (_13477_, _13476_, _02445_);
  or (_13478_, _13477_, _13473_);
  or (_13479_, _13478_, _02421_);
  and (_13480_, _13479_, _02458_);
  and (_13481_, _13480_, _13469_);
  or (_13482_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_13483_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and (_13484_, _13483_, _02445_);
  and (_13485_, _13484_, _13482_);
  or (_13486_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_13487_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and (_13488_, _13487_, _02393_);
  and (_13489_, _13488_, _13486_);
  or (_13490_, _13489_, _13485_);
  or (_13491_, _13490_, _02459_);
  or (_13492_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_13493_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and (_13494_, _13493_, _02445_);
  and (_13495_, _13494_, _13492_);
  or (_13496_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_13497_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and (_13498_, _13497_, _02393_);
  and (_13499_, _13498_, _13496_);
  or (_13500_, _13499_, _13495_);
  or (_13501_, _13500_, _02421_);
  and (_13502_, _13501_, _02414_);
  and (_13503_, _13502_, _13491_);
  or (_13504_, _13503_, _13481_);
  or (_13505_, _13504_, _02398_);
  and (_13506_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and (_13507_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_13508_, _13507_, _13506_);
  and (_13509_, _13508_, _02393_);
  and (_13510_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and (_13511_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_13512_, _13511_, _13510_);
  and (_13513_, _13512_, _02445_);
  or (_13514_, _13513_, _13509_);
  or (_13515_, _13514_, _02459_);
  and (_13516_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and (_13517_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_13518_, _13517_, _13516_);
  and (_13519_, _13518_, _02393_);
  and (_13520_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and (_13521_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_13522_, _13521_, _13520_);
  and (_13523_, _13522_, _02445_);
  or (_13524_, _13523_, _13519_);
  or (_13525_, _13524_, _02421_);
  and (_13526_, _13525_, _02458_);
  and (_13527_, _13526_, _13515_);
  or (_13528_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_13529_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and (_13530_, _13529_, _13528_);
  and (_13531_, _13530_, _02393_);
  or (_13532_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_13533_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and (_13534_, _13533_, _13532_);
  and (_13535_, _13534_, _02445_);
  or (_13536_, _13535_, _13531_);
  or (_13537_, _13536_, _02459_);
  or (_13538_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_13539_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and (_13540_, _13539_, _13538_);
  and (_13541_, _13540_, _02393_);
  or (_13542_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_13543_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and (_13544_, _13543_, _13542_);
  and (_13545_, _13544_, _02445_);
  or (_13546_, _13545_, _13541_);
  or (_13547_, _13546_, _02421_);
  and (_13548_, _13547_, _02414_);
  and (_13549_, _13548_, _13537_);
  or (_13550_, _13549_, _13527_);
  or (_13551_, _13550_, _02496_);
  and (_13552_, _13551_, _13505_);
  and (_13553_, _13552_, _02546_);
  or (_13554_, _13553_, _13459_);
  and (_13555_, _13554_, _02646_);
  and (_13556_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and (_13557_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_13558_, _13557_, _13556_);
  and (_13559_, _13558_, _02445_);
  and (_13560_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and (_13561_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_13562_, _13561_, _13560_);
  and (_13563_, _13562_, _02393_);
  or (_13564_, _13563_, _13559_);
  or (_13565_, _13564_, _02459_);
  and (_13566_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and (_13567_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_13568_, _13567_, _13566_);
  and (_13569_, _13568_, _02445_);
  and (_13570_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and (_13571_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_13572_, _13571_, _13570_);
  and (_13573_, _13572_, _02393_);
  or (_13574_, _13573_, _13569_);
  or (_13575_, _13574_, _02421_);
  and (_13576_, _13575_, _02458_);
  and (_13577_, _13576_, _13565_);
  or (_13578_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_13579_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and (_13580_, _13579_, _02393_);
  and (_13581_, _13580_, _13578_);
  or (_13582_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_13583_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and (_13584_, _13583_, _02445_);
  and (_13585_, _13584_, _13582_);
  or (_13586_, _13585_, _13581_);
  or (_13587_, _13586_, _02459_);
  or (_13588_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_13589_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and (_13590_, _13589_, _02393_);
  and (_13591_, _13590_, _13588_);
  or (_13592_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_13593_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and (_13594_, _13593_, _02445_);
  and (_13595_, _13594_, _13592_);
  or (_13596_, _13595_, _13591_);
  or (_13597_, _13596_, _02421_);
  and (_13598_, _13597_, _02414_);
  and (_13599_, _13598_, _13587_);
  or (_13600_, _13599_, _13577_);
  or (_13601_, _13600_, _02398_);
  and (_13602_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and (_13603_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_13604_, _13603_, _02393_);
  or (_13605_, _13604_, _13602_);
  and (_13606_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and (_13607_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_13608_, _13607_, _02445_);
  or (_13609_, _13608_, _13606_);
  and (_13610_, _13609_, _13605_);
  or (_13611_, _13610_, _02459_);
  and (_13612_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and (_13613_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_13614_, _13613_, _02393_);
  or (_13615_, _13614_, _13612_);
  and (_13616_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and (_13617_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_13618_, _13617_, _02445_);
  or (_13619_, _13618_, _13616_);
  and (_13620_, _13619_, _13615_);
  or (_13621_, _13620_, _02421_);
  and (_13622_, _13621_, _02458_);
  and (_13623_, _13622_, _13611_);
  or (_13624_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_13625_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and (_13626_, _13625_, _13624_);
  or (_13627_, _13626_, _02445_);
  or (_13628_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_13629_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and (_13630_, _13629_, _13628_);
  or (_13631_, _13630_, _02393_);
  and (_13632_, _13631_, _13627_);
  or (_13633_, _13632_, _02459_);
  or (_13634_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_13635_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and (_13636_, _13635_, _13634_);
  or (_13637_, _13636_, _02445_);
  or (_13638_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_13639_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and (_13640_, _13639_, _13638_);
  or (_13641_, _13640_, _02393_);
  and (_13642_, _13641_, _13637_);
  or (_13643_, _13642_, _02421_);
  and (_13644_, _13643_, _02414_);
  and (_13645_, _13644_, _13633_);
  or (_13646_, _13645_, _13623_);
  or (_13647_, _13646_, _02496_);
  and (_13648_, _13647_, _02546_);
  and (_13649_, _13648_, _13601_);
  and (_13650_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and (_13651_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_13652_, _13651_, _13650_);
  and (_13653_, _13652_, _02393_);
  and (_13654_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and (_13655_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_13656_, _13655_, _13654_);
  and (_13657_, _13656_, _02445_);
  or (_13658_, _13657_, _13653_);
  and (_13659_, _13658_, _02421_);
  and (_13660_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and (_13661_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_13662_, _13661_, _13660_);
  and (_13663_, _13662_, _02393_);
  and (_13664_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and (_13665_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_13666_, _13665_, _13664_);
  and (_13667_, _13666_, _02445_);
  or (_13668_, _13667_, _13663_);
  and (_13669_, _13668_, _02459_);
  or (_13670_, _13669_, _02414_);
  or (_13671_, _13670_, _13659_);
  or (_13672_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_13673_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and (_13674_, _13673_, _13672_);
  and (_13675_, _13674_, _02393_);
  or (_13676_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_13677_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and (_13678_, _13677_, _13676_);
  and (_13679_, _13678_, _02445_);
  or (_13680_, _13679_, _13675_);
  and (_13681_, _13680_, _02421_);
  or (_13682_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_13683_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and (_13684_, _13683_, _13682_);
  and (_13685_, _13684_, _02393_);
  or (_13686_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_13687_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and (_13688_, _13687_, _13686_);
  and (_13689_, _13688_, _02445_);
  or (_13690_, _13689_, _13685_);
  and (_13691_, _13690_, _02459_);
  or (_13692_, _13691_, _02458_);
  or (_13693_, _13692_, _13681_);
  and (_13694_, _13693_, _13671_);
  or (_13695_, _13694_, _02496_);
  and (_13696_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  and (_13697_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or (_13698_, _13697_, _13696_);
  and (_13699_, _13698_, _02393_);
  and (_13700_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  and (_13701_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or (_13702_, _13701_, _13700_);
  and (_13703_, _13702_, _02445_);
  or (_13704_, _13703_, _13699_);
  and (_13705_, _13704_, _02421_);
  and (_13706_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  and (_13707_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or (_13708_, _13707_, _13706_);
  and (_13709_, _13708_, _02393_);
  and (_13710_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  and (_13711_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or (_13712_, _13711_, _13710_);
  and (_13713_, _13712_, _02445_);
  or (_13714_, _13713_, _13709_);
  and (_13715_, _13714_, _02459_);
  or (_13716_, _13715_, _02414_);
  or (_13717_, _13716_, _13705_);
  or (_13718_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or (_13719_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  and (_13720_, _13719_, _13718_);
  and (_13721_, _13720_, _02393_);
  or (_13722_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  or (_13723_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  and (_13724_, _13723_, _13722_);
  and (_13725_, _13724_, _02445_);
  or (_13726_, _13725_, _13721_);
  and (_13727_, _13726_, _02421_);
  or (_13728_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or (_13729_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  and (_13730_, _13729_, _13728_);
  and (_13731_, _13730_, _02393_);
  or (_13732_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or (_13733_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  and (_13734_, _13733_, _13732_);
  and (_13735_, _13734_, _02445_);
  or (_13736_, _13735_, _13731_);
  and (_13737_, _13736_, _02459_);
  or (_13738_, _13737_, _02458_);
  or (_13739_, _13738_, _13727_);
  and (_13740_, _13739_, _13717_);
  or (_13741_, _13740_, _02398_);
  and (_13742_, _13741_, _13695_);
  and (_13743_, _13742_, _02400_);
  or (_13744_, _13743_, _13649_);
  and (_13745_, _13744_, _02405_);
  or (_13746_, _13745_, _13555_);
  and (_13747_, _13746_, _02444_);
  or (_13748_, _13747_, _13365_);
  or (_13749_, _13748_, _02443_);
  or (_13750_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_13751_, _13750_, _22762_);
  and (_04033_, _13751_, _13749_);
  and (_13752_, _05336_, _24329_);
  not (_13753_, _13752_);
  and (_13754_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  and (_13755_, _13752_, _23946_);
  or (_04045_, _13755_, _13754_);
  and (_13756_, _06886_, _01808_);
  not (_13757_, _13756_);
  and (_13758_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_13759_, _13756_, _23946_);
  or (_04049_, _13759_, _13758_);
  nand (_13760_, _24352_, _22767_);
  or (_13761_, _22767_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_13762_, _13761_, _22762_);
  and (_26864_[3], _13762_, _13760_);
  and (_13763_, _24201_, _24005_);
  not (_13764_, _13763_);
  and (_13765_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and (_13766_, _13763_, _23707_);
  or (_04080_, _13766_, _13765_);
  and (_13767_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_13768_, _13756_, _23707_);
  or (_04090_, _13768_, _13767_);
  and (_13769_, _05336_, _25078_);
  not (_13770_, _13769_);
  and (_13771_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  and (_13772_, _13769_, _23747_);
  or (_27091_, _13772_, _13771_);
  and (_13773_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  and (_13774_, _13769_, _23898_);
  or (_04098_, _13774_, _13773_);
  and (_13775_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_13776_, _13756_, _24050_);
  or (_04111_, _13776_, _13775_);
  and (_13777_, _05336_, _24282_);
  not (_13778_, _13777_);
  and (_13779_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_13780_, _13777_, _23824_);
  or (_04114_, _13780_, _13779_);
  and (_13781_, _10347_, _23649_);
  and (_13782_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or (_04117_, _13782_, _13781_);
  and (_13783_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  and (_13784_, _13752_, _23824_);
  or (_04120_, _13784_, _13783_);
  and (_13785_, _05336_, _23752_);
  not (_13786_, _13785_);
  and (_13787_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_13788_, _13785_, _23707_);
  or (_04125_, _13788_, _13787_);
  and (_13789_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_13790_, _13785_, _23649_);
  or (_04133_, _13790_, _13789_);
  and (_13791_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and (_13792_, _12935_, _24050_);
  or (_04140_, _13792_, _13791_);
  or (_13793_, _24436_, _23837_);
  or (_13794_, _22767_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_13795_, _13794_, _22762_);
  and (_26864_[2], _13795_, _13793_);
  nand (_13796_, _24486_, _22767_);
  or (_13797_, _22767_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_13799_, _13797_, _22762_);
  and (_26864_[6], _13799_, _13796_);
  and (_13800_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  and (_13801_, _12941_, _23898_);
  or (_27100_, _13801_, _13800_);
  and (_13802_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  and (_13803_, _12970_, _24050_);
  or (_04171_, _13803_, _13802_);
  and (_13804_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  and (_13805_, _12970_, _23747_);
  or (_04174_, _13805_, _13804_);
  and (_13806_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_13807_, _12906_, _23778_);
  or (_04193_, _13807_, _13806_);
  and (_13808_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_13809_, _12974_, _23898_);
  or (_04195_, _13809_, _13808_);
  and (_13810_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and (_13811_, _12980_, _24050_);
  or (_04199_, _13811_, _13810_);
  and (_13812_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_13813_, _12980_, _23778_);
  or (_04203_, _13813_, _13812_);
  and (_13814_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_13815_, _13785_, _23778_);
  or (_04209_, _13815_, _13814_);
  and (_13816_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_13817_, _12906_, _23898_);
  or (_04212_, _13817_, _13816_);
  and (_13818_, _05336_, _23656_);
  not (_13819_, _13818_);
  and (_13820_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  and (_13821_, _13818_, _23747_);
  or (_04214_, _13821_, _13820_);
  and (_13822_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  and (_13823_, _13818_, _23778_);
  or (_04217_, _13823_, _13822_);
  and (_13824_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_13825_, _13777_, _23649_);
  or (_04225_, _13825_, _13824_);
  and (_13826_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_13827_, _12935_, _23778_);
  or (_04238_, _13827_, _13826_);
  and (_13828_, _06886_, _24329_);
  not (_13829_, _13828_);
  and (_13830_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  and (_13831_, _13828_, _23707_);
  or (_04246_, _13831_, _13830_);
  and (_13832_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_13833_, _12974_, _23946_);
  or (_04258_, _13833_, _13832_);
  and (_13834_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_13835_, _13756_, _23778_);
  or (_04270_, _13835_, _13834_);
  and (_13836_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  and (_13837_, _13769_, _23946_);
  or (_04275_, _13837_, _13836_);
  and (_13838_, _05125_, _23898_);
  and (_13839_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  or (_04330_, _13839_, _13838_);
  and (_13840_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_13841_, _13785_, _23747_);
  or (_04332_, _13841_, _13840_);
  and (_13842_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_13843_, _13785_, _23898_);
  or (_04345_, _13843_, _13842_);
  and (_13844_, _08043_, _23747_);
  and (_13845_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_27211_, _13845_, _13844_);
  and (_13846_, _05288_, _23824_);
  and (_13847_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or (_27056_, _13847_, _13846_);
  and (_13848_, _05288_, _23778_);
  and (_13849_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or (_04352_, _13849_, _13848_);
  and (_13850_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_13851_, _13756_, _23747_);
  or (_04355_, _13851_, _13850_);
  and (_13852_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and (_13853_, _13785_, _23824_);
  or (_04359_, _13853_, _13852_);
  and (_13854_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and (_13855_, _01967_, _23946_);
  or (_04364_, _13855_, _13854_);
  and (_13856_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_13857_, _13756_, _23824_);
  or (_04371_, _13857_, _13856_);
  and (_13858_, _12733_, _23707_);
  and (_13859_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  or (_04379_, _13859_, _13858_);
  and (_13860_, _05288_, _23747_);
  and (_13861_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or (_04382_, _13861_, _13860_);
  and (_13862_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_13863_, _13785_, _23946_);
  or (_04385_, _13863_, _13862_);
  and (_13864_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_13865_, _13756_, _23898_);
  or (_27012_, _13865_, _13864_);
  and (_13866_, _05125_, _23946_);
  and (_13867_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or (_27059_, _13867_, _13866_);
  and (_13868_, _05125_, _23747_);
  and (_13869_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  or (_04400_, _13869_, _13868_);
  and (_13870_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and (_13871_, _08351_, _23778_);
  or (_04409_, _13871_, _13870_);
  and (_13872_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and (_13873_, _13785_, _24050_);
  or (_04412_, _13873_, _13872_);
  and (_13874_, _12733_, _24050_);
  and (_13875_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  or (_04419_, _13875_, _13874_);
  and (_13876_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  and (_13877_, _13752_, _23778_);
  or (_04422_, _13877_, _13876_);
  and (_13878_, _05008_, _23747_);
  and (_13879_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_04446_, _13879_, _13878_);
  and (_13880_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  and (_13881_, _13828_, _23898_);
  or (_04450_, _13881_, _13880_);
  and (_13882_, _05008_, _23707_);
  and (_13883_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_27062_, _13883_, _13882_);
  and (_13884_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  and (_13885_, _13752_, _23898_);
  or (_04456_, _13885_, _13884_);
  and (_13886_, _05008_, _24050_);
  and (_13887_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_27061_, _13887_, _13886_);
  and (_13888_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  and (_13889_, _13828_, _23778_);
  or (_27010_, _13889_, _13888_);
  and (_13890_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_13891_, _13777_, _23898_);
  or (_04468_, _13891_, _13890_);
  and (_13892_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_13893_, _13777_, _23747_);
  or (_04472_, _13893_, _13892_);
  and (_13894_, _06886_, _23752_);
  not (_13895_, _13894_);
  and (_13896_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_13897_, _13894_, _23707_);
  or (_04482_, _13897_, _13896_);
  and (_13898_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and (_13899_, _13777_, _23946_);
  or (_04489_, _13899_, _13898_);
  and (_13900_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  and (_13901_, _02245_, _24050_);
  or (_04492_, _13901_, _13900_);
  and (_13902_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_13903_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or (_13904_, _13903_, _13902_);
  and (_13905_, _13904_, _02393_);
  and (_13906_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_13907_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_13908_, _13907_, _13906_);
  and (_13909_, _13908_, _02445_);
  or (_13910_, _13909_, _13905_);
  and (_13911_, _13910_, _02421_);
  and (_13912_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_13913_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_13914_, _13913_, _13912_);
  and (_13915_, _13914_, _02393_);
  and (_13916_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_13917_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or (_13918_, _13917_, _13916_);
  and (_13919_, _13918_, _02445_);
  or (_13920_, _13919_, _13915_);
  and (_13921_, _13920_, _02459_);
  or (_13922_, _13921_, _13911_);
  and (_13923_, _13922_, _02458_);
  or (_13924_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_13925_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_13926_, _13925_, _13924_);
  and (_13927_, _13926_, _02393_);
  or (_13928_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_13929_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and (_13930_, _13929_, _13928_);
  and (_13931_, _13930_, _02445_);
  or (_13932_, _13931_, _13927_);
  and (_13933_, _13932_, _02421_);
  or (_13934_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or (_13935_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_13936_, _13935_, _13934_);
  and (_13937_, _13936_, _02393_);
  or (_13938_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or (_13939_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_13940_, _13939_, _13938_);
  and (_13941_, _13940_, _02445_);
  or (_13942_, _13941_, _13937_);
  and (_13943_, _13942_, _02459_);
  or (_13944_, _13943_, _13933_);
  and (_13945_, _13944_, _02414_);
  or (_13946_, _13945_, _13923_);
  and (_13947_, _13946_, _02398_);
  and (_13948_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and (_13949_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or (_13950_, _13949_, _13948_);
  and (_13951_, _13950_, _02393_);
  and (_13952_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and (_13953_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_13954_, _13953_, _13952_);
  and (_13955_, _13954_, _02445_);
  or (_13956_, _13955_, _13951_);
  and (_13957_, _13956_, _02421_);
  and (_13958_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and (_13959_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or (_13960_, _13959_, _13958_);
  and (_13961_, _13960_, _02393_);
  and (_13962_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and (_13963_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_13964_, _13963_, _13962_);
  and (_13965_, _13964_, _02445_);
  or (_13966_, _13965_, _13961_);
  and (_13967_, _13966_, _02459_);
  or (_13968_, _13967_, _13957_);
  and (_13969_, _13968_, _02458_);
  or (_13970_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or (_13971_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and (_13972_, _13971_, _02445_);
  and (_13973_, _13972_, _13970_);
  or (_13974_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_13975_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and (_13976_, _13975_, _02393_);
  and (_13977_, _13976_, _13974_);
  or (_13978_, _13977_, _13973_);
  and (_13979_, _13978_, _02421_);
  or (_13980_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or (_13981_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and (_13982_, _13981_, _02445_);
  and (_13983_, _13982_, _13980_);
  or (_13984_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_13985_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and (_13986_, _13985_, _02393_);
  and (_13987_, _13986_, _13984_);
  or (_13988_, _13987_, _13983_);
  and (_13989_, _13988_, _02459_);
  or (_13990_, _13989_, _13979_);
  and (_13991_, _13990_, _02414_);
  or (_13992_, _13991_, _13969_);
  and (_13993_, _13992_, _02496_);
  or (_13994_, _13993_, _13947_);
  and (_13995_, _13994_, _02400_);
  and (_13996_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_13997_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or (_13998_, _13997_, _13996_);
  and (_13999_, _13998_, _02393_);
  and (_14000_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_14001_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or (_14002_, _14001_, _14000_);
  and (_14003_, _14002_, _02445_);
  or (_14004_, _14003_, _13999_);
  or (_14005_, _14004_, _02459_);
  and (_14006_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_14007_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or (_14008_, _14007_, _14006_);
  and (_14009_, _14008_, _02393_);
  and (_14010_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_14011_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or (_14012_, _14011_, _14010_);
  and (_14013_, _14012_, _02445_);
  or (_14014_, _14013_, _14009_);
  or (_14015_, _14014_, _02421_);
  and (_14016_, _14015_, _02458_);
  and (_14017_, _14016_, _14005_);
  or (_14018_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or (_14019_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_14020_, _14019_, _02445_);
  and (_14021_, _14020_, _14018_);
  or (_14022_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or (_14023_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_14024_, _14023_, _02393_);
  and (_14025_, _14024_, _14022_);
  or (_14026_, _14025_, _14021_);
  or (_14027_, _14026_, _02459_);
  or (_14028_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or (_14029_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_14030_, _14029_, _02445_);
  and (_14031_, _14030_, _14028_);
  or (_14032_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or (_14033_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_14034_, _14033_, _02393_);
  and (_14035_, _14034_, _14032_);
  or (_14036_, _14035_, _14031_);
  or (_14037_, _14036_, _02421_);
  and (_14038_, _14037_, _02414_);
  and (_14039_, _14038_, _14027_);
  or (_14040_, _14039_, _14017_);
  and (_14041_, _14040_, _02496_);
  and (_14042_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and (_14043_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_14044_, _14043_, _14042_);
  and (_14045_, _14044_, _02393_);
  and (_14046_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and (_14047_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_14048_, _14047_, _14046_);
  and (_14049_, _14048_, _02445_);
  or (_14050_, _14049_, _14045_);
  or (_14051_, _14050_, _02459_);
  and (_14052_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and (_14053_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_14054_, _14053_, _14052_);
  and (_14055_, _14054_, _02393_);
  and (_14056_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and (_14057_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_14058_, _14057_, _14056_);
  and (_14059_, _14058_, _02445_);
  or (_14060_, _14059_, _14055_);
  or (_14061_, _14060_, _02421_);
  and (_14062_, _14061_, _02458_);
  and (_14063_, _14062_, _14051_);
  or (_14064_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_14065_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and (_14066_, _14065_, _14064_);
  and (_14067_, _14066_, _02393_);
  or (_14068_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_14069_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and (_14070_, _14069_, _14068_);
  and (_14071_, _14070_, _02445_);
  or (_14072_, _14071_, _14067_);
  or (_14073_, _14072_, _02459_);
  or (_14074_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_14075_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and (_14076_, _14075_, _14074_);
  and (_14077_, _14076_, _02393_);
  or (_14078_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_14079_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and (_14080_, _14079_, _14078_);
  and (_14081_, _14080_, _02445_);
  or (_14082_, _14081_, _14077_);
  or (_14083_, _14082_, _02421_);
  and (_14084_, _14083_, _02414_);
  and (_14085_, _14084_, _14073_);
  or (_14086_, _14085_, _14063_);
  and (_14087_, _14086_, _02398_);
  or (_14088_, _14087_, _14041_);
  and (_14089_, _14088_, _02546_);
  or (_14090_, _14089_, _13995_);
  and (_14091_, _14090_, _02646_);
  or (_14092_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_14093_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and (_14094_, _14093_, _02445_);
  and (_14095_, _14094_, _14092_);
  or (_14096_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_14097_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and (_14098_, _14097_, _02393_);
  and (_14099_, _14098_, _14096_);
  or (_14100_, _14099_, _14095_);
  and (_14101_, _14100_, _02459_);
  or (_14102_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_14103_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and (_14104_, _14103_, _02445_);
  and (_14105_, _14104_, _14102_);
  or (_14106_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_14107_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and (_14108_, _14107_, _02393_);
  and (_14109_, _14108_, _14106_);
  or (_14110_, _14109_, _14105_);
  and (_14111_, _14110_, _02421_);
  or (_14112_, _14111_, _14101_);
  and (_14113_, _14112_, _02414_);
  and (_14114_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and (_14115_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_14116_, _14115_, _14114_);
  and (_14117_, _14116_, _02393_);
  and (_14118_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and (_14119_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_14120_, _14119_, _14118_);
  and (_14121_, _14120_, _02445_);
  or (_14122_, _14121_, _14117_);
  and (_14123_, _14122_, _02459_);
  and (_14124_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and (_14125_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_14126_, _14125_, _14124_);
  and (_14127_, _14126_, _02393_);
  and (_14128_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and (_14129_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_14130_, _14129_, _14128_);
  and (_14131_, _14130_, _02445_);
  or (_14132_, _14131_, _14127_);
  and (_14133_, _14132_, _02421_);
  or (_14134_, _14133_, _14123_);
  and (_14135_, _14134_, _02458_);
  or (_14136_, _14135_, _14113_);
  and (_14137_, _14136_, _02496_);
  or (_14138_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or (_14139_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and (_14140_, _14139_, _14138_);
  and (_14141_, _14140_, _02393_);
  or (_14142_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_14143_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_14144_, _14143_, _14142_);
  and (_14145_, _14144_, _02445_);
  or (_14146_, _14145_, _14141_);
  and (_14147_, _14146_, _02459_);
  or (_14148_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or (_14149_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and (_14150_, _14149_, _14148_);
  and (_14151_, _14150_, _02393_);
  or (_14152_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_14153_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_14154_, _14153_, _14152_);
  and (_14155_, _14154_, _02445_);
  or (_14156_, _14155_, _14151_);
  and (_14157_, _14156_, _02421_);
  or (_14158_, _14157_, _14147_);
  and (_14159_, _14158_, _02414_);
  and (_14160_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_14161_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_14162_, _14161_, _14160_);
  and (_14163_, _14162_, _02393_);
  and (_14164_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_14165_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or (_14166_, _14165_, _14164_);
  and (_14167_, _14166_, _02445_);
  or (_14168_, _14167_, _14163_);
  and (_14169_, _14168_, _02459_);
  and (_14170_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_14171_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or (_14172_, _14171_, _14170_);
  and (_14173_, _14172_, _02393_);
  and (_14174_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_14175_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_14176_, _14175_, _14174_);
  and (_14177_, _14176_, _02445_);
  or (_14178_, _14177_, _14173_);
  and (_14179_, _14178_, _02421_);
  or (_14180_, _14179_, _14169_);
  and (_14181_, _14180_, _02458_);
  or (_14182_, _14181_, _14159_);
  and (_14183_, _14182_, _02398_);
  or (_14184_, _14183_, _14137_);
  and (_14185_, _14184_, _02400_);
  and (_14186_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and (_14187_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_14188_, _14187_, _14186_);
  and (_14189_, _14188_, _02393_);
  and (_14190_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and (_14191_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_14192_, _14191_, _14190_);
  and (_14193_, _14192_, _02445_);
  or (_14194_, _14193_, _14189_);
  or (_14195_, _14194_, _02459_);
  and (_14196_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and (_14197_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_14198_, _14197_, _14196_);
  and (_14199_, _14198_, _02393_);
  and (_14200_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and (_14201_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_14202_, _14201_, _14200_);
  and (_14203_, _14202_, _02445_);
  or (_14204_, _14203_, _14199_);
  or (_14205_, _14204_, _02421_);
  and (_14206_, _14205_, _02458_);
  and (_14207_, _14206_, _14195_);
  or (_14208_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_14209_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and (_14210_, _14209_, _14208_);
  and (_14211_, _14210_, _02393_);
  or (_14212_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_14213_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and (_14214_, _14213_, _14212_);
  and (_14215_, _14214_, _02445_);
  or (_14216_, _14215_, _14211_);
  or (_14217_, _14216_, _02459_);
  or (_14218_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_14219_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and (_14220_, _14219_, _14218_);
  and (_14221_, _14220_, _02393_);
  or (_14222_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_14223_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and (_14224_, _14223_, _14222_);
  and (_14225_, _14224_, _02445_);
  or (_14226_, _14225_, _14221_);
  or (_14227_, _14226_, _02421_);
  and (_14228_, _14227_, _02414_);
  and (_14229_, _14228_, _14217_);
  or (_14230_, _14229_, _14207_);
  and (_14231_, _14230_, _02398_);
  and (_14232_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and (_14233_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_14234_, _14233_, _14232_);
  and (_14235_, _14234_, _02393_);
  and (_14236_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and (_14237_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_14238_, _14237_, _14236_);
  and (_14239_, _14238_, _02445_);
  or (_14240_, _14239_, _14235_);
  or (_14241_, _14240_, _02459_);
  and (_14242_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and (_14243_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_14244_, _14243_, _14242_);
  and (_14245_, _14244_, _02393_);
  and (_14246_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and (_14247_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_14248_, _14247_, _14246_);
  and (_14249_, _14248_, _02445_);
  or (_14250_, _14249_, _14245_);
  or (_14251_, _14250_, _02421_);
  and (_14252_, _14251_, _02458_);
  and (_14253_, _14252_, _14241_);
  or (_14254_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_14255_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and (_14256_, _14255_, _02445_);
  and (_14257_, _14256_, _14254_);
  or (_14258_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_14259_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and (_14260_, _14259_, _02393_);
  and (_14261_, _14260_, _14258_);
  or (_14262_, _14261_, _14257_);
  or (_14263_, _14262_, _02459_);
  or (_14264_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_14265_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and (_14266_, _14265_, _02445_);
  and (_14267_, _14266_, _14264_);
  or (_14268_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_14269_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and (_14270_, _14269_, _02393_);
  and (_14271_, _14270_, _14268_);
  or (_14272_, _14271_, _14267_);
  or (_14273_, _14272_, _02421_);
  and (_14274_, _14273_, _02414_);
  and (_14275_, _14274_, _14263_);
  or (_14276_, _14275_, _14253_);
  and (_14277_, _14276_, _02496_);
  or (_14278_, _14277_, _14231_);
  and (_14279_, _14278_, _02546_);
  or (_14280_, _14279_, _14185_);
  and (_14281_, _14280_, _02405_);
  or (_14282_, _14281_, _14091_);
  and (_14283_, _14282_, _26777_);
  and (_14284_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and (_14285_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_14286_, _14285_, _14284_);
  and (_14287_, _14286_, _02393_);
  and (_14288_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and (_14289_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_14290_, _14289_, _14288_);
  and (_14291_, _14290_, _02445_);
  or (_14292_, _14291_, _14287_);
  and (_14293_, _14292_, _02421_);
  and (_14294_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and (_14295_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_14296_, _14295_, _14294_);
  and (_14297_, _14296_, _02393_);
  and (_14298_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and (_14299_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_14300_, _14299_, _14298_);
  and (_14301_, _14300_, _02445_);
  or (_14302_, _14301_, _14297_);
  and (_14303_, _14302_, _02459_);
  or (_14304_, _14303_, _02414_);
  or (_14305_, _14304_, _14293_);
  or (_14306_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_14307_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and (_14308_, _14307_, _14306_);
  and (_14309_, _14308_, _02393_);
  or (_14310_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_14311_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and (_14312_, _14311_, _14310_);
  and (_14313_, _14312_, _02445_);
  or (_14314_, _14313_, _14309_);
  and (_14315_, _14314_, _02421_);
  or (_14316_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_14317_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and (_14318_, _14317_, _14316_);
  and (_14319_, _14318_, _02393_);
  or (_14320_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_14321_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and (_14322_, _14321_, _14320_);
  and (_14323_, _14322_, _02445_);
  or (_14324_, _14323_, _14319_);
  and (_14325_, _14324_, _02459_);
  or (_14326_, _14325_, _02458_);
  or (_14327_, _14326_, _14315_);
  and (_14328_, _14327_, _14305_);
  or (_14329_, _14328_, _02496_);
  and (_14330_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_14331_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_14332_, _14331_, _14330_);
  and (_14333_, _14332_, _02393_);
  and (_14334_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_14335_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_14336_, _14335_, _14334_);
  and (_14337_, _14336_, _02445_);
  or (_14338_, _14337_, _14333_);
  and (_14339_, _14338_, _02421_);
  and (_14340_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_14341_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_14342_, _14341_, _14340_);
  and (_14343_, _14342_, _02393_);
  and (_14344_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_14345_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_14346_, _14345_, _14344_);
  and (_14347_, _14346_, _02445_);
  or (_14348_, _14347_, _14343_);
  and (_14349_, _14348_, _02459_);
  or (_14350_, _14349_, _02414_);
  or (_14351_, _14350_, _14339_);
  or (_14352_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_14353_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_14354_, _14353_, _02445_);
  and (_14355_, _14354_, _14352_);
  or (_14356_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_14357_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_14358_, _14357_, _02393_);
  and (_14359_, _14358_, _14356_);
  or (_14360_, _14359_, _14355_);
  and (_14361_, _14360_, _02421_);
  or (_14362_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_14363_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_14364_, _14363_, _02445_);
  and (_14365_, _14364_, _14362_);
  or (_14366_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_14367_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_14368_, _14367_, _02393_);
  and (_14369_, _14368_, _14366_);
  or (_14370_, _14369_, _14365_);
  and (_14371_, _14370_, _02459_);
  or (_14372_, _14371_, _02458_);
  or (_14373_, _14372_, _14361_);
  and (_14374_, _14373_, _14351_);
  or (_14375_, _14374_, _02398_);
  and (_14376_, _14375_, _14329_);
  and (_14377_, _14376_, _02400_);
  and (_14378_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and (_14379_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_14380_, _14379_, _14378_);
  and (_14381_, _14380_, _02393_);
  and (_14382_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and (_14383_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_14384_, _14383_, _14382_);
  and (_14385_, _14384_, _02445_);
  or (_14386_, _14385_, _14381_);
  or (_14387_, _14386_, _02459_);
  and (_14388_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and (_14389_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_14390_, _14389_, _14388_);
  and (_14391_, _14390_, _02393_);
  and (_14392_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and (_14393_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_14394_, _14393_, _14392_);
  and (_14395_, _14394_, _02445_);
  or (_14396_, _14395_, _14391_);
  or (_14397_, _14396_, _02421_);
  and (_14398_, _14397_, _02458_);
  and (_14399_, _14398_, _14387_);
  or (_14400_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_14401_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and (_14402_, _14401_, _02445_);
  and (_14403_, _14402_, _14400_);
  or (_14404_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_14405_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and (_14406_, _14405_, _02393_);
  and (_14407_, _14406_, _14404_);
  or (_14408_, _14407_, _14403_);
  or (_14409_, _14408_, _02459_);
  or (_14410_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_14411_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and (_14412_, _14411_, _02445_);
  and (_14413_, _14412_, _14410_);
  or (_14414_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_14415_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and (_14416_, _14415_, _02393_);
  and (_14417_, _14416_, _14414_);
  or (_14418_, _14417_, _14413_);
  or (_14419_, _14418_, _02421_);
  and (_14420_, _14419_, _02414_);
  and (_14421_, _14420_, _14409_);
  or (_14422_, _14421_, _14399_);
  or (_14423_, _14422_, _02398_);
  and (_14424_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_14425_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_14426_, _14425_, _14424_);
  and (_14427_, _14426_, _02393_);
  and (_14428_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and (_14429_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_14430_, _14429_, _14428_);
  and (_14431_, _14430_, _02445_);
  or (_14432_, _14431_, _14427_);
  or (_14433_, _14432_, _02459_);
  and (_14434_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and (_14435_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_14436_, _14435_, _14434_);
  and (_14437_, _14436_, _02393_);
  and (_14438_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and (_14439_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_14440_, _14439_, _14438_);
  and (_14441_, _14440_, _02445_);
  or (_14442_, _14441_, _14437_);
  or (_14443_, _14442_, _02421_);
  and (_14444_, _14443_, _02458_);
  and (_14445_, _14444_, _14433_);
  or (_14446_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_14447_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and (_14448_, _14447_, _14446_);
  and (_14449_, _14448_, _02393_);
  or (_14451_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_14452_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and (_14453_, _14452_, _14451_);
  and (_14454_, _14453_, _02445_);
  or (_14455_, _14454_, _14449_);
  or (_14456_, _14455_, _02459_);
  or (_14457_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_14458_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and (_14459_, _14458_, _14457_);
  and (_14460_, _14459_, _02393_);
  or (_14461_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_14462_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and (_14463_, _14462_, _14461_);
  and (_14464_, _14463_, _02445_);
  or (_14465_, _14464_, _14460_);
  or (_14466_, _14465_, _02421_);
  and (_14467_, _14466_, _02414_);
  and (_14468_, _14467_, _14456_);
  or (_14469_, _14468_, _14445_);
  or (_14470_, _14469_, _02496_);
  and (_14471_, _14470_, _14423_);
  and (_14472_, _14471_, _02546_);
  or (_14473_, _14472_, _14377_);
  and (_14474_, _14473_, _02646_);
  and (_14475_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and (_14476_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_14477_, _14476_, _14475_);
  and (_14478_, _14477_, _02445_);
  and (_14479_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and (_14480_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_14481_, _14480_, _14479_);
  and (_14482_, _14481_, _02393_);
  or (_14483_, _14482_, _14478_);
  or (_14484_, _14483_, _02459_);
  and (_14485_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and (_14486_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_14487_, _14486_, _14485_);
  and (_14488_, _14487_, _02445_);
  and (_14489_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and (_14490_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_14491_, _14490_, _14489_);
  and (_14492_, _14491_, _02393_);
  or (_14493_, _14492_, _14488_);
  or (_14494_, _14493_, _02421_);
  and (_14495_, _14494_, _02458_);
  and (_14496_, _14495_, _14484_);
  or (_14497_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_14498_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and (_14499_, _14498_, _02393_);
  and (_14500_, _14499_, _14497_);
  or (_14501_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_14502_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and (_14503_, _14502_, _02445_);
  and (_14504_, _14503_, _14501_);
  or (_14505_, _14504_, _14500_);
  or (_14506_, _14505_, _02459_);
  or (_14507_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_14508_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and (_14509_, _14508_, _02393_);
  and (_14510_, _14509_, _14507_);
  or (_14511_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_14512_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and (_14513_, _14512_, _02445_);
  and (_14514_, _14513_, _14511_);
  or (_14515_, _14514_, _14510_);
  or (_14516_, _14515_, _02421_);
  and (_14517_, _14516_, _02414_);
  and (_14518_, _14517_, _14506_);
  or (_14519_, _14518_, _14496_);
  or (_14520_, _14519_, _02398_);
  and (_14521_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and (_14522_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_14523_, _14522_, _02393_);
  or (_14524_, _14523_, _14521_);
  and (_14525_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and (_14526_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_14527_, _14526_, _02445_);
  or (_14528_, _14527_, _14525_);
  and (_14529_, _14528_, _14524_);
  or (_14530_, _14529_, _02459_);
  and (_14531_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and (_14532_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_14533_, _14532_, _02393_);
  or (_14534_, _14533_, _14531_);
  and (_14535_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and (_14536_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_14537_, _14536_, _02445_);
  or (_14538_, _14537_, _14535_);
  and (_14539_, _14538_, _14534_);
  or (_14540_, _14539_, _02421_);
  and (_14541_, _14540_, _02458_);
  and (_14542_, _14541_, _14530_);
  or (_14543_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_14544_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and (_14545_, _14544_, _14543_);
  or (_14546_, _14545_, _02445_);
  or (_14547_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_14548_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and (_14549_, _14548_, _14547_);
  or (_14550_, _14549_, _02393_);
  and (_14551_, _14550_, _14546_);
  or (_14552_, _14551_, _02459_);
  or (_14553_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_14554_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and (_14555_, _14554_, _14553_);
  or (_14556_, _14555_, _02445_);
  or (_14557_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_14558_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and (_14559_, _14558_, _14557_);
  or (_14560_, _14559_, _02393_);
  and (_14561_, _14560_, _14556_);
  or (_14562_, _14561_, _02421_);
  and (_14563_, _14562_, _02414_);
  and (_14564_, _14563_, _14552_);
  or (_14565_, _14564_, _14542_);
  or (_14566_, _14565_, _02496_);
  and (_14567_, _14566_, _02546_);
  and (_14568_, _14567_, _14520_);
  and (_14569_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and (_14570_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_14571_, _14570_, _14569_);
  and (_14572_, _14571_, _02393_);
  and (_14573_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and (_14574_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_14575_, _14574_, _14573_);
  and (_14576_, _14575_, _02445_);
  or (_14577_, _14576_, _14572_);
  and (_14578_, _14577_, _02421_);
  and (_14579_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and (_14580_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_14581_, _14580_, _14579_);
  and (_14582_, _14581_, _02393_);
  and (_14583_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and (_14584_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_14585_, _14584_, _14583_);
  and (_14586_, _14585_, _02445_);
  or (_14587_, _14586_, _14582_);
  and (_14588_, _14587_, _02459_);
  or (_14589_, _14588_, _02414_);
  or (_14590_, _14589_, _14578_);
  or (_14591_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_14592_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and (_14593_, _14592_, _14591_);
  and (_14594_, _14593_, _02393_);
  or (_14595_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_14596_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and (_14597_, _14596_, _14595_);
  and (_14598_, _14597_, _02445_);
  or (_14599_, _14598_, _14594_);
  and (_14600_, _14599_, _02421_);
  or (_14602_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_14603_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and (_14604_, _14603_, _14602_);
  and (_14605_, _14604_, _02393_);
  or (_14606_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_14607_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and (_14608_, _14607_, _14606_);
  and (_14609_, _14608_, _02445_);
  or (_14610_, _14609_, _14605_);
  and (_14611_, _14610_, _02459_);
  or (_14612_, _14611_, _02458_);
  or (_14613_, _14612_, _14600_);
  and (_14614_, _14613_, _14590_);
  or (_14615_, _14614_, _02496_);
  and (_14616_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  and (_14617_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or (_14618_, _14617_, _14616_);
  and (_14619_, _14618_, _02393_);
  and (_14620_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  and (_14621_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or (_14622_, _14621_, _14620_);
  and (_14623_, _14622_, _02445_);
  or (_14624_, _14623_, _14619_);
  and (_14625_, _14624_, _02421_);
  and (_14626_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  and (_14627_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or (_14628_, _14627_, _14626_);
  and (_14629_, _14628_, _02393_);
  and (_14630_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  and (_14631_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or (_14632_, _14631_, _14630_);
  and (_14633_, _14632_, _02445_);
  or (_14634_, _14633_, _14629_);
  and (_14635_, _14634_, _02459_);
  or (_14636_, _14635_, _02414_);
  or (_14637_, _14636_, _14625_);
  or (_14638_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or (_14639_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  and (_14640_, _14639_, _14638_);
  and (_14641_, _14640_, _02393_);
  or (_14642_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or (_14643_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  and (_14644_, _14643_, _14642_);
  and (_14645_, _14644_, _02445_);
  or (_14646_, _14645_, _14641_);
  and (_14647_, _14646_, _02421_);
  or (_14648_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or (_14649_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  and (_14650_, _14649_, _14648_);
  and (_14651_, _14650_, _02393_);
  or (_14652_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or (_14653_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  and (_14654_, _14653_, _14652_);
  and (_14655_, _14654_, _02445_);
  or (_14656_, _14655_, _14651_);
  and (_14657_, _14656_, _02459_);
  or (_14658_, _14657_, _02458_);
  or (_14659_, _14658_, _14647_);
  and (_14660_, _14659_, _14637_);
  or (_14661_, _14660_, _02398_);
  and (_14662_, _14661_, _14615_);
  and (_14663_, _14662_, _02400_);
  or (_14664_, _14663_, _14568_);
  and (_14665_, _14664_, _02405_);
  or (_14666_, _14665_, _14474_);
  and (_14667_, _14666_, _02444_);
  or (_14668_, _14667_, _14283_);
  or (_14669_, _14668_, _02443_);
  or (_14670_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_14671_, _14670_, _22762_);
  and (_04499_, _14671_, _14669_);
  and (_14672_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_14673_, _13777_, _24050_);
  or (_04502_, _14673_, _14672_);
  and (_14674_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_14675_, _02204_, _23898_);
  or (_04503_, _14675_, _14674_);
  and (_14676_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and (_14677_, _13763_, _24050_);
  or (_27245_, _14677_, _14676_);
  and (_14678_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_14679_, _02204_, _23707_);
  or (_04512_, _14679_, _14678_);
  and (_14680_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and (_14681_, _13777_, _23707_);
  or (_27090_, _14681_, _14680_);
  and (_14682_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_14683_, _25763_, _23747_);
  or (_04530_, _14683_, _14682_);
  and (_14684_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  and (_14685_, _13769_, _23778_);
  or (_04534_, _14685_, _14684_);
  and (_14686_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  and (_14687_, _13828_, _23649_);
  or (_04539_, _14687_, _14686_);
  and (_14688_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_14689_, _25763_, _23707_);
  or (_04542_, _14689_, _14688_);
  nor (_14690_, t2ex_i, rst);
  and (_04546_, _14690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  and (_14691_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  and (_14692_, _13769_, _23824_);
  or (_04548_, _14692_, _14691_);
  and (_14693_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_14694_, _25763_, _24050_);
  or (_04550_, _14694_, _14693_);
  and (_14695_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  and (_14696_, _13769_, _23649_);
  or (_04553_, _14696_, _14695_);
  and (_14697_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  and (_14698_, _13828_, _23747_);
  or (_27011_, _14698_, _14697_);
  and (_14699_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  and (_14700_, _25542_, _23898_);
  or (_04562_, _14700_, _14699_);
  and (_14701_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  and (_14702_, _13769_, _24050_);
  or (_27092_, _14702_, _14701_);
  and (_14703_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  and (_14704_, _13828_, _23824_);
  or (_04566_, _14704_, _14703_);
  and (_14705_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  and (_14706_, _25252_, _23649_);
  or (_27044_, _14706_, _14705_);
  and (_14707_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  and (_14708_, _13769_, _23707_);
  or (_04573_, _14708_, _14707_);
  and (_14709_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_14710_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_14711_, _22770_, _14710_);
  or (_14712_, _14711_, _14709_);
  and (_26882_[15], _14712_, _22762_);
  and (_14713_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  and (_14714_, _25252_, _23824_);
  or (_04577_, _14714_, _14713_);
  and (_14715_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  and (_14716_, _13818_, _23898_);
  or (_04580_, _14716_, _14715_);
  and (_14717_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_14718_, _24767_, _23778_);
  or (_04583_, _14718_, _14717_);
  not (_14719_, _24174_);
  and (_14720_, _14719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_14721_, _24145_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_14722_, _14721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_14723_, _14722_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_14724_, _14723_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_14725_, _24173_, _24178_);
  and (_14726_, _14725_, _14724_);
  and (_14727_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_14728_, _14727_, _14726_);
  nor (_14729_, _14728_, _24127_);
  or (_14730_, _14729_, _14720_);
  and (_14731_, _14730_, _24166_);
  and (_14732_, _24121_, _23738_);
  or (_04585_, _14732_, _14731_);
  and (_14733_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and (_14734_, _25252_, _23707_);
  or (_04587_, _14734_, _14733_);
  and (_14735_, _24121_, _24685_);
  nor (_14736_, _24145_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_14737_, _14736_, _14721_);
  and (_14738_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_14739_, _14738_, _14737_);
  nand (_14740_, _14739_, _24174_);
  or (_14741_, _24174_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_14742_, _14741_, _14740_);
  and (_14743_, _14742_, _24166_);
  or (_04590_, _14743_, _14735_);
  and (_14744_, _08799_, _24050_);
  and (_14745_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or (_04592_, _14745_, _14744_);
  and (_14746_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_14747_, _24767_, _23707_);
  or (_04597_, _14747_, _14746_);
  and (_14748_, _24852_, _23778_);
  and (_14749_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or (_04610_, _14749_, _14748_);
  nor (_26897_[1], _00392_, rst);
  and (_14750_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  and (_14751_, _13818_, _23824_);
  or (_04614_, _14751_, _14750_);
  and (_14752_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_14753_, _24767_, _23649_);
  or (_04617_, _14753_, _14752_);
  and (_14754_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  and (_14755_, _13818_, _23649_);
  or (_04620_, _14755_, _14754_);
  or (_14756_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_14757_, _14756_, _22762_);
  or (_14758_, _02037_, _23642_);
  and (_04622_, _14758_, _14757_);
  and (_14759_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_14760_, _24127_, _23772_);
  nor (_14761_, _24159_, _24155_);
  and (_14762_, _14761_, _24157_);
  nor (_14763_, _14761_, _24157_);
  or (_14764_, _14763_, _14762_);
  or (_14765_, _14764_, _24127_);
  and (_14766_, _14765_, _14760_);
  and (_14767_, _14766_, _24166_);
  or (_04624_, _14767_, _14759_);
  and (_14768_, _24226_, _23824_);
  and (_14769_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  or (_04626_, _14769_, _14768_);
  and (_14770_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  and (_14771_, _13818_, _23946_);
  or (_27093_, _14771_, _14770_);
  and (_14772_, _24194_, _23824_);
  and (_14773_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_27047_, _14773_, _14772_);
  and (_14774_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  and (_14775_, _13818_, _24050_);
  or (_27094_, _14775_, _14774_);
  and (_14776_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_14777_, _13894_, _23824_);
  or (_04635_, _14777_, _14776_);
  and (_14778_, _02313_, _23824_);
  and (_14779_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_04638_, _14779_, _14778_);
  and (_14780_, _08043_, _23649_);
  and (_14781_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_04640_, _14781_, _14780_);
  and (_14782_, _26113_, _26110_);
  nor (_14783_, _09920_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_14784_, _14783_, _14782_);
  and (_14785_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_14786_, _14785_, _04864_);
  nor (_14787_, _14786_, _14784_);
  nor (_14788_, _14787_, _24299_);
  and (_14789_, _24299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_14790_, _14789_, _14788_);
  and (_14791_, _14790_, _24294_);
  and (_14792_, _24293_, _23738_);
  or (_14793_, _14792_, _14791_);
  and (_04642_, _14793_, _22762_);
  and (_14794_, _24194_, _23946_);
  and (_14795_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_04645_, _14795_, _14794_);
  and (_14796_, _02313_, _23898_);
  and (_14797_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_04647_, _14797_, _14796_);
  and (_14798_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and (_14799_, _13894_, _23898_);
  or (_04649_, _14799_, _14798_);
  and (_14800_, _24081_, _24050_);
  and (_14801_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_04651_, _14801_, _14800_);
  and (_14802_, _02313_, _23778_);
  and (_14803_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_04653_, _14803_, _14802_);
  and (_14804_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  and (_14805_, _13818_, _23707_);
  or (_04655_, _14805_, _14804_);
  or (_14806_, _04891_, _23816_);
  or (_14807_, _04880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_14808_, _14807_, _26097_);
  nor (_14809_, _14808_, _04881_);
  and (_14810_, _04864_, _24307_);
  or (_14811_, _14810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  not (_14812_, _04866_);
  and (_14813_, _14812_, _04860_);
  and (_14814_, _14813_, _14811_);
  and (_14815_, _24307_, _24300_);
  and (_14816_, _14815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_14817_, _14816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_14818_, _04874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_14819_, _14818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_14820_, _14819_, _14817_);
  or (_14821_, _14820_, _14814_);
  or (_14822_, _14821_, _14809_);
  or (_14823_, _14822_, _24299_);
  and (_14824_, _14823_, _24294_);
  and (_14825_, _14824_, _14806_);
  and (_14826_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_14827_, _14826_, _14825_);
  and (_04657_, _14827_, _22762_);
  or (_14828_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_14829_, _14828_, _22762_);
  or (_14830_, _24079_, _23816_);
  and (_04659_, _14830_, _14829_);
  and (_14831_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and (_14832_, _13894_, _23778_);
  or (_04662_, _14832_, _14831_);
  and (_14833_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  and (_14834_, _13752_, _23747_);
  or (_04664_, _14834_, _14833_);
  and (_14835_, _23898_, _23755_);
  and (_14836_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or (_04670_, _14836_, _14835_);
  and (_14837_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  and (_14838_, _13752_, _23649_);
  or (_04672_, _14838_, _14837_);
  and (_14839_, _08799_, _23946_);
  and (_14840_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or (_04687_, _14840_, _14839_);
  and (_14841_, _23833_, _23707_);
  and (_14842_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_04689_, _14842_, _14841_);
  and (_14843_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  and (_14844_, _13752_, _24050_);
  or (_04692_, _14844_, _14843_);
  and (_14845_, _02313_, _23707_);
  and (_14846_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_04697_, _14846_, _14845_);
  and (_14847_, _02200_, _23747_);
  and (_14848_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_04699_, _14848_, _14847_);
  and (_14849_, _02200_, _23946_);
  and (_14850_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_27167_, _14850_, _14849_);
  and (_14851_, _24331_, _23747_);
  and (_14852_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_04710_, _14852_, _14851_);
  and (_14853_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  and (_14854_, _13752_, _23707_);
  or (_04713_, _14854_, _14853_);
  or (_14855_, _24464_, _23837_);
  or (_14856_, _22767_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_14857_, _14856_, _22762_);
  and (_26864_[4], _14857_, _14855_);
  and (_14858_, _02313_, _23946_);
  and (_14859_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_04716_, _14859_, _14858_);
  and (_14860_, _24331_, _23898_);
  and (_14861_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_04719_, _14861_, _14860_);
  and (_14862_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_14863_, _12980_, _23898_);
  or (_04722_, _14863_, _14862_);
  and (_14864_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_14865_, _12980_, _23824_);
  or (_04731_, _14865_, _14864_);
  and (_14866_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_04733_, _14866_, _05664_);
  and (_14867_, _05350_, _23946_);
  and (_14868_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or (_27065_, _14868_, _14867_);
  and (_14869_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_14870_, _13894_, _23946_);
  or (_04739_, _14870_, _14869_);
  and (_14871_, _02313_, _23747_);
  and (_14872_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_27156_, _14872_, _14871_);
  and (_14873_, _04811_, _24050_);
  and (_14874_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  or (_04747_, _14874_, _14873_);
  and (_14875_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and (_14876_, _12980_, _23747_);
  or (_04750_, _14876_, _14875_);
  and (_14877_, _04811_, _23649_);
  and (_14878_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or (_04753_, _14878_, _14877_);
  and (_14879_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and (_14880_, _12980_, _23946_);
  or (_04755_, _14880_, _14879_);
  and (_14881_, _05281_, _23649_);
  and (_14882_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_04759_, _14882_, _14881_);
  and (_14883_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_14884_, _13894_, _23649_);
  or (_04765_, _14884_, _14883_);
  and (_14885_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_14886_, _13894_, _23747_);
  or (_04777_, _14886_, _14885_);
  and (_14887_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_14888_, _12980_, _23707_);
  or (_27095_, _14888_, _14887_);
  and (_14889_, _02321_, _23824_);
  and (_14890_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  or (_04779_, _14890_, _14889_);
  and (_14891_, _02321_, _23747_);
  and (_14892_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or (_27139_, _14892_, _14891_);
  and (_14893_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_14894_, _12974_, _23778_);
  or (_04784_, _14894_, _14893_);
  and (_14895_, _02370_, _23707_);
  and (_14896_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_27067_, _14896_, _14895_);
  and (_14897_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and (_14898_, _12974_, _23824_);
  or (_04796_, _14898_, _14897_);
  and (_14899_, _04922_, _23824_);
  and (_14900_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or (_04798_, _14900_, _14899_);
  and (_14901_, _25739_, _23707_);
  and (_14902_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or (_04803_, _14902_, _14901_);
  and (_14903_, _06886_, _23656_);
  not (_14904_, _14903_);
  and (_14905_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  and (_14906_, _14903_, _23747_);
  or (_04808_, _14906_, _14905_);
  and (_14907_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  and (_14908_, _14903_, _23824_);
  or (_04815_, _14908_, _14907_);
  and (_14909_, _02321_, _23946_);
  and (_14910_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or (_04818_, _14910_, _14909_);
  and (_14911_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_14912_, _12974_, _23747_);
  or (_04824_, _14912_, _14911_);
  and (_14913_, _04922_, _24050_);
  and (_14914_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  or (_04827_, _14914_, _14913_);
  and (_14915_, _02321_, _23707_);
  and (_14916_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or (_27140_, _14916_, _14915_);
  and (_14917_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_14918_, _12974_, _24050_);
  or (_04837_, _14918_, _14917_);
  and (_14919_, _25748_, _23778_);
  and (_14920_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or (_04841_, _14920_, _14919_);
  and (_14921_, _09913_, _24050_);
  and (_14922_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_04844_, _14922_, _14921_);
  and (_14923_, _02321_, _24050_);
  and (_14924_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or (_04847_, _14924_, _14923_);
  and (_14925_, _24852_, _23946_);
  and (_14926_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or (_04849_, _14926_, _14925_);
  and (_14927_, _25748_, _23946_);
  and (_14928_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_04865_, _14928_, _14927_);
  and (_14929_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_14930_, _12974_, _23707_);
  or (_04868_, _14930_, _14929_);
  and (_14931_, _25748_, _23747_);
  and (_14932_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_04870_, _14932_, _14931_);
  and (_14933_, _07743_, _23824_);
  and (_14934_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  or (_04875_, _14934_, _14933_);
  and (_14935_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  and (_14936_, _12970_, _23778_);
  or (_27097_, _14936_, _14935_);
  and (_14937_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  and (_14939_, _14903_, _23649_);
  or (_04884_, _14939_, _14937_);
  and (_14940_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  and (_14941_, _12970_, _23824_);
  or (_04889_, _14941_, _14940_);
  and (_14942_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  and (_14943_, _14903_, _24050_);
  or (_04893_, _14943_, _14942_);
  and (_14944_, _24639_, _23898_);
  and (_14945_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_04899_, _14945_, _14944_);
  and (_14946_, _05350_, _23778_);
  and (_14947_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  or (_04902_, _14947_, _14946_);
  and (_14948_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  and (_14949_, _14903_, _23946_);
  or (_04904_, _14949_, _14948_);
  and (_14950_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  and (_14951_, _12970_, _23649_);
  or (_04906_, _14951_, _14950_);
  and (_14952_, _02200_, _24050_);
  and (_14953_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_04910_, _14953_, _14952_);
  and (_14954_, _09913_, _23649_);
  and (_14955_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_04912_, _14955_, _14954_);
  and (_14956_, _23911_, _23664_);
  and (_14957_, _14956_, _23649_);
  not (_14958_, _14956_);
  and (_14959_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_04916_, _14959_, _14957_);
  and (_14960_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  and (_14961_, _12970_, _23946_);
  or (_04921_, _14961_, _14960_);
  and (_14962_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  and (_14963_, _12970_, _23707_);
  or (_04923_, _14963_, _14962_);
  and (_14964_, _24639_, _23946_);
  and (_14965_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_27169_, _14965_, _14964_);
  and (_14966_, _14956_, _23707_);
  and (_14967_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_04930_, _14967_, _14966_);
  and (_14968_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  and (_14969_, _12941_, _23778_);
  or (_04932_, _14969_, _14968_);
  and (_14970_, _24639_, _23824_);
  and (_14971_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_04933_, _14971_, _14970_);
  and (_14972_, _12782_, _23946_);
  and (_14973_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_04951_, _14973_, _14972_);
  and (_14974_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  and (_14975_, _12941_, _23824_);
  or (_04954_, _14975_, _14974_);
  and (_14976_, _24639_, _23747_);
  and (_14977_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_04960_, _14977_, _14976_);
  and (_14978_, _08799_, _23649_);
  and (_14979_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  or (_04963_, _14979_, _14978_);
  and (_14980_, _23946_, _23665_);
  and (_14981_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or (_04971_, _14981_, _14980_);
  and (_14982_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  and (_14983_, _12941_, _23747_);
  or (_27101_, _14983_, _14982_);
  and (_14984_, _23824_, _23665_);
  and (_14985_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  or (_04975_, _14985_, _14984_);
  and (_14986_, _02107_, _23747_);
  and (_14987_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  or (_04986_, _14987_, _14986_);
  and (_14988_, _03300_, _23649_);
  and (_14989_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_04988_, _14989_, _14988_);
  and (_14990_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  and (_14991_, _12941_, _23946_);
  or (_04990_, _14991_, _14990_);
  and (_14992_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  and (_14993_, _12941_, _23707_);
  or (_04997_, _14993_, _14992_);
  and (_14994_, _02107_, _23824_);
  and (_14995_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or (_04999_, _14995_, _14994_);
  and (_14996_, _06886_, _25078_);
  not (_14997_, _14996_);
  and (_14998_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  and (_14999_, _14996_, _23946_);
  or (_05002_, _14999_, _14998_);
  and (_15000_, _01971_, _23747_);
  and (_15001_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  or (_05004_, _15001_, _15000_);
  and (_15002_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and (_15003_, _12935_, _23898_);
  or (_05010_, _15003_, _15002_);
  and (_15004_, _01808_, _23664_);
  and (_15005_, _15004_, _23824_);
  not (_15006_, _15004_);
  and (_15007_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_05015_, _15007_, _15005_);
  and (_15008_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  and (_15009_, _14996_, _23649_);
  or (_05021_, _15009_, _15008_);
  and (_15010_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  and (_15011_, _14996_, _23747_);
  or (_05040_, _15011_, _15010_);
  and (_15012_, _23664_, _23069_);
  and (_15013_, _15012_, _23778_);
  not (_15014_, _15012_);
  and (_15015_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_05043_, _15015_, _15013_);
  and (_15016_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_15017_, _12935_, _23824_);
  or (_05046_, _15017_, _15016_);
  and (_15018_, _02107_, _23707_);
  and (_15019_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or (_05048_, _15019_, _15018_);
  and (_15020_, _15004_, _24050_);
  and (_15021_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_05051_, _15021_, _15020_);
  and (_15022_, _15012_, _23946_);
  and (_15023_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_05056_, _15023_, _15022_);
  and (_15024_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and (_15025_, _12935_, _23747_);
  or (_05059_, _15025_, _15024_);
  and (_15026_, _15012_, _23824_);
  and (_15027_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_05062_, _15027_, _15026_);
  and (_15028_, _02107_, _24050_);
  and (_15029_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  or (_05069_, _15029_, _15028_);
  and (_15030_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and (_15031_, _12935_, _23946_);
  or (_05071_, _15031_, _15030_);
  and (_15032_, _12733_, _23898_);
  and (_15033_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  or (_05076_, _15033_, _15032_);
  and (_15034_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_15035_, _12935_, _23707_);
  or (_05078_, _15035_, _15034_);
  and (_15036_, _05042_, _23898_);
  and (_15037_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_27134_, _15037_, _15036_);
  and (_15038_, _02107_, _23946_);
  and (_15039_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  or (_05082_, _15039_, _15038_);
  and (_15040_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_15041_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or (_15042_, _15041_, _15040_);
  and (_15043_, _15042_, _02393_);
  and (_15044_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and (_15045_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_15046_, _15045_, _15044_);
  and (_15047_, _15046_, _02445_);
  or (_15048_, _15047_, _15043_);
  and (_15049_, _15048_, _02421_);
  and (_15050_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_15051_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or (_15052_, _15051_, _15050_);
  and (_15053_, _15052_, _02393_);
  and (_15054_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and (_15055_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_15056_, _15055_, _15054_);
  and (_15057_, _15056_, _02445_);
  or (_15058_, _15057_, _15053_);
  and (_15059_, _15058_, _02459_);
  or (_15060_, _15059_, _15049_);
  and (_15061_, _15060_, _02458_);
  or (_15062_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or (_15063_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_15064_, _15063_, _15062_);
  and (_15065_, _15064_, _02393_);
  or (_15066_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or (_15067_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_15068_, _15067_, _15066_);
  and (_15069_, _15068_, _02445_);
  or (_15070_, _15069_, _15065_);
  and (_15071_, _15070_, _02421_);
  or (_15072_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_15073_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and (_15074_, _15073_, _15072_);
  and (_15075_, _15074_, _02393_);
  or (_15076_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or (_15077_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_15078_, _15077_, _15076_);
  and (_15079_, _15078_, _02445_);
  or (_15080_, _15079_, _15075_);
  and (_15081_, _15080_, _02459_);
  or (_15082_, _15081_, _15071_);
  and (_15083_, _15082_, _02414_);
  or (_15084_, _15083_, _15061_);
  and (_15085_, _15084_, _02398_);
  and (_15086_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and (_15087_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_15088_, _15087_, _15086_);
  and (_15089_, _15088_, _02393_);
  and (_15090_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and (_15091_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_15092_, _15091_, _15090_);
  and (_15093_, _15092_, _02445_);
  or (_15094_, _15093_, _15089_);
  and (_15095_, _15094_, _02421_);
  and (_15096_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and (_15097_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_15098_, _15097_, _15096_);
  and (_15099_, _15098_, _02393_);
  and (_15100_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and (_15101_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_15102_, _15101_, _15100_);
  and (_15103_, _15102_, _02445_);
  or (_15104_, _15103_, _15099_);
  and (_15105_, _15104_, _02459_);
  or (_15106_, _15105_, _15095_);
  and (_15107_, _15106_, _02458_);
  or (_15108_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_15109_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and (_15110_, _15109_, _02445_);
  and (_15111_, _15110_, _15108_);
  or (_15112_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_15113_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and (_15114_, _15113_, _02393_);
  and (_15115_, _15114_, _15112_);
  or (_15116_, _15115_, _15111_);
  and (_15117_, _15116_, _02421_);
  or (_15118_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_15119_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and (_15120_, _15119_, _02445_);
  and (_15121_, _15120_, _15118_);
  or (_15122_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_15123_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and (_15124_, _15123_, _02393_);
  and (_15125_, _15124_, _15122_);
  or (_15126_, _15125_, _15121_);
  and (_15127_, _15126_, _02459_);
  or (_15128_, _15127_, _15117_);
  and (_15129_, _15128_, _02414_);
  or (_15130_, _15129_, _15107_);
  and (_15131_, _15130_, _02496_);
  or (_15133_, _15131_, _15085_);
  and (_15134_, _15133_, _02400_);
  and (_15135_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_15136_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or (_15137_, _15136_, _15135_);
  and (_15138_, _15137_, _02393_);
  and (_15139_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_15140_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or (_15141_, _15140_, _15139_);
  and (_15142_, _15141_, _02445_);
  or (_15143_, _15142_, _15138_);
  or (_15144_, _15143_, _02459_);
  and (_15145_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_15146_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or (_15147_, _15146_, _15145_);
  and (_15148_, _15147_, _02393_);
  and (_15149_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_15150_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or (_15151_, _15150_, _15149_);
  and (_15152_, _15151_, _02445_);
  or (_15154_, _15152_, _15148_);
  or (_15155_, _15154_, _02421_);
  and (_15156_, _15155_, _02458_);
  and (_15157_, _15156_, _15144_);
  or (_15158_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or (_15159_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_15160_, _15159_, _02445_);
  and (_15161_, _15160_, _15158_);
  or (_15162_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or (_15163_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_15164_, _15163_, _02393_);
  and (_15165_, _15164_, _15162_);
  or (_15166_, _15165_, _15161_);
  or (_15167_, _15166_, _02459_);
  or (_15168_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or (_15169_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_15170_, _15169_, _02445_);
  and (_15171_, _15170_, _15168_);
  or (_15172_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or (_15173_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_15174_, _15173_, _02393_);
  and (_15175_, _15174_, _15172_);
  or (_15176_, _15175_, _15171_);
  or (_15177_, _15176_, _02421_);
  and (_15178_, _15177_, _02414_);
  and (_15179_, _15178_, _15167_);
  or (_15180_, _15179_, _15157_);
  and (_15181_, _15180_, _02496_);
  and (_15182_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and (_15183_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_15184_, _15183_, _15182_);
  and (_15185_, _15184_, _02393_);
  and (_15186_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and (_15187_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_15188_, _15187_, _15186_);
  and (_15189_, _15188_, _02445_);
  or (_15190_, _15189_, _15185_);
  or (_15191_, _15190_, _02459_);
  and (_15192_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and (_15193_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_15194_, _15193_, _15192_);
  and (_15195_, _15194_, _02393_);
  and (_15196_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and (_15197_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_15198_, _15197_, _15196_);
  and (_15199_, _15198_, _02445_);
  or (_15200_, _15199_, _15195_);
  or (_15201_, _15200_, _02421_);
  and (_15202_, _15201_, _02458_);
  and (_15203_, _15202_, _15191_);
  or (_15204_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_15205_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and (_15206_, _15205_, _15204_);
  and (_15207_, _15206_, _02393_);
  or (_15208_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_15209_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and (_15210_, _15209_, _15208_);
  and (_15211_, _15210_, _02445_);
  or (_15212_, _15211_, _15207_);
  or (_15213_, _15212_, _02459_);
  or (_15214_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_15215_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and (_15216_, _15215_, _15214_);
  and (_15217_, _15216_, _02393_);
  or (_15218_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_15219_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and (_15220_, _15219_, _15218_);
  and (_15221_, _15220_, _02445_);
  or (_15222_, _15221_, _15217_);
  or (_15223_, _15222_, _02421_);
  and (_15224_, _15223_, _02414_);
  and (_15225_, _15224_, _15213_);
  or (_15226_, _15225_, _15203_);
  and (_15227_, _15226_, _02398_);
  or (_15228_, _15227_, _15181_);
  and (_15229_, _15228_, _02546_);
  or (_15230_, _15229_, _15134_);
  and (_15231_, _15230_, _02646_);
  and (_15232_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and (_15233_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_15234_, _15233_, _15232_);
  and (_15235_, _15234_, _02445_);
  and (_15236_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and (_15237_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_15238_, _15237_, _15236_);
  and (_15239_, _15238_, _02393_);
  or (_15240_, _15239_, _15235_);
  or (_15241_, _15240_, _02459_);
  and (_15242_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and (_15243_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_15244_, _15243_, _15242_);
  and (_15245_, _15244_, _02445_);
  and (_15246_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and (_15247_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_15248_, _15247_, _15246_);
  and (_15249_, _15248_, _02393_);
  or (_15250_, _15249_, _15245_);
  or (_15251_, _15250_, _02421_);
  and (_15252_, _15251_, _02458_);
  and (_15253_, _15252_, _15241_);
  or (_15254_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_15255_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and (_15256_, _15255_, _02393_);
  and (_15257_, _15256_, _15254_);
  or (_15258_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_15259_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and (_15260_, _15259_, _02445_);
  and (_15261_, _15260_, _15258_);
  or (_15262_, _15261_, _15257_);
  or (_15263_, _15262_, _02459_);
  or (_15264_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_15265_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and (_15266_, _15265_, _02393_);
  and (_15267_, _15266_, _15264_);
  or (_15268_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_15269_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and (_15270_, _15269_, _02445_);
  and (_15271_, _15270_, _15268_);
  or (_15272_, _15271_, _15267_);
  or (_15273_, _15272_, _02421_);
  and (_15274_, _15273_, _02414_);
  and (_15275_, _15274_, _15263_);
  or (_15276_, _15275_, _15253_);
  or (_15277_, _15276_, _02398_);
  and (_15278_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and (_15279_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_15280_, _15279_, _02393_);
  or (_15281_, _15280_, _15278_);
  and (_15282_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_15283_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_15284_, _15283_, _02445_);
  or (_15285_, _15284_, _15282_);
  and (_15286_, _15285_, _15281_);
  or (_15287_, _15286_, _02459_);
  and (_15288_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and (_15289_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_15290_, _15289_, _02393_);
  or (_15291_, _15290_, _15288_);
  and (_15292_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and (_15293_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_15294_, _15293_, _02445_);
  or (_15295_, _15294_, _15292_);
  and (_15296_, _15295_, _15291_);
  or (_15297_, _15296_, _02421_);
  and (_15298_, _15297_, _02458_);
  and (_15299_, _15298_, _15287_);
  or (_15300_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_15301_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and (_15302_, _15301_, _15300_);
  or (_15303_, _15302_, _02445_);
  or (_15304_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_15305_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and (_15306_, _15305_, _15304_);
  or (_15307_, _15306_, _02393_);
  and (_15308_, _15307_, _15303_);
  or (_15309_, _15308_, _02459_);
  or (_15310_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_15311_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_15312_, _15311_, _15310_);
  or (_15313_, _15312_, _02445_);
  or (_15314_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_15315_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and (_15316_, _15315_, _15314_);
  or (_15317_, _15316_, _02393_);
  and (_15318_, _15317_, _15313_);
  or (_15319_, _15318_, _02421_);
  and (_15320_, _15319_, _02414_);
  and (_15321_, _15320_, _15309_);
  or (_15322_, _15321_, _15299_);
  or (_15323_, _15322_, _02496_);
  and (_15324_, _15323_, _02546_);
  and (_15325_, _15324_, _15277_);
  and (_15326_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  and (_15327_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or (_15328_, _15327_, _15326_);
  and (_15329_, _15328_, _02393_);
  and (_15330_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  and (_15331_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or (_15332_, _15331_, _15330_);
  and (_15333_, _15332_, _02445_);
  or (_15334_, _15333_, _15329_);
  and (_15335_, _15334_, _02421_);
  and (_15336_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  and (_15337_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or (_15338_, _15337_, _15336_);
  and (_15339_, _15338_, _02393_);
  and (_15340_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  and (_15341_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or (_15342_, _15341_, _15340_);
  and (_15343_, _15342_, _02445_);
  or (_15344_, _15343_, _15339_);
  and (_15345_, _15344_, _02459_);
  or (_15346_, _15345_, _15335_);
  and (_15347_, _15346_, _02458_);
  or (_15348_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or (_15349_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  and (_15350_, _15349_, _15348_);
  and (_15351_, _15350_, _02393_);
  or (_15352_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or (_15353_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  and (_15354_, _15353_, _15352_);
  and (_15355_, _15354_, _02445_);
  or (_15356_, _15355_, _15351_);
  and (_15357_, _15356_, _02421_);
  or (_15358_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or (_15359_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  and (_15360_, _15359_, _15358_);
  and (_15361_, _15360_, _02393_);
  or (_15362_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or (_15363_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  and (_15364_, _15363_, _15362_);
  and (_15365_, _15364_, _02445_);
  or (_15366_, _15365_, _15361_);
  and (_15367_, _15366_, _02459_);
  or (_15368_, _15367_, _15357_);
  and (_15369_, _15368_, _02414_);
  or (_15370_, _15369_, _15347_);
  and (_15371_, _15370_, _02496_);
  and (_15372_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_15373_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_15374_, _15373_, _15372_);
  and (_15375_, _15374_, _02393_);
  and (_15376_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_15377_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or (_15378_, _15377_, _15376_);
  and (_15379_, _15378_, _02445_);
  or (_15380_, _15379_, _15375_);
  and (_15381_, _15380_, _02421_);
  and (_15382_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_15383_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or (_15384_, _15383_, _15382_);
  and (_15385_, _15384_, _02393_);
  and (_15386_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_15387_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_15388_, _15387_, _15386_);
  and (_15389_, _15388_, _02445_);
  or (_15390_, _15389_, _15385_);
  and (_15391_, _15390_, _02459_);
  or (_15392_, _15391_, _15381_);
  and (_15393_, _15392_, _02458_);
  or (_15394_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_15395_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_15396_, _15395_, _15394_);
  and (_15397_, _15396_, _02393_);
  or (_15398_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or (_15399_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_15400_, _15399_, _15398_);
  and (_15401_, _15400_, _02445_);
  or (_15402_, _15401_, _15397_);
  and (_15403_, _15402_, _02421_);
  or (_15404_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_15405_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_15406_, _15405_, _15404_);
  and (_15407_, _15406_, _02393_);
  or (_15408_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or (_15409_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_15410_, _15409_, _15408_);
  and (_15411_, _15410_, _02445_);
  or (_15412_, _15411_, _15407_);
  and (_15413_, _15412_, _02459_);
  or (_15414_, _15413_, _15403_);
  and (_15415_, _15414_, _02414_);
  or (_15416_, _15415_, _15393_);
  and (_15417_, _15416_, _02398_);
  or (_15418_, _15417_, _15371_);
  and (_15419_, _15418_, _02400_);
  or (_15420_, _15419_, _15325_);
  and (_15421_, _15420_, _02405_);
  or (_15422_, _15421_, _15231_);
  and (_15423_, _15422_, _26777_);
  and (_15424_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and (_15425_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_15426_, _15425_, _15424_);
  and (_15427_, _15426_, _02445_);
  and (_15428_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and (_15429_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_15430_, _15429_, _15428_);
  and (_15431_, _15430_, _02393_);
  or (_15432_, _15431_, _15427_);
  or (_15433_, _15432_, _02459_);
  and (_15434_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and (_15435_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_15436_, _15435_, _15434_);
  and (_15437_, _15436_, _02445_);
  and (_15438_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and (_15439_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_15440_, _15439_, _15438_);
  and (_15441_, _15440_, _02393_);
  or (_15442_, _15441_, _15437_);
  or (_15443_, _15442_, _02421_);
  and (_15444_, _15443_, _02458_);
  and (_15445_, _15444_, _15433_);
  or (_15446_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_15447_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and (_15448_, _15447_, _02393_);
  and (_15449_, _15448_, _15446_);
  or (_15450_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_15451_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and (_15452_, _15451_, _02445_);
  and (_15453_, _15452_, _15450_);
  or (_15454_, _15453_, _15449_);
  or (_15455_, _15454_, _02459_);
  or (_15456_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_15457_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and (_15458_, _15457_, _02393_);
  and (_15459_, _15458_, _15456_);
  or (_15460_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_15461_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and (_15462_, _15461_, _02445_);
  and (_15463_, _15462_, _15460_);
  or (_15464_, _15463_, _15459_);
  or (_15465_, _15464_, _02421_);
  and (_15466_, _15465_, _02414_);
  and (_15467_, _15466_, _15455_);
  or (_15468_, _15467_, _15445_);
  and (_15469_, _15468_, _02496_);
  and (_15470_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and (_15471_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_15472_, _15471_, _02393_);
  or (_15473_, _15472_, _15470_);
  and (_15474_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and (_15475_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_15476_, _15475_, _02445_);
  or (_15477_, _15476_, _15474_);
  and (_15478_, _15477_, _15473_);
  or (_15479_, _15478_, _02459_);
  and (_15480_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and (_15481_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_15482_, _15481_, _02393_);
  or (_15483_, _15482_, _15480_);
  and (_15484_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and (_15485_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_15486_, _15485_, _02445_);
  or (_15487_, _15486_, _15484_);
  and (_15488_, _15487_, _15483_);
  or (_15489_, _15488_, _02421_);
  and (_15490_, _15489_, _02458_);
  and (_15491_, _15490_, _15479_);
  or (_15492_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_15493_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and (_15494_, _15493_, _15492_);
  or (_15495_, _15494_, _02445_);
  or (_15496_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_15497_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and (_15498_, _15497_, _15496_);
  or (_15499_, _15498_, _02393_);
  and (_15500_, _15499_, _15495_);
  or (_15501_, _15500_, _02459_);
  or (_15502_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_15503_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and (_15504_, _15503_, _15502_);
  or (_15505_, _15504_, _02445_);
  or (_15506_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_15507_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and (_15508_, _15507_, _15506_);
  or (_15509_, _15508_, _02393_);
  and (_15510_, _15509_, _15505_);
  or (_15511_, _15510_, _02421_);
  and (_15512_, _15511_, _02414_);
  and (_15513_, _15512_, _15501_);
  or (_15514_, _15513_, _15491_);
  and (_15515_, _15514_, _02398_);
  or (_15516_, _15515_, _15469_);
  and (_15517_, _15516_, _02546_);
  and (_15518_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and (_15519_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_15520_, _15519_, _15518_);
  and (_15521_, _15520_, _02393_);
  and (_15522_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and (_15523_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_15524_, _15523_, _15522_);
  and (_15525_, _15524_, _02445_);
  or (_15526_, _15525_, _15521_);
  and (_15527_, _15526_, _02421_);
  and (_15528_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and (_15529_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_15530_, _15529_, _15528_);
  and (_15531_, _15530_, _02393_);
  and (_15532_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and (_15533_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_15534_, _15533_, _15532_);
  and (_15535_, _15534_, _02445_);
  or (_15536_, _15535_, _15531_);
  and (_15537_, _15536_, _02459_);
  or (_15538_, _15537_, _15527_);
  and (_15539_, _15538_, _02458_);
  or (_15540_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_15541_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and (_15542_, _15541_, _15540_);
  and (_15543_, _15542_, _02393_);
  or (_15544_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_15545_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and (_15546_, _15545_, _15544_);
  and (_15547_, _15546_, _02445_);
  or (_15548_, _15547_, _15543_);
  and (_15549_, _15548_, _02421_);
  or (_15550_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_15551_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and (_15552_, _15551_, _15550_);
  and (_15553_, _15552_, _02393_);
  or (_15554_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_15555_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and (_15556_, _15555_, _15554_);
  and (_15557_, _15556_, _02445_);
  or (_15558_, _15557_, _15553_);
  and (_15559_, _15558_, _02459_);
  or (_15560_, _15559_, _15549_);
  and (_15561_, _15560_, _02414_);
  or (_15562_, _15561_, _15539_);
  and (_15563_, _15562_, _02398_);
  and (_15564_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_15565_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_15566_, _15565_, _15564_);
  and (_15567_, _15566_, _02393_);
  and (_15568_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_15569_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_15570_, _15569_, _15568_);
  and (_15571_, _15570_, _02445_);
  or (_15572_, _15571_, _15567_);
  and (_15573_, _15572_, _02421_);
  and (_15574_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_15575_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_15576_, _15575_, _15574_);
  and (_15577_, _15576_, _02393_);
  and (_15578_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_15579_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_15580_, _15579_, _15578_);
  and (_15581_, _15580_, _02445_);
  or (_15582_, _15581_, _15577_);
  and (_15583_, _15582_, _02459_);
  or (_15584_, _15583_, _15573_);
  and (_15585_, _15584_, _02458_);
  or (_15586_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_15587_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_15588_, _15587_, _15586_);
  and (_15589_, _15588_, _02393_);
  or (_15590_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_15591_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_15592_, _15591_, _15590_);
  and (_15593_, _15592_, _02445_);
  or (_15594_, _15593_, _15589_);
  and (_15595_, _15594_, _02421_);
  or (_15596_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_15597_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_15598_, _15597_, _15596_);
  and (_15599_, _15598_, _02393_);
  or (_15600_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_15601_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_15602_, _15601_, _15600_);
  and (_15603_, _15602_, _02445_);
  or (_15604_, _15603_, _15599_);
  and (_15605_, _15604_, _02459_);
  or (_15606_, _15605_, _15595_);
  and (_15607_, _15606_, _02414_);
  or (_15608_, _15607_, _15585_);
  and (_15609_, _15608_, _02496_);
  or (_15610_, _15609_, _15563_);
  and (_15611_, _15610_, _02400_);
  or (_15612_, _15611_, _15517_);
  and (_15613_, _15612_, _02646_);
  or (_15614_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_15615_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and (_15616_, _15615_, _02445_);
  and (_15617_, _15616_, _15614_);
  or (_15618_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or (_15619_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and (_15620_, _15619_, _02393_);
  and (_15621_, _15620_, _15618_);
  or (_15622_, _15621_, _15617_);
  and (_15623_, _15622_, _02459_);
  or (_15624_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_15625_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and (_15626_, _15625_, _02445_);
  and (_15627_, _15626_, _15624_);
  or (_15628_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or (_15629_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and (_15630_, _15629_, _02393_);
  and (_15631_, _15630_, _15628_);
  or (_15632_, _15631_, _15627_);
  and (_15633_, _15632_, _02421_);
  or (_15634_, _15633_, _15623_);
  and (_15635_, _15634_, _02414_);
  and (_15636_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and (_15637_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or (_15638_, _15637_, _15636_);
  and (_15639_, _15638_, _02393_);
  and (_15640_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and (_15641_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or (_15642_, _15641_, _15640_);
  and (_15643_, _15642_, _02445_);
  or (_15644_, _15643_, _15639_);
  and (_15645_, _15644_, _02459_);
  and (_15646_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and (_15647_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_15648_, _15647_, _15646_);
  and (_15649_, _15648_, _02393_);
  and (_15650_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and (_15651_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_15652_, _15651_, _15650_);
  and (_15653_, _15652_, _02445_);
  or (_15654_, _15653_, _15649_);
  and (_15655_, _15654_, _02421_);
  or (_15656_, _15655_, _15645_);
  and (_15657_, _15656_, _02458_);
  or (_15658_, _15657_, _15635_);
  and (_15659_, _15658_, _02496_);
  or (_15660_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_15661_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and (_15662_, _15661_, _15660_);
  and (_15663_, _15662_, _02393_);
  or (_15664_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_15665_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and (_15666_, _15665_, _15664_);
  and (_15667_, _15666_, _02445_);
  or (_15668_, _15667_, _15663_);
  and (_15669_, _15668_, _02459_);
  or (_15670_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_15671_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and (_15672_, _15671_, _15670_);
  and (_15673_, _15672_, _02393_);
  or (_15674_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_15675_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and (_15676_, _15675_, _15674_);
  and (_15677_, _15676_, _02445_);
  or (_15678_, _15677_, _15673_);
  and (_15679_, _15678_, _02421_);
  or (_15680_, _15679_, _15669_);
  and (_15681_, _15680_, _02414_);
  and (_15682_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and (_15683_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_15684_, _15683_, _15682_);
  and (_15685_, _15684_, _02393_);
  and (_15686_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and (_15687_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_15688_, _15687_, _15686_);
  and (_15689_, _15688_, _02445_);
  or (_15690_, _15689_, _15685_);
  and (_15691_, _15690_, _02459_);
  and (_15692_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and (_15693_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_15694_, _15693_, _15692_);
  and (_15695_, _15694_, _02393_);
  and (_15696_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and (_15697_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_15698_, _15697_, _15696_);
  and (_15699_, _15698_, _02445_);
  or (_15700_, _15699_, _15695_);
  and (_15701_, _15700_, _02421_);
  or (_15702_, _15701_, _15691_);
  and (_15703_, _15702_, _02458_);
  or (_15704_, _15703_, _15681_);
  and (_15705_, _15704_, _02398_);
  or (_15706_, _15705_, _15659_);
  and (_15707_, _15706_, _02400_);
  and (_15708_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and (_15709_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_15710_, _15709_, _15708_);
  and (_15711_, _15710_, _02393_);
  and (_15712_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and (_15713_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_15714_, _15713_, _15712_);
  and (_15715_, _15714_, _02445_);
  or (_15716_, _15715_, _15711_);
  or (_15717_, _15716_, _02459_);
  and (_15718_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and (_15719_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_15720_, _15719_, _15718_);
  and (_15721_, _15720_, _02393_);
  and (_15722_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and (_15723_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_15724_, _15723_, _15722_);
  and (_15725_, _15724_, _02445_);
  or (_15726_, _15725_, _15721_);
  or (_15727_, _15726_, _02421_);
  and (_15728_, _15727_, _02458_);
  and (_15729_, _15728_, _15717_);
  or (_15730_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_15731_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and (_15732_, _15731_, _15730_);
  and (_15733_, _15732_, _02393_);
  or (_15734_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_15735_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and (_15736_, _15735_, _15734_);
  and (_15737_, _15736_, _02445_);
  or (_15738_, _15737_, _15733_);
  or (_15739_, _15738_, _02459_);
  or (_15740_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_15741_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and (_15742_, _15741_, _15740_);
  and (_15743_, _15742_, _02393_);
  or (_15744_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_15745_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and (_15746_, _15745_, _15744_);
  and (_15747_, _15746_, _02445_);
  or (_15748_, _15747_, _15743_);
  or (_15749_, _15748_, _02421_);
  and (_15750_, _15749_, _02414_);
  and (_15751_, _15750_, _15739_);
  or (_15752_, _15751_, _15729_);
  and (_15753_, _15752_, _02398_);
  and (_15754_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and (_15755_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_15756_, _15755_, _15754_);
  and (_15757_, _15756_, _02393_);
  and (_15758_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and (_15759_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_15760_, _15759_, _15758_);
  and (_15761_, _15760_, _02445_);
  or (_15762_, _15761_, _15757_);
  or (_15763_, _15762_, _02459_);
  and (_15764_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and (_15765_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_15766_, _15765_, _15764_);
  and (_15767_, _15766_, _02393_);
  and (_15768_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and (_15769_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_15770_, _15769_, _15768_);
  and (_15771_, _15770_, _02445_);
  or (_15772_, _15771_, _15767_);
  or (_15773_, _15772_, _02421_);
  and (_15774_, _15773_, _02458_);
  and (_15775_, _15774_, _15763_);
  or (_15776_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_15777_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and (_15778_, _15777_, _02445_);
  and (_15779_, _15778_, _15776_);
  or (_15780_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_15781_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and (_15782_, _15781_, _02393_);
  and (_15783_, _15782_, _15780_);
  or (_15785_, _15783_, _15779_);
  or (_15786_, _15785_, _02459_);
  or (_15787_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_15788_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and (_15789_, _15788_, _02445_);
  and (_15790_, _15789_, _15787_);
  or (_15791_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_15792_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and (_15793_, _15792_, _02393_);
  and (_15794_, _15793_, _15791_);
  or (_15795_, _15794_, _15790_);
  or (_15796_, _15795_, _02421_);
  and (_15797_, _15796_, _02414_);
  and (_15798_, _15797_, _15786_);
  or (_15799_, _15798_, _15775_);
  and (_15800_, _15799_, _02496_);
  or (_15801_, _15800_, _15753_);
  and (_15802_, _15801_, _02546_);
  or (_15803_, _15802_, _15707_);
  and (_15804_, _15803_, _02405_);
  or (_15805_, _15804_, _15613_);
  and (_15806_, _15805_, _02444_);
  or (_15807_, _15806_, _15423_);
  or (_15808_, _15807_, _02443_);
  or (_15809_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_15810_, _15809_, _22762_);
  and (_05084_, _15810_, _15808_);
  and (_15811_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  and (_15812_, _14996_, _24050_);
  or (_05092_, _15812_, _15811_);
  and (_15813_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  and (_15814_, _14903_, _23778_);
  or (_05094_, _15814_, _15813_);
  and (_15815_, _08360_, _23707_);
  and (_15816_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or (_05103_, _15816_, _15815_);
  and (_15817_, _08360_, _23649_);
  and (_15818_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  or (_05106_, _15818_, _15817_);
  and (_15819_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_15820_, _12927_, _23898_);
  or (_05108_, _15820_, _15819_);
  and (_15821_, _08198_, _23824_);
  and (_15822_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_05112_, _15822_, _15821_);
  and (_15823_, _05701_, _23824_);
  and (_15824_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_05115_, _15824_, _15823_);
  and (_15825_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_15826_, _12927_, _23824_);
  or (_27104_, _15826_, _15825_);
  nand (_15827_, _24402_, _22767_);
  or (_15828_, _22767_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_15829_, _15828_, _22762_);
  and (_26864_[0], _15829_, _15827_);
  and (_15830_, _01808_, _24356_);
  and (_15831_, _15830_, _23946_);
  not (_15832_, _15830_);
  and (_15833_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or (_05123_, _15833_, _15831_);
  and (_15834_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  and (_15835_, _14996_, _23707_);
  or (_05124_, _15835_, _15834_);
  and (_15836_, _15830_, _23649_);
  and (_15837_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  or (_05136_, _15837_, _15836_);
  and (_15838_, _15830_, _23747_);
  and (_15839_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or (_05150_, _15839_, _15838_);
  and (_15840_, _15830_, _23824_);
  and (_15841_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  or (_05155_, _15841_, _15840_);
  and (_15842_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and (_15843_, _12829_, _23707_);
  or (_05179_, _15843_, _15842_);
  and (_15844_, _02107_, _23778_);
  and (_15845_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or (_27165_, _15845_, _15844_);
  and (_15846_, _06886_, _24282_);
  not (_15847_, _15846_);
  and (_15848_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_15849_, _15846_, _23649_);
  or (_27005_, _15849_, _15848_);
  and (_15850_, _23752_, _23076_);
  and (_15851_, _15850_, _23824_);
  not (_15852_, _15850_);
  and (_15853_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or (_05185_, _15853_, _15851_);
  and (_15854_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_15855_, _15846_, _24050_);
  or (_27006_, _15855_, _15854_);
  not (_15856_, _26110_);
  nor (_15857_, _15856_, _24299_);
  or (_15858_, _15857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_15859_, _26114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_15860_, _15859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_15861_, _15860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_15862_, _15861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_15863_, _15862_, _26100_);
  nand (_15864_, _15863_, _12811_);
  or (_15865_, _15864_, _24299_);
  and (_15866_, _15865_, _15858_);
  or (_15867_, _15866_, _24293_);
  nand (_15868_, _24293_, _23772_);
  and (_15869_, _15868_, _22762_);
  and (_05196_, _15869_, _15867_);
  and (_15870_, _15830_, _23707_);
  and (_15871_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  or (_05198_, _15871_, _15870_);
  and (_15872_, _15830_, _24050_);
  and (_15873_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or (_05202_, _15873_, _15872_);
  nand (_15874_, _24508_, _22767_);
  or (_15875_, _22767_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_15876_, _15875_, _22762_);
  and (_26864_[7], _15876_, _15874_);
  and (_15877_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and (_15878_, _15846_, _23946_);
  or (_05220_, _15878_, _15877_);
  and (_15879_, _12733_, _23946_);
  and (_15880_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or (_05225_, _15880_, _15879_);
  and (_15881_, _15830_, _23898_);
  and (_15882_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or (_05232_, _15882_, _15881_);
  and (_15883_, _15830_, _23778_);
  and (_15884_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  or (_27164_, _15884_, _15883_);
  and (_15885_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  and (_15886_, _14996_, _23778_);
  or (_27007_, _15886_, _15885_);
  and (_15887_, _05187_, _23946_);
  and (_15888_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_05274_, _15888_, _15887_);
  and (_15889_, _05187_, _23649_);
  and (_15890_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_05280_, _15890_, _15889_);
  and (_15891_, _05187_, _23747_);
  and (_15892_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_05287_, _15892_, _15891_);
  and (_15893_, _15850_, _23649_);
  and (_15894_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or (_05300_, _15894_, _15893_);
  and (_15895_, _24201_, _23784_);
  not (_15896_, _15895_);
  and (_15897_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  and (_15898_, _15895_, _23707_);
  or (_05306_, _15898_, _15897_);
  and (_15899_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_15900_, _15846_, _23707_);
  or (_05312_, _15900_, _15899_);
  and (_15901_, _05114_, _23778_);
  and (_15902_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_05321_, _15902_, _15901_);
  and (_15903_, _05187_, _23707_);
  and (_15904_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_05341_, _15904_, _15903_);
  and (_15905_, _05187_, _24050_);
  and (_15906_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_27099_, _15906_, _15905_);
  and (_15907_, _06886_, _23911_);
  not (_15908_, _15907_);
  and (_15909_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_15910_, _15907_, _23707_);
  or (_27003_, _15910_, _15909_);
  and (_15911_, _24358_, _23707_);
  and (_15912_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or (_05370_, _15912_, _15911_);
  and (_15913_, _24331_, _23946_);
  and (_15914_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_05383_, _15914_, _15913_);
  and (_15915_, _24358_, _24050_);
  and (_15916_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or (_05386_, _15916_, _15915_);
  and (_15917_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  and (_15918_, _15895_, _24050_);
  or (_05389_, _15918_, _15917_);
  and (_15919_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and (_15920_, _15846_, _23824_);
  or (_05406_, _15920_, _15919_);
  and (_15921_, _05187_, _23898_);
  and (_15922_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_05408_, _15922_, _15921_);
  and (_15923_, _05187_, _23778_);
  and (_15924_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_05418_, _15924_, _15923_);
  and (_15925_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_15926_, _15846_, _23898_);
  or (_05421_, _15926_, _15925_);
  and (_15927_, _04811_, _23747_);
  and (_15928_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  or (_05423_, _15928_, _15927_);
  and (_15929_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and (_15930_, _01967_, _23898_);
  or (_27233_, _15930_, _15929_);
  and (_15931_, _23790_, _23778_);
  and (_15932_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  or (_27252_, _15932_, _15931_);
  and (_15933_, _05114_, _23649_);
  and (_15934_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_05451_, _15934_, _15933_);
  and (_15935_, _05114_, _23747_);
  and (_15936_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_05456_, _15936_, _15935_);
  and (_15937_, _05114_, _23824_);
  and (_15938_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_05465_, _15938_, _15937_);
  and (_15939_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_15940_, _15907_, _23898_);
  or (_05473_, _15940_, _15939_);
  and (_15941_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and (_15942_, _15907_, _23778_);
  or (_05476_, _15942_, _15941_);
  and (_15943_, _09913_, _23707_);
  and (_15944_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_05479_, _15944_, _15943_);
  and (_15945_, _05114_, _24050_);
  and (_15946_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_05498_, _15946_, _15945_);
  and (_15947_, _05114_, _23946_);
  and (_15948_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_05503_, _15948_, _15947_);
  and (_15949_, _08360_, _23898_);
  and (_15950_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  or (_27086_, _15950_, _15949_);
  and (_15951_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and (_15952_, _15907_, _23649_);
  or (_27001_, _15952_, _15951_);
  and (_15953_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_15954_, _15907_, _23747_);
  or (_27000_, _15954_, _15953_);
  and (_15955_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  and (_15956_, _05337_, _23898_);
  or (_05542_, _15956_, _15955_);
  and (_15957_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and (_15958_, _12927_, _23707_);
  or (_05543_, _15958_, _15957_);
  and (_15959_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  and (_15960_, _08477_, _23898_);
  or (_05546_, _15960_, _15959_);
  and (_15961_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and (_15962_, _05398_, _24050_);
  or (_05549_, _15962_, _15961_);
  and (_15963_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and (_15964_, _05358_, _23778_);
  or (_05557_, _15964_, _15963_);
  and (_15965_, _05371_, _23824_);
  and (_15966_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_05568_, _15966_, _15965_);
  and (_15967_, _08360_, _23778_);
  and (_15968_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or (_05570_, _15968_, _15967_);
  and (_15969_, _05371_, _23649_);
  and (_15970_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_05573_, _15970_, _15969_);
  and (_15971_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_15972_, _13777_, _23778_);
  or (_05577_, _15972_, _15971_);
  and (_15973_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  and (_15974_, _05358_, _23747_);
  or (_05584_, _15974_, _15973_);
  and (_15975_, _06886_, _24010_);
  not (_15976_, _15975_);
  and (_15977_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  and (_15978_, _15975_, _23747_);
  or (_05589_, _15978_, _15977_);
  and (_15979_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  and (_15980_, _05354_, _23824_);
  or (_05598_, _15980_, _15979_);
  and (_15981_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_15982_, _05705_, _23898_);
  or (_05622_, _15982_, _15981_);
  and (_15983_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  and (_15984_, _05358_, _23824_);
  or (_05625_, _15984_, _15983_);
  and (_15985_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  and (_15986_, _05354_, _24050_);
  or (_05633_, _15986_, _15985_);
  and (_15987_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  and (_15988_, _12829_, _23824_);
  or (_05639_, _15988_, _15987_);
  and (_15989_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  and (_15990_, _05358_, _23649_);
  or (_05643_, _15990_, _15989_);
  and (_15991_, _04760_, _24085_);
  not (_15992_, _15991_);
  and (_15993_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  and (_15994_, _15991_, _24050_);
  or (_05659_, _15994_, _15993_);
  and (_15995_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  and (_15996_, _15991_, _23747_);
  or (_05661_, _15996_, _15995_);
  and (_15997_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and (_15998_, _12829_, _23898_);
  or (_27224_, _15998_, _15997_);
  and (_15999_, _24699_, _23778_);
  and (_16000_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or (_27189_, _16000_, _15999_);
  nand (_16001_, _25172_, _23662_);
  or (_16002_, _16001_, _00875_);
  not (_16003_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_16004_, _16001_, _16003_);
  and (_16005_, _16004_, _24069_);
  and (_16006_, _16005_, _16002_);
  nor (_16007_, _24068_, _16003_);
  and (_16008_, _00265_, _25163_);
  and (_16009_, _16008_, _24654_);
  nand (_16010_, _16009_, _23594_);
  or (_16011_, _16009_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_16012_, _16011_, _24645_);
  and (_16013_, _16012_, _16010_);
  or (_16014_, _16013_, _16007_);
  or (_16015_, _16014_, _16006_);
  and (_05678_, _16015_, _22762_);
  and (_16016_, _15850_, _23747_);
  and (_16017_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or (_05689_, _16017_, _16016_);
  and (_16018_, _04760_, _23986_);
  not (_16019_, _16018_);
  and (_16020_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  and (_16021_, _16018_, _23898_);
  or (_05700_, _16021_, _16020_);
  and (_16022_, _24370_, _23903_);
  and (_16023_, _16022_, _23649_);
  not (_16024_, _16022_);
  and (_16025_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_05707_, _16025_, _16023_);
  and (_16026_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_16027_, _12927_, _24050_);
  or (_05754_, _16027_, _16026_);
  and (_16028_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_16029_, _05398_, _23778_);
  or (_05769_, _16029_, _16028_);
  and (_16030_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  and (_16031_, _15991_, _23649_);
  or (_05784_, _16031_, _16030_);
  and (_16032_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and (_16033_, _12927_, _23649_);
  or (_05788_, _16033_, _16032_);
  and (_16034_, _05701_, _23946_);
  and (_16035_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_27087_, _16035_, _16034_);
  and (_16036_, _06665_, _24050_);
  and (_16037_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  or (_27089_, _16037_, _16036_);
  and (_16038_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_16039_, _12927_, _23946_);
  or (_05804_, _16039_, _16038_);
  and (_16040_, _24050_, _23833_);
  and (_16041_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_05815_, _16041_, _16040_);
  and (_16042_, _05371_, _23946_);
  and (_16043_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_05842_, _16043_, _16042_);
  and (_16044_, _05180_, _23898_);
  and (_16045_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_05849_, _16045_, _16044_);
  and (_16046_, _12733_, _23778_);
  and (_16047_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or (_05854_, _16047_, _16046_);
  and (_16048_, _04760_, _24010_);
  not (_16049_, _16048_);
  and (_16050_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  and (_16051_, _16048_, _23778_);
  or (_05862_, _16051_, _16050_);
  and (_16052_, _24121_, _23939_);
  nand (_16053_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_16054_, _16053_, _24127_);
  nor (_16055_, _24151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_16056_, _16055_, _12951_);
  nand (_16057_, _16056_, _12956_);
  or (_16058_, _12956_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_16059_, _16058_, _16057_);
  or (_16060_, _16059_, _16054_);
  and (_16061_, _16060_, _24166_);
  or (_05875_, _16061_, _16052_);
  and (_16062_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_16063_, _11746_, _24050_);
  or (_27029_, _16063_, _16062_);
  and (_16064_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_16065_, _11746_, _23824_);
  or (_27027_, _16065_, _16064_);
  and (_16066_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  and (_16067_, _15895_, _23778_);
  or (_27222_, _16067_, _16066_);
  and (_16068_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  and (_16069_, _16048_, _23898_);
  or (_05899_, _16069_, _16068_);
  and (_16070_, _15012_, _23707_);
  and (_16071_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_05905_, _16071_, _16070_);
  and (_16072_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  and (_16073_, _11729_, _23707_);
  or (_05907_, _16073_, _16072_);
  and (_16074_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  and (_16075_, _11729_, _23898_);
  or (_05915_, _16075_, _16074_);
  and (_16076_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_16077_, _11693_, _24050_);
  or (_05949_, _16077_, _16076_);
  and (_16078_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_16079_, _11693_, _23824_);
  or (_05956_, _16079_, _16078_);
  and (_16080_, _12782_, _23649_);
  and (_16081_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_05964_, _16081_, _16080_);
  and (_16082_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_16083_, _11693_, _23778_);
  or (_05968_, _16083_, _16082_);
  and (_16084_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  and (_16085_, _15975_, _23824_);
  or (_05971_, _16085_, _16084_);
  and (_16086_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_16087_, _11652_, _23707_);
  or (_05974_, _16087_, _16086_);
  and (_16088_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_16089_, _11652_, _23649_);
  or (_27025_, _16089_, _16088_);
  and (_16090_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  and (_16091_, _10494_, _23946_);
  or (_05987_, _16091_, _16090_);
  and (_16092_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  and (_16093_, _15975_, _23898_);
  or (_05991_, _16093_, _16092_);
  and (_16094_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and (_16095_, _10494_, _23824_);
  or (_05995_, _16095_, _16094_);
  and (_16096_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  and (_16097_, _08375_, _23707_);
  or (_06009_, _16097_, _16096_);
  and (_16098_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  and (_16099_, _08375_, _23824_);
  or (_06016_, _16099_, _16098_);
  and (_16100_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_16101_, _06896_, _23747_);
  or (_06023_, _16101_, _16100_);
  and (_16102_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  and (_16103_, _15975_, _24050_);
  or (_06031_, _16103_, _16102_);
  and (_16104_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  and (_16105_, _15975_, _23946_);
  or (_06041_, _16105_, _16104_);
  and (_16106_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  and (_16107_, _07551_, _23747_);
  or (_27019_, _16107_, _16106_);
  and (_16108_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  and (_16109_, _07525_, _24050_);
  or (_06051_, _16109_, _16108_);
  and (_16110_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  and (_16111_, _07525_, _23824_);
  or (_27018_, _16111_, _16110_);
  and (_16112_, _05180_, _23747_);
  and (_16113_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_27131_, _16113_, _16112_);
  and (_16114_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_16115_, _06927_, _23707_);
  or (_06077_, _16115_, _16114_);
  and (_16116_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_16117_, _06927_, _23747_);
  or (_06085_, _16117_, _16116_);
  and (_16118_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  and (_16119_, _16048_, _23824_);
  or (_06088_, _16119_, _16118_);
  and (_16120_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  and (_16121_, _16048_, _23649_);
  or (_06093_, _16121_, _16120_);
  and (_16122_, _06886_, _24085_);
  not (_16123_, _16122_);
  and (_16124_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  and (_16125_, _16122_, _23946_);
  or (_06098_, _16125_, _16124_);
  and (_16126_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_16127_, _06900_, _23707_);
  or (_06100_, _16127_, _16126_);
  and (_16128_, _24086_, _23778_);
  and (_16129_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_27254_, _16129_, _16128_);
  and (_16130_, _02359_, _23649_);
  and (_16131_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  or (_06103_, _16131_, _16130_);
  and (_16132_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_16133_, _06900_, _23649_);
  or (_27021_, _16133_, _16132_);
  and (_16134_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  and (_16135_, _16122_, _23649_);
  or (_06109_, _16135_, _16134_);
  and (_16136_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_16137_, _06896_, _23898_);
  or (_06112_, _16137_, _16136_);
  and (_16138_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  and (_16139_, _04748_, _23898_);
  or (_06116_, _16139_, _16138_);
  and (_16140_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  and (_16141_, _16018_, _23824_);
  or (_06121_, _16141_, _16140_);
  and (_16142_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  and (_16143_, _11729_, _23747_);
  or (_06123_, _16143_, _16142_);
  and (_16144_, _15012_, _24050_);
  and (_16145_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_06131_, _16145_, _16144_);
  and (_16146_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_16147_, _11693_, _23649_);
  or (_06134_, _16147_, _16146_);
  and (_16148_, _06639_, _23649_);
  and (_16149_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_06141_, _16149_, _16148_);
  and (_16150_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_16151_, _11652_, _23898_);
  or (_06151_, _16151_, _16150_);
  and (_16152_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  and (_16153_, _08375_, _23649_);
  or (_27023_, _16153_, _16152_);
  and (_16154_, _06639_, _24050_);
  and (_16155_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_06160_, _16155_, _16154_);
  and (_16156_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  and (_16157_, _08375_, _23778_);
  or (_06163_, _16157_, _16156_);
  and (_16158_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_16159_, _06896_, _23946_);
  or (_06168_, _16159_, _16158_);
  and (_16160_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_16161_, _06900_, _23778_);
  or (_06171_, _16161_, _16160_);
  and (_16162_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  and (_16163_, _16122_, _23707_);
  or (_06176_, _16163_, _16162_);
  and (_16164_, _06639_, _23946_);
  and (_16165_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_06178_, _16165_, _16164_);
  and (_16166_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  and (_16167_, _07551_, _23946_);
  or (_06180_, _16167_, _16166_);
  and (_16168_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  and (_16169_, _07551_, _23898_);
  or (_06184_, _16169_, _16168_);
  and (_16170_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_16171_, _06927_, _23778_);
  or (_06205_, _16171_, _16170_);
  or (_26862_[0], _05000_, _12899_);
  and (_16172_, _24283_, _23747_);
  and (_16173_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  or (_06233_, _16173_, _16172_);
  and (_16174_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_16175_, _11746_, _23747_);
  or (_27028_, _16175_, _16174_);
  and (_16176_, _23992_, _23824_);
  and (_16177_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_26944_, _16177_, _16176_);
  and (_16178_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_16179_, _11652_, _23946_);
  or (_06254_, _16179_, _16178_);
  and (_16180_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  and (_16181_, _10494_, _24050_);
  or (_06257_, _16181_, _16180_);
  and (_16182_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  and (_16183_, _16122_, _23778_);
  or (_06264_, _16183_, _16182_);
  and (_16184_, _25439_, _24118_);
  nand (_16185_, _16184_, _23594_);
  or (_16186_, _16184_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_16187_, _16186_, _24645_);
  and (_16188_, _16187_, _16185_);
  or (_16189_, _25447_, _23738_);
  or (_16190_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_16191_, _16190_, _24069_);
  and (_16192_, _16191_, _16189_);
  and (_16193_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_16194_, _16193_, rst);
  or (_16195_, _16194_, _16192_);
  or (_06267_, _16195_, _16188_);
  and (_16196_, _06886_, _23784_);
  not (_16197_, _16196_);
  and (_16198_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_16199_, _16196_, _23707_);
  or (_06271_, _16199_, _16198_);
  and (_16200_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  and (_16201_, _07525_, _23747_);
  or (_06273_, _16201_, _16200_);
  and (_16202_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_16203_, _06927_, _23649_);
  or (_06276_, _16203_, _16202_);
  and (_16204_, _25350_, _24296_);
  nand (_16205_, _16204_, _23594_);
  or (_16206_, _16204_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_16207_, _16206_, _24645_);
  and (_16208_, _16207_, _16205_);
  or (_16209_, _25359_, _23642_);
  or (_16210_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_16211_, _16210_, _24069_);
  and (_16212_, _16211_, _16209_);
  nor (_16213_, _24068_, _06249_);
  or (_16214_, _16213_, rst);
  or (_16215_, _16214_, _16212_);
  or (_06280_, _16215_, _16208_);
  and (_16216_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and (_16217_, _11729_, _23649_);
  or (_06289_, _16217_, _16216_);
  and (_16218_, _25260_, _24705_);
  nand (_16219_, _16218_, _23594_);
  or (_16220_, _16218_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_16221_, _16220_, _24645_);
  and (_16222_, _16221_, _16219_);
  or (_16223_, _25267_, _24043_);
  or (_16224_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_16225_, _16224_, _24069_);
  and (_16226_, _16225_, _16223_);
  nor (_16227_, _24068_, _06185_);
  or (_16228_, _16227_, rst);
  or (_16229_, _16228_, _16226_);
  or (_06293_, _16229_, _16222_);
  and (_16230_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_16231_, _06900_, _23898_);
  or (_27020_, _16231_, _16230_);
  and (_16232_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  and (_16233_, _16122_, _23824_);
  or (_26997_, _16233_, _16232_);
  and (_16234_, _25164_, _24296_);
  nand (_16235_, _16234_, _23594_);
  or (_16237_, _16234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_16238_, _16237_, _24645_);
  and (_16239_, _16238_, _16235_);
  or (_16240_, _25174_, _23642_);
  or (_16241_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_16242_, _16241_, _24069_);
  and (_16243_, _16242_, _16240_);
  nor (_16244_, _24068_, _06149_);
  or (_16245_, _16244_, rst);
  or (_16246_, _16245_, _16243_);
  or (_06326_, _16246_, _16239_);
  and (_16247_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  and (_16248_, _12728_, _24050_);
  or (_06332_, _16248_, _16247_);
  and (_16249_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_16250_, _12906_, _23824_);
  or (_06338_, _16250_, _16249_);
  and (_16251_, _05710_, _23707_);
  and (_16252_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  or (_06342_, _16252_, _16251_);
  and (_16253_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and (_16254_, _13756_, _23649_);
  or (_06360_, _16254_, _16253_);
  and (_16255_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  and (_16256_, _14903_, _23707_);
  or (_06364_, _16256_, _16255_);
  and (_16257_, _05710_, _24050_);
  and (_16258_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  or (_06368_, _16258_, _16257_);
  and (_16259_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  and (_16260_, _14903_, _23898_);
  or (_06370_, _16260_, _16259_);
  and (_16261_, _05710_, _23946_);
  and (_16262_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  or (_27163_, _16262_, _16261_);
  and (_16263_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_16264_, _15907_, _23946_);
  or (_27002_, _16264_, _16263_);
  and (_16265_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_16266_, _16196_, _23824_);
  or (_06386_, _16266_, _16265_);
  and (_16267_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  and (_16268_, _15975_, _23778_);
  or (_06391_, _16268_, _16267_);
  and (_16269_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  and (_16270_, _16122_, _23747_);
  or (_06395_, _16270_, _16269_);
  and (_16271_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_16272_, _16196_, _23946_);
  or (_06398_, _16272_, _16271_);
  and (_16273_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_16274_, _16196_, _23898_);
  or (_06401_, _16274_, _16273_);
  and (_16275_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_16276_, _16196_, _23778_);
  or (_06403_, _16276_, _16275_);
  and (_16277_, _06506_, _23991_);
  not (_16278_, _16277_);
  and (_16279_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  and (_16280_, _16277_, _23824_);
  or (_06415_, _16280_, _16279_);
  and (_16281_, _06506_, _23903_);
  not (_16282_, _16281_);
  and (_16283_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  and (_16284_, _16281_, _23824_);
  or (_26995_, _16284_, _16283_);
  and (_16285_, _06506_, _24005_);
  not (_16286_, _16285_);
  and (_16287_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and (_16288_, _16285_, _23649_);
  or (_06430_, _16288_, _16287_);
  and (_16289_, _06506_, _23986_);
  not (_16290_, _16289_);
  and (_16291_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and (_16292_, _16289_, _23649_);
  or (_26991_, _16292_, _16291_);
  and (_16293_, _06506_, _23069_);
  not (_16294_, _16293_);
  and (_16295_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  and (_16296_, _16293_, _24050_);
  or (_06440_, _16296_, _16295_);
  and (_16297_, _06639_, _23778_);
  and (_16298_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_06446_, _16298_, _16297_);
  and (_16299_, _06506_, _24329_);
  not (_16300_, _16299_);
  and (_16301_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and (_16302_, _16299_, _23747_);
  or (_06450_, _16302_, _16301_);
  and (_16303_, _06506_, _23752_);
  not (_16304_, _16303_);
  and (_16305_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  and (_16306_, _16303_, _23778_);
  or (_06457_, _16306_, _16305_);
  and (_16307_, _06506_, _23656_);
  not (_16308_, _16307_);
  and (_16309_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and (_16310_, _16307_, _23747_);
  or (_06461_, _16310_, _16309_);
  and (_16311_, _06506_, _24085_);
  not (_16312_, _16311_);
  and (_16313_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and (_16314_, _16311_, _24050_);
  or (_06468_, _16314_, _16313_);
  and (_16315_, _06639_, _23898_);
  and (_16316_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_06470_, _16316_, _16315_);
  and (_16317_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_16318_, _16196_, _23649_);
  or (_06473_, _16318_, _16317_);
  and (_16319_, _04760_, _24275_);
  not (_16320_, _16319_);
  and (_16321_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  and (_16322_, _16319_, _24050_);
  or (_06484_, _16322_, _16321_);
  and (_16323_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_16324_, _16196_, _23747_);
  or (_06492_, _16324_, _16323_);
  and (_16325_, _04760_, _23903_);
  not (_16326_, _16325_);
  and (_16327_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and (_16328_, _16325_, _23946_);
  or (_26968_, _16328_, _16327_);
  and (_16329_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and (_16330_, _16325_, _23898_);
  or (_06512_, _16330_, _16329_);
  and (_16331_, _04760_, _24005_);
  not (_16332_, _16331_);
  and (_16333_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  and (_16334_, _16331_, _23946_);
  or (_06516_, _16334_, _16333_);
  and (_16335_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  and (_16336_, _16018_, _23707_);
  or (_06519_, _16336_, _16335_);
  and (_16337_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  and (_16338_, _16018_, _23747_);
  or (_06521_, _16338_, _16337_);
  and (_16339_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and (_16340_, _07513_, _24050_);
  or (_06523_, _16340_, _16339_);
  and (_16341_, _23992_, _23747_);
  and (_16342_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_06526_, _16342_, _16341_);
  and (_16343_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and (_16344_, _04761_, _23747_);
  or (_06528_, _16344_, _16343_);
  and (_16345_, _23992_, _23649_);
  and (_16346_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_06535_, _16346_, _16345_);
  and (_16347_, _24050_, _23992_);
  and (_16348_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_06537_, _16348_, _16347_);
  and (_16349_, _24275_, _23906_);
  and (_16350_, _16349_, _23778_);
  not (_16351_, _16349_);
  and (_16352_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  or (_06543_, _16352_, _16350_);
  and (_16353_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  and (_16354_, _13828_, _24050_);
  or (_06546_, _16354_, _16353_);
  and (_16355_, _05714_, _23707_);
  and (_16356_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  or (_27160_, _16356_, _16355_);
  and (_16357_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  and (_16358_, _14996_, _23824_);
  or (_06549_, _16358_, _16357_);
  and (_16359_, _06506_, _24275_);
  not (_16360_, _16359_);
  and (_16361_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and (_16362_, _16359_, _23824_);
  or (_06556_, _16362_, _16361_);
  and (_16363_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and (_16364_, _16359_, _23649_);
  or (_06560_, _16364_, _16363_);
  and (_16365_, _05710_, _23778_);
  and (_16366_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  or (_06562_, _16366_, _16365_);
  and (_16367_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and (_16368_, _16359_, _23747_);
  or (_06565_, _16368_, _16367_);
  and (_16369_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and (_16370_, _16359_, _23898_);
  or (_06571_, _16370_, _16369_);
  and (_16371_, _06506_, _23784_);
  not (_16372_, _16371_);
  and (_16373_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  and (_16374_, _16371_, _23747_);
  or (_06591_, _16374_, _16373_);
  and (_16375_, _04760_, _23991_);
  not (_16376_, _16375_);
  and (_16377_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and (_16378_, _16375_, _23898_);
  or (_06595_, _16378_, _16377_);
  and (_16379_, _08167_, _23778_);
  and (_16380_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or (_06601_, _16380_, _16379_);
  and (_16381_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and (_16382_, _04761_, _23707_);
  or (_26962_, _16382_, _16381_);
  and (_16383_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  and (_16384_, _08477_, _23946_);
  or (_06611_, _16384_, _16383_);
  and (_16385_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and (_16386_, _06507_, _24050_);
  or (_26979_, _16386_, _16385_);
  and (_16387_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and (_16388_, _16359_, _24050_);
  or (_06617_, _16388_, _16387_);
  and (_16389_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and (_16390_, _15907_, _24050_);
  or (_06631_, _16390_, _16389_);
  and (_16391_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_16392_, _16196_, _24050_);
  or (_06633_, _16392_, _16391_);
  and (_16393_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  and (_16394_, _16281_, _23747_);
  or (_06635_, _16394_, _16393_);
  and (_16395_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  and (_16396_, _16303_, _23898_);
  or (_06638_, _16396_, _16395_);
  and (_16397_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and (_16398_, _16359_, _23707_);
  or (_06640_, _16398_, _16397_);
  and (_16399_, _08167_, _23824_);
  and (_16400_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  or (_06642_, _16400_, _16399_);
  and (_16401_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and (_16402_, _16311_, _23707_);
  or (_06645_, _16402_, _16401_);
  and (_16403_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  and (_16404_, _16319_, _23824_);
  or (_06648_, _16404_, _16403_);
  and (_16405_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  and (_16406_, _10331_, _23824_);
  or (_06660_, _16406_, _16405_);
  and (_16407_, _05710_, _23747_);
  and (_16408_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  or (_27161_, _16408_, _16407_);
  and (_16409_, _05710_, _23824_);
  and (_16410_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  or (_06664_, _16410_, _16409_);
  and (_16411_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  and (_16412_, _16277_, _23946_);
  or (_26996_, _16412_, _16411_);
  and (_16413_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and (_16414_, _10331_, _23898_);
  or (_26982_, _16414_, _16413_);
  and (_16415_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and (_16416_, _06507_, _23824_);
  or (_06679_, _16416_, _16415_);
  and (_16417_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and (_16418_, _06507_, _23778_);
  or (_06684_, _16418_, _16417_);
  and (_16419_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and (_16420_, _06507_, _23946_);
  or (_06689_, _16420_, _16419_);
  and (_16421_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  and (_16422_, _16277_, _23649_);
  or (_06695_, _16422_, _16421_);
  and (_16423_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and (_16424_, _06507_, _23707_);
  or (_06702_, _16424_, _16423_);
  and (_16425_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  and (_16426_, _08477_, _23649_);
  or (_06705_, _16426_, _16425_);
  and (_16427_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  and (_16428_, _16277_, _23747_);
  or (_06707_, _16428_, _16427_);
  and (_16429_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and (_16430_, _04761_, _23824_);
  or (_06709_, _16430_, _16429_);
  and (_16431_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and (_16432_, _04761_, _24050_);
  or (_06711_, _16432_, _16431_);
  and (_16433_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and (_16434_, _04761_, _23946_);
  or (_06714_, _16434_, _16433_);
  and (_16435_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and (_16436_, _07513_, _23824_);
  or (_26964_, _16436_, _16435_);
  and (_16437_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and (_16438_, _07513_, _23778_);
  or (_06721_, _16438_, _16437_);
  or (_16439_, _16001_, _26565_);
  not (_16440_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_16441_, _16001_, _16440_);
  and (_16442_, _16441_, _24069_);
  and (_16443_, _16442_, _16439_);
  nor (_16444_, _24068_, _16440_);
  or (_16445_, _16001_, _23711_);
  and (_16446_, _16441_, _24645_);
  and (_16447_, _16446_, _16445_);
  or (_16448_, _16447_, _16444_);
  or (_16449_, _16448_, _16443_);
  and (_06742_, _16449_, _22762_);
  or (_16450_, _16001_, _00451_);
  not (_16451_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_16452_, _16001_, _16451_);
  and (_16453_, _16452_, _24069_);
  and (_16454_, _16453_, _16450_);
  nor (_16456_, _24068_, _16451_);
  and (_16457_, _16008_, _24291_);
  nand (_16458_, _16457_, _23594_);
  or (_16459_, _16457_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_16460_, _16459_, _24645_);
  and (_16461_, _16460_, _16458_);
  or (_16462_, _16461_, _16456_);
  or (_16463_, _16462_, _16454_);
  and (_06744_, _16463_, _22762_);
  or (_16464_, _16001_, _00373_);
  not (_16465_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_16466_, _16001_, _16465_);
  and (_16467_, _16466_, _24069_);
  and (_16468_, _16467_, _16464_);
  nor (_16469_, _24068_, _16465_);
  and (_16470_, _16008_, _24067_);
  nand (_16471_, _16470_, _23594_);
  or (_16472_, _16470_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_16473_, _16472_, _24645_);
  and (_16474_, _16473_, _16471_);
  or (_16475_, _16474_, _16469_);
  or (_16476_, _16475_, _16468_);
  and (_06745_, _16476_, _22762_);
  and (_16477_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and (_16478_, _07513_, _23649_);
  or (_06748_, _16478_, _16477_);
  or (_16479_, _16001_, _00545_);
  not (_16480_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_16481_, _16001_, _16480_);
  and (_16482_, _16481_, _24069_);
  and (_16483_, _16482_, _16479_);
  nor (_16484_, _24068_, _16480_);
  and (_16485_, _16008_, _24118_);
  nand (_16486_, _16485_, _23594_);
  or (_16487_, _16485_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_16488_, _16487_, _24645_);
  and (_16489_, _16488_, _16486_);
  or (_16490_, _16489_, _16484_);
  or (_16491_, _16490_, _16483_);
  and (_06752_, _16491_, _22762_);
  and (_16492_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  and (_16493_, _16018_, _23778_);
  or (_06754_, _16493_, _16492_);
  and (_16494_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  and (_16495_, _16277_, _24050_);
  or (_06758_, _16495_, _16494_);
  and (_16496_, _05714_, _23824_);
  and (_16497_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  or (_27159_, _16497_, _16496_);
  or (_16498_, _16001_, _00708_);
  not (_16499_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_16500_, _16001_, _16499_);
  and (_16501_, _16500_, _24069_);
  and (_16502_, _16501_, _16498_);
  nor (_16503_, _24068_, _16499_);
  and (_16504_, _16008_, _24125_);
  nand (_16505_, _16504_, _23594_);
  or (_16506_, _16504_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_16507_, _16506_, _24645_);
  and (_16508_, _16507_, _16505_);
  or (_16509_, _16508_, _16503_);
  or (_16510_, _16509_, _16502_);
  and (_06760_, _16510_, _22762_);
  or (_16511_, _16001_, _00620_);
  not (_16512_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_16513_, _16001_, _16512_);
  and (_16514_, _16513_, _24069_);
  and (_16515_, _16514_, _16511_);
  nor (_16516_, _24068_, _16512_);
  not (_16517_, _16008_);
  or (_16518_, _16517_, _24751_);
  and (_16519_, _16518_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_16520_, _23065_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_16521_, _16520_, _24745_);
  and (_16522_, _16521_, _16008_);
  or (_16523_, _16522_, _16519_);
  and (_16524_, _16523_, _24645_);
  or (_16525_, _16524_, _16516_);
  or (_16526_, _16525_, _16515_);
  and (_06762_, _16526_, _22762_);
  and (_16527_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  and (_16528_, _16277_, _23707_);
  or (_06765_, _16528_, _16527_);
  or (_16529_, _16001_, _00794_);
  not (_16530_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_16531_, _16001_, _16530_);
  and (_16532_, _16531_, _24069_);
  and (_16533_, _16532_, _16529_);
  nor (_16534_, _24068_, _16530_);
  and (_16535_, _16008_, _24705_);
  nand (_16536_, _16535_, _23594_);
  or (_16537_, _16535_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_16538_, _16537_, _24645_);
  and (_16539_, _16538_, _16536_);
  or (_16540_, _16539_, _16534_);
  or (_16541_, _16540_, _16533_);
  and (_06767_, _16541_, _22762_);
  and (_16542_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  and (_16543_, _16331_, _23824_);
  or (_06770_, _16543_, _16542_);
  and (_16544_, _24639_, _23778_);
  and (_16545_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_06777_, _16545_, _16544_);
  and (_16546_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and (_16547_, _16375_, _23778_);
  or (_06782_, _16547_, _16546_);
  and (_16548_, _05714_, _23898_);
  and (_16549_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  or (_06784_, _16549_, _16548_);
  and (_16550_, _01810_, _23707_);
  and (_16551_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_06787_, _16551_, _16550_);
  and (_16552_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and (_16553_, _16325_, _23707_);
  or (_06790_, _16553_, _16552_);
  and (_16554_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and (_16555_, _16375_, _23946_);
  or (_06793_, _16555_, _16554_);
  and (_16556_, _24121_, _26750_);
  nand (_16557_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_16558_, _16557_, _24127_);
  nor (_16559_, _12952_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or (_16560_, _16559_, _24154_);
  nand (_16561_, _16560_, _12956_);
  or (_16562_, _12956_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_16563_, _16562_, _16561_);
  or (_16564_, _16563_, _16558_);
  and (_16565_, _16564_, _24166_);
  or (_06794_, _16565_, _16556_);
  and (_16566_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  and (_16567_, _16319_, _23898_);
  or (_06802_, _16567_, _16566_);
  and (_16568_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  and (_16569_, _16319_, _23649_);
  or (_06812_, _16569_, _16568_);
  and (_16570_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  and (_16571_, _16371_, _23824_);
  or (_26973_, _16571_, _16570_);
  and (_16572_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and (_16573_, _16311_, _23778_);
  or (_06824_, _16573_, _16572_);
  and (_16574_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  and (_16575_, _16371_, _24050_);
  or (_06831_, _16575_, _16574_);
  and (_16576_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and (_16577_, _16311_, _23747_);
  or (_06833_, _16577_, _16576_);
  and (_16578_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  and (_16579_, _16281_, _24050_);
  or (_06837_, _16579_, _16578_);
  and (_16580_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  and (_16581_, _16281_, _23946_);
  or (_06859_, _16581_, _16580_);
  and (_16582_, _06506_, _25078_);
  not (_16583_, _16582_);
  and (_16584_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and (_16585_, _16582_, _24050_);
  or (_06864_, _16585_, _16584_);
  or (_16586_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_16587_, _16586_, _22762_);
  nand (_16588_, _24078_, _23702_);
  and (_06866_, _16588_, _16587_);
  and (_16589_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  and (_16590_, _16281_, _23649_);
  or (_06869_, _16590_, _16589_);
  and (_16591_, _02200_, _23707_);
  and (_16592_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_27168_, _16592_, _16591_);
  and (_16593_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  and (_16594_, _16303_, _24050_);
  or (_06885_, _16594_, _16593_);
  and (_16595_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  and (_16596_, _16303_, _23747_);
  or (_06887_, _16596_, _16595_);
  and (_16597_, _05714_, _23649_);
  and (_16598_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  or (_06891_, _16598_, _16597_);
  and (_16599_, _06506_, _01808_);
  not (_16600_, _16599_);
  and (_16601_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  and (_16602_, _16599_, _23898_);
  or (_26987_, _16602_, _16601_);
  and (_16603_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and (_16604_, _16299_, _23707_);
  or (_06901_, _16604_, _16603_);
  and (_16605_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  and (_16606_, _16277_, _23898_);
  or (_06911_, _16606_, _16605_);
  and (_16607_, _16349_, _23898_);
  and (_16608_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  or (_06913_, _16608_, _16607_);
  and (_16609_, _05714_, _23747_);
  and (_16610_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  or (_06915_, _16610_, _16609_);
  and (_16611_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  and (_16612_, _16277_, _23778_);
  or (_06917_, _16612_, _16611_);
  and (_16613_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and (_16614_, _16289_, _23778_);
  or (_06923_, _16614_, _16613_);
  and (_16615_, _05350_, _23747_);
  and (_16616_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or (_06925_, _16616_, _16615_);
  and (_16617_, _16349_, _23747_);
  and (_16618_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or (_06926_, _16618_, _16617_);
  and (_16619_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and (_16620_, _16285_, _24050_);
  or (_06929_, _16620_, _16619_);
  and (_16621_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  and (_16622_, _16281_, _23707_);
  or (_06932_, _16622_, _16621_);
  and (_16623_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and (_16624_, _16359_, _23778_);
  or (_06938_, _16624_, _16623_);
  and (_06939_, _26682_, _22762_);
  and (_06960_, _26727_, _22762_);
  and (_16625_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_16626_, _16359_, _23946_);
  or (_06965_, _16626_, _16625_);
  and (_16627_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  and (_16628_, _16122_, _23898_);
  or (_06969_, _16628_, _16627_);
  and (_16629_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  and (_16630_, _16122_, _24050_);
  or (_06972_, _16630_, _16629_);
  and (_16631_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  and (_16632_, _15975_, _23707_);
  or (_06974_, _16632_, _16631_);
  and (_16633_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  and (_16634_, _15975_, _23649_);
  or (_26998_, _16634_, _16633_);
  and (_16635_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_16636_, _15907_, _23824_);
  or (_26999_, _16636_, _16635_);
  and (_16637_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_16638_, _15846_, _23747_);
  or (_27004_, _16638_, _16637_);
  and (_16639_, _06646_, _23649_);
  and (_16640_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_06986_, _16640_, _16639_);
  and (_16641_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_16642_, _15846_, _23778_);
  or (_06994_, _16642_, _16641_);
  and (_16643_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  and (_16644_, _14996_, _23898_);
  or (_06999_, _16644_, _16643_);
  and (_16645_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_16646_, _16285_, _23946_);
  or (_07013_, _16646_, _16645_);
  and (_16647_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and (_16648_, _13894_, _24050_);
  or (_07018_, _16648_, _16647_);
  and (_16649_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  and (_16650_, _13828_, _23946_);
  or (_07022_, _16650_, _16649_);
  and (_16651_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  and (_16652_, _16281_, _23898_);
  or (_26994_, _16652_, _16651_);
  and (_16653_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  and (_16654_, _12728_, _23747_);
  or (_07053_, _16654_, _16653_);
  and (_16655_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  and (_16656_, _06888_, _23747_);
  or (_07055_, _16656_, _16655_);
  and (_16657_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and (_16658_, _06918_, _23778_);
  or (_27015_, _16658_, _16657_);
  and (_16659_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  and (_16660_, _16281_, _23778_);
  or (_07061_, _16660_, _16659_);
  and (_16661_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and (_16662_, _16285_, _23707_);
  or (_07081_, _16662_, _16661_);
  and (_16663_, _12782_, _23747_);
  and (_16664_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_07086_, _16664_, _16663_);
  and (_16665_, _06646_, _23707_);
  and (_16666_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_07089_, _16666_, _16665_);
  and (_16667_, _06646_, _24050_);
  and (_16668_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_07092_, _16668_, _16667_);
  and (_16669_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and (_16670_, _16289_, _23946_);
  or (_07098_, _16670_, _16669_);
  and (_16671_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and (_16672_, _16289_, _23707_);
  or (_07106_, _16672_, _16671_);
  and (_16673_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and (_16674_, _16289_, _24050_);
  or (_07110_, _16674_, _16673_);
  and (_16675_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and (_16676_, _16285_, _23747_);
  or (_07150_, _16676_, _16675_);
  and (_16677_, _06755_, _23707_);
  and (_16678_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_27158_, _16678_, _16677_);
  and (_16679_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and (_16680_, _16285_, _23824_);
  or (_07173_, _16680_, _16679_);
  and (_16681_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and (_16682_, _16285_, _23898_);
  or (_26993_, _16682_, _16681_);
  and (_16683_, _06755_, _24050_);
  and (_16684_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_07191_, _16684_, _16683_);
  and (_16685_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and (_16686_, _16285_, _23778_);
  or (_07195_, _16686_, _16685_);
  and (_16687_, _10347_, _24050_);
  and (_16688_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  or (_07203_, _16688_, _16687_);
  nand (_07218_, _00077_, _22762_);
  nand (_07222_, _00112_, _22762_);
  nor (_07226_, _00029_, rst);
  nor (_07228_, _00046_, rst);
  nand (_07231_, _00147_, _22762_);
  nor (_07237_, _26788_, rst);
  nor (_07241_, _26826_, rst);
  and (_16689_, _05350_, _23649_);
  and (_16690_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  or (_07244_, _16690_, _16689_);
  and (_16691_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  and (_16692_, _16293_, _23707_);
  or (_07246_, _16692_, _16691_);
  and (_16693_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and (_16694_, _24692_, _23778_);
  or (_07250_, _16694_, _16693_);
  and (_16695_, _06646_, _23898_);
  and (_16696_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_07253_, _16696_, _16695_);
  and (_16697_, _06646_, _23778_);
  and (_16698_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_07278_, _16698_, _16697_);
  and (_16699_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and (_16700_, _01967_, _23778_);
  or (_07282_, _16700_, _16699_);
  and (_16701_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and (_16702_, _16289_, _23898_);
  or (_07287_, _16702_, _16701_);
  and (_16703_, _15850_, _24050_);
  and (_16704_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  or (_07290_, _16704_, _16703_);
  nand (_16705_, _25644_, _24598_);
  or (_26862_[2], _16705_, _04996_);
  and (_16706_, _25649_, _23898_);
  and (_16707_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_07300_, _16707_, _16706_);
  and (_16708_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and (_16709_, _16289_, _23747_);
  or (_07305_, _16709_, _16708_);
  and (_16710_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and (_16711_, _16289_, _23824_);
  or (_07310_, _16711_, _16710_);
  nor (_26885_[4], _25919_, rst);
  and (_26886_[7], _26752_, _22762_);
  and (_16712_, _06755_, _23824_);
  and (_16713_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_07338_, _16713_, _16712_);
  and (_16714_, _23946_, _23833_);
  and (_16715_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_07342_, _16715_, _16714_);
  and (_26884_, _26777_, _22762_);
  and (_16716_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  and (_16717_, _16293_, _23747_);
  or (_26989_, _16717_, _16716_);
  and (_16718_, _06755_, _23898_);
  and (_16719_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_07359_, _16719_, _16718_);
  and (_16720_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and (_16721_, _16293_, _23824_);
  or (_07363_, _16721_, _16720_);
  and (_16722_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and (_16723_, _16293_, _23898_);
  or (_07390_, _16723_, _16722_);
  and (_16724_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  and (_16725_, _16293_, _23778_);
  or (_07396_, _16725_, _16724_);
  and (_16726_, _24699_, _24050_);
  and (_16727_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  or (_07402_, _16727_, _16726_);
  and (_16728_, _08167_, _23649_);
  and (_16729_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  or (_07408_, _16729_, _16728_);
  and (_16730_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_16731_, _06918_, _23946_);
  or (_07416_, _16731_, _16730_);
  and (_16732_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_16733_, _06918_, _23747_);
  or (_07425_, _16733_, _16732_);
  and (_16734_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  and (_16735_, _16293_, _23946_);
  or (_07428_, _16735_, _16734_);
  and (_16736_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and (_16737_, _06918_, _23824_);
  or (_27016_, _16737_, _16736_);
  and (_16738_, _06755_, _23649_);
  and (_16739_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_07435_, _16739_, _16738_);
  and (_16740_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  and (_16741_, _16293_, _23649_);
  or (_26990_, _16741_, _16740_);
  and (_16742_, _04760_, _24329_);
  not (_16743_, _16742_);
  and (_16744_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  and (_16745_, _16742_, _23946_);
  or (_07441_, _16745_, _16744_);
  and (_16746_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  and (_16747_, _16742_, _23747_);
  or (_07445_, _16747_, _16746_);
  and (_16748_, _04760_, _23752_);
  not (_16749_, _16748_);
  and (_16750_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and (_16751_, _16748_, _23649_);
  or (_07453_, _16751_, _16750_);
  and (_16752_, _04760_, _23656_);
  not (_16753_, _16752_);
  and (_16754_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  and (_16755_, _16752_, _23747_);
  or (_07481_, _16755_, _16754_);
  and (_16756_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  and (_16757_, _16599_, _23649_);
  or (_07485_, _16757_, _16756_);
  and (_16758_, _04760_, _25078_);
  not (_16759_, _16758_);
  and (_16760_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  and (_16761_, _16758_, _23747_);
  or (_07487_, _16761_, _16760_);
  and (_16762_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  and (_16763_, _16599_, _23747_);
  or (_07491_, _16763_, _16762_);
  and (_16764_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  and (_16765_, _16599_, _23824_);
  or (_07495_, _16765_, _16764_);
  and (_16766_, _04760_, _24282_);
  not (_16767_, _16766_);
  and (_16768_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and (_16769_, _16766_, _23649_);
  or (_07498_, _16769_, _16768_);
  and (_16770_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and (_16771_, _16766_, _23824_);
  or (_26951_, _16771_, _16770_);
  and (_16772_, _04760_, _23911_);
  not (_16773_, _16772_);
  and (_16774_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and (_16775_, _16772_, _23649_);
  or (_26948_, _16775_, _16774_);
  and (_16776_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  and (_16777_, _15991_, _23898_);
  or (_07507_, _16777_, _16776_);
  and (_16778_, _06651_, _23778_);
  and (_16779_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  or (_27152_, _16779_, _16778_);
  and (_16780_, _04760_, _23784_);
  not (_16781_, _16780_);
  and (_16782_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and (_16783_, _16780_, _24050_);
  or (_07520_, _16783_, _16782_);
  and (_16784_, _06511_, _23707_);
  and (_16785_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_07523_, _16785_, _16784_);
  and (_16786_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and (_16787_, _16780_, _23778_);
  or (_07529_, _16787_, _16786_);
  and (_16788_, _16022_, _24050_);
  and (_16789_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_07531_, _16789_, _16788_);
  and (_16790_, _16349_, _23946_);
  and (_16791_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or (_07532_, _16791_, _16790_);
  and (_16792_, _15850_, _23946_);
  and (_16793_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or (_07535_, _16793_, _16792_);
  and (_16794_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  and (_16795_, _16599_, _23707_);
  or (_07538_, _16795_, _16794_);
  and (_16796_, _23992_, _23946_);
  and (_16797_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_07540_, _16797_, _16796_);
  and (_16798_, _08307_, _24067_);
  nand (_16799_, _16798_, _23594_);
  or (_16800_, _16798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_16801_, _16800_, _12774_);
  and (_16802_, _16801_, _16799_);
  and (_16803_, _08313_, _23892_);
  or (_16804_, _16803_, _16802_);
  and (_07546_, _16804_, _22762_);
  and (_16805_, _08307_, _24678_);
  nand (_16806_, _16805_, _23594_);
  or (_16807_, _16805_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_16808_, _16807_, _12774_);
  and (_16809_, _16808_, _16806_);
  and (_16810_, _08313_, _24685_);
  or (_16811_, _16810_, _16809_);
  and (_07549_, _16811_, _22762_);
  and (_16812_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  and (_16813_, _16048_, _23747_);
  or (_26946_, _16813_, _16812_);
  and (_16814_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  and (_16815_, _16599_, _24050_);
  or (_07561_, _16815_, _16814_);
  and (_16816_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  and (_16817_, _16599_, _23946_);
  or (_26988_, _16817_, _16816_);
  and (_16818_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  and (_16819_, _15991_, _23946_);
  or (_07564_, _16819_, _16818_);
  and (_16820_, _08307_, _24296_);
  nand (_16821_, _16820_, _23594_);
  or (_16822_, _16820_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_16823_, _16822_, _12774_);
  and (_16824_, _16823_, _16821_);
  and (_16825_, _08313_, _23642_);
  or (_16826_, _16825_, _16824_);
  and (_07565_, _16826_, _22762_);
  and (_16827_, _16349_, _23649_);
  and (_16828_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  or (_07567_, _16828_, _16827_);
  and (_16829_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  and (_16830_, _15991_, _23707_);
  or (_07569_, _16830_, _16829_);
  not (_16831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_16832_, _01999_, _16831_);
  or (_16833_, _16832_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_16834_, _16833_, _08307_);
  nand (_16835_, _05826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_16836_, _16835_, _08307_);
  or (_16837_, _16836_, _05827_);
  and (_16838_, _16837_, _16834_);
  or (_16839_, _16838_, _08313_);
  or (_16840_, _12774_, _24043_);
  and (_16841_, _16840_, _22762_);
  and (_07571_, _16841_, _16839_);
  and (_16842_, _08307_, _24125_);
  nand (_16843_, _16842_, _23594_);
  or (_16844_, _16842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_16845_, _16844_, _12774_);
  and (_16846_, _16845_, _16843_);
  and (_16847_, _08313_, _23939_);
  or (_16848_, _16847_, _16846_);
  and (_07573_, _16848_, _22762_);
  and (_16849_, _08307_, _24118_);
  nand (_16850_, _16849_, _23594_);
  or (_16851_, _16849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_16852_, _16851_, _12774_);
  and (_16853_, _16852_, _16850_);
  and (_16854_, _08313_, _23738_);
  or (_16855_, _16854_, _16853_);
  and (_07575_, _16855_, _22762_);
  and (_16856_, _24050_, _24006_);
  and (_16857_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  or (_07579_, _16857_, _16856_);
  and (_16858_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and (_16859_, _16748_, _24050_);
  or (_26960_, _16859_, _16858_);
  and (_16860_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and (_16861_, _16748_, _23778_);
  or (_07587_, _16861_, _16860_);
  and (_16862_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_16863_, _16862_, _02041_);
  and (_16864_, _02009_, _01988_);
  or (_16865_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_16866_, _16865_, _12758_);
  or (_16867_, _16866_, _02001_);
  or (_16868_, _16867_, _16863_);
  nor (_16869_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_16870_, _16869_, _12764_);
  and (_16871_, _16870_, _16868_);
  and (_16872_, _01978_, _23892_);
  and (_16873_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_16874_, _16873_, _16872_);
  or (_16875_, _16874_, _16871_);
  and (_07593_, _16875_, _22762_);
  and (_16876_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_16877_, _16876_, _02041_);
  and (_16878_, _02009_, _01987_);
  nor (_16879_, _16878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor (_16880_, _16879_, _16864_);
  or (_16881_, _16880_, _02001_);
  or (_16882_, _16881_, _16877_);
  or (_16883_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_16884_, _16883_, _01979_);
  and (_16885_, _16884_, _16882_);
  and (_16886_, _01978_, _24685_);
  and (_16887_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_16888_, _16887_, _16886_);
  or (_16889_, _16888_, _16885_);
  and (_07596_, _16889_, _22762_);
  and (_16890_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  and (_16891_, _16752_, _23946_);
  or (_07598_, _16891_, _16890_);
  and (_16892_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  and (_16893_, _16752_, _23778_);
  or (_07602_, _16893_, _16892_);
  and (_16894_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  and (_16895_, _16758_, _23946_);
  or (_07604_, _16895_, _16894_);
  and (_16896_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  and (_16897_, _16758_, _23898_);
  or (_07607_, _16897_, _16896_);
  nor (_16898_, _02025_, _12687_);
  nand (_16899_, _16898_, _02041_);
  and (_16900_, _02009_, _01992_);
  and (_16901_, _16900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_16902_, _16900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_16903_, _16902_, _16901_);
  and (_16904_, _16903_, _02002_);
  nand (_16905_, _16904_, _16899_);
  nand (_16906_, _02001_, _12687_);
  and (_16907_, _16906_, _01979_);
  and (_16908_, _16907_, _16905_);
  and (_16909_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_16910_, _16909_, _16908_);
  and (_16911_, _01978_, _23642_);
  or (_16912_, _16911_, _16910_);
  and (_07609_, _16912_, _22762_);
  and (_16913_, _06651_, _23747_);
  and (_16914_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  or (_07611_, _16914_, _16913_);
  and (_16915_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and (_16916_, _16766_, _24050_);
  or (_07614_, _16916_, _16915_);
  and (_16917_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and (_16918_, _16299_, _24050_);
  or (_07617_, _16918_, _16917_);
  nor (_16919_, _02018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_16920_, _16919_, _02019_);
  not (_16921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_16922_, _02025_, _16921_);
  nand (_16923_, _16922_, _02041_);
  and (_16924_, _16923_, _02002_);
  nand (_16925_, _16924_, _16920_);
  nand (_16926_, _02001_, _16921_);
  and (_16927_, _16926_, _01979_);
  and (_16928_, _16927_, _16925_);
  and (_16929_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_16930_, _16929_, _16928_);
  and (_16931_, _01978_, _24043_);
  or (_16932_, _16931_, _16930_);
  and (_07620_, _16932_, _22762_);
  and (_16933_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_16934_, _16901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_16935_, _16934_, _02018_);
  and (_16936_, _02026_, _02009_);
  and (_16937_, _16936_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_16938_, _16937_, _01996_);
  or (_16939_, _16938_, _02001_);
  or (_16940_, _16939_, _16935_);
  or (_16941_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_16942_, _16941_, _01979_);
  and (_16943_, _16942_, _16940_);
  or (_16944_, _16943_, _16933_);
  and (_16945_, _01978_, _23939_);
  or (_16946_, _16945_, _16944_);
  and (_07622_, _16946_, _22762_);
  and (_16947_, _16349_, _23707_);
  and (_16948_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  or (_07625_, _16948_, _16947_);
  and (_16949_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and (_16950_, _16772_, _23898_);
  or (_07627_, _16950_, _16949_);
  not (_16951_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_16952_, _02025_, _16951_);
  nand (_16953_, _16952_, _02041_);
  and (_16954_, _02009_, _01990_);
  nor (_16955_, _16954_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_16956_, _16955_, _16900_);
  and (_16957_, _16956_, _02002_);
  nand (_16958_, _16957_, _16953_);
  and (_16959_, _02001_, _16951_);
  nor (_16960_, _16959_, _12764_);
  and (_16961_, _16960_, _16958_);
  and (_16962_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_16963_, _16962_, _16961_);
  and (_16964_, _01978_, _23738_);
  or (_16965_, _16964_, _16963_);
  and (_07630_, _16965_, _22762_);
  and (_16966_, _06651_, _23824_);
  and (_16967_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  or (_07633_, _16967_, _16966_);
  and (_16968_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and (_16969_, _16780_, _23747_);
  or (_07635_, _16969_, _16968_);
  and (_16970_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and (_16971_, _16299_, _23946_);
  or (_07638_, _16971_, _16970_);
  and (_16972_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and (_16973_, _16299_, _23649_);
  or (_07640_, _16973_, _16972_);
  and (_16974_, _16349_, _23824_);
  and (_16975_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  or (_07644_, _16975_, _16974_);
  and (_16976_, _01977_, _23738_);
  and (_16977_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_16978_, _16977_, _02041_);
  and (_16979_, _02009_, _01982_);
  or (_16980_, _16979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_16981_, _16980_, _12742_);
  or (_16982_, _16981_, _02001_);
  or (_16983_, _16982_, _16978_);
  or (_16984_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_16985_, _16984_, _01979_);
  and (_16986_, _16985_, _16983_);
  and (_16987_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_16988_, _16987_, _16986_);
  or (_16989_, _16988_, _16976_);
  and (_07646_, _16989_, _22762_);
  and (_16990_, _01977_, _23816_);
  and (_16991_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_16992_, _16991_, _02041_);
  not (_16993_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand (_16994_, _02009_, _01981_);
  and (_16995_, _16994_, _16993_);
  nor (_16996_, _16995_, _16979_);
  or (_16997_, _16996_, _02001_);
  or (_16998_, _16997_, _16992_);
  or (_16999_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_17000_, _16999_, _01979_);
  and (_17001_, _17000_, _16998_);
  and (_17002_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_17003_, _17002_, _17001_);
  or (_17004_, _17003_, _16990_);
  and (_07651_, _17004_, _22762_);
  and (_17005_, _23992_, _23707_);
  and (_17006_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_07654_, _17006_, _17005_);
  and (_17007_, _02001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_17008_, _12708_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_17009_, _16994_, _02002_);
  and (_17010_, _17009_, _17008_);
  or (_17011_, _17010_, _17007_);
  or (_17012_, _17011_, _01977_);
  and (_17013_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_17014_, _17013_, _16936_);
  and (_17015_, _17014_, _01996_);
  or (_17016_, _17015_, _17012_);
  or (_17017_, _02017_, _23892_);
  and (_17018_, _17017_, _17016_);
  or (_17019_, _17018_, _01978_);
  not (_17020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand (_17021_, _01978_, _17020_);
  and (_17022_, _17021_, _22762_);
  and (_07656_, _17022_, _17019_);
  and (_17023_, _06651_, _23898_);
  and (_17024_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  or (_07658_, _17024_, _17023_);
  and (_17025_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  and (_17026_, _16048_, _23946_);
  or (_07680_, _17026_, _17025_);
  and (_17027_, _12782_, _23707_);
  and (_17028_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_07688_, _17028_, _17027_);
  and (_17029_, _24086_, _23649_);
  and (_17030_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_07690_, _17030_, _17029_);
  and (_17031_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  and (_17032_, _16599_, _23778_);
  or (_07694_, _17032_, _17031_);
  and (_17033_, _01977_, _24043_);
  and (_17034_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_17035_, _17034_, _02041_);
  and (_17036_, _02009_, _01985_);
  nor (_17037_, _17036_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_17038_, _17037_, _02043_);
  or (_17039_, _17038_, _02001_);
  or (_17040_, _17039_, _17035_);
  or (_17041_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_17042_, _17041_, _01979_);
  and (_17043_, _17042_, _17040_);
  and (_17044_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_17045_, _17044_, _17043_);
  or (_17046_, _17045_, _17033_);
  and (_07697_, _17046_, _22762_);
  and (_17047_, _01977_, _23939_);
  and (_17048_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_17049_, _17048_, _02041_);
  and (_17050_, _02009_, _01984_);
  nor (_17051_, _17050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_17052_, _17051_, _17036_);
  or (_17053_, _17052_, _02001_);
  or (_17054_, _17053_, _17049_);
  or (_17055_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_17056_, _17055_, _01979_);
  and (_17057_, _17056_, _17054_);
  and (_17058_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_17059_, _17058_, _17057_);
  or (_17060_, _17059_, _17047_);
  and (_07699_, _17060_, _22762_);
  and (_17061_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and (_17062_, _16772_, _23946_);
  or (_07702_, _17062_, _17061_);
  nor (_26861_[2], _24574_, rst);
  and (_17063_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  and (_17064_, _15991_, _23824_);
  or (_07705_, _17064_, _17063_);
  and (_17065_, _02345_, _24050_);
  and (_17066_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_07708_, _17066_, _17065_);
  and (_17067_, _16349_, _24050_);
  and (_17068_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  or (_07712_, _17068_, _17067_);
  or (_17069_, _12675_, _24043_);
  nor (_17070_, _02078_, _16921_);
  and (_17071_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_17072_, _17071_, _17070_);
  or (_17073_, _17072_, _02073_);
  and (_17074_, _17073_, _22762_);
  and (_07716_, _17074_, _17069_);
  and (_17075_, _06511_, _23824_);
  and (_17076_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_07719_, _17076_, _17075_);
  and (_17077_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  and (_17078_, _16752_, _23898_);
  or (_07724_, _17078_, _17077_);
  and (_17079_, _06511_, _23898_);
  and (_17080_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_07729_, _17080_, _17079_);
  and (_17081_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  and (_17082_, _16048_, _24050_);
  or (_26947_, _17082_, _17081_);
  and (_17083_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and (_17084_, _16299_, _23778_);
  or (_07739_, _17084_, _17083_);
  and (_17085_, _05281_, _23898_);
  and (_17086_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_07741_, _17086_, _17085_);
  and (_17087_, _01810_, _23824_);
  and (_17088_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_07744_, _17088_, _17087_);
  and (_17089_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and (_17090_, _13763_, _23946_);
  or (_07746_, _17090_, _17089_);
  and (_17091_, _24201_, _23986_);
  not (_17092_, _17091_);
  and (_17093_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and (_17094_, _17091_, _23707_);
  or (_07750_, _17094_, _17093_);
  and (_17095_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  and (_17096_, _17091_, _23898_);
  or (_07752_, _17096_, _17095_);
  and (_17097_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  and (_17098_, _16303_, _23707_);
  or (_07765_, _17098_, _17097_);
  nor (_17099_, _02078_, _16951_);
  and (_17100_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_17101_, _17100_, _17099_);
  and (_17102_, _17101_, _12675_);
  and (_17103_, _02073_, _23738_);
  or (_17104_, _17103_, _17102_);
  and (_07767_, _17104_, _22762_);
  or (_17105_, _12675_, _23816_);
  nor (_17106_, _02078_, _12754_);
  and (_17107_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_17108_, _17107_, _17106_);
  or (_17109_, _17108_, _02073_);
  and (_17110_, _17109_, _22762_);
  and (_07769_, _17110_, _17105_);
  and (_17111_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  and (_17112_, _02306_, _23747_);
  or (_07771_, _17112_, _17111_);
  or (_17113_, _12675_, _23892_);
  and (_17114_, _17113_, _22762_);
  and (_17115_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_17116_, _02079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_17117_, _17116_, _17115_);
  or (_17118_, _17117_, _02073_);
  and (_07773_, _17118_, _17114_);
  and (_17119_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and (_17120_, _07492_, _23707_);
  or (_07775_, _17120_, _17119_);
  and (_17121_, _06511_, _23747_);
  and (_17122_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_07777_, _17122_, _17121_);
  or (_17123_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_17124_, _02079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_17125_, _17124_, _17123_);
  or (_17126_, _17125_, _02073_);
  nand (_17127_, _02073_, _23772_);
  and (_17128_, _17127_, _22762_);
  and (_07779_, _17128_, _17126_);
  and (_17129_, _06511_, _23946_);
  and (_17130_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_07781_, _17130_, _17129_);
  and (_17131_, _06511_, _23649_);
  and (_17132_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_07797_, _17132_, _17131_);
  and (_17133_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and (_17134_, _02298_, _23898_);
  or (_07800_, _17134_, _17133_);
  or (_17135_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_17136_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_17137_, _17136_, _17135_);
  or (_17138_, _17137_, _02077_);
  nand (_17139_, _02077_, _23772_);
  and (_17140_, _17139_, _17138_);
  or (_17141_, _17140_, _02073_);
  or (_17142_, _12675_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_17143_, _17142_, _22762_);
  and (_07802_, _17143_, _17141_);
  and (_17144_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  and (_17145_, _24692_, _23824_);
  or (_07805_, _17145_, _17144_);
  and (_17146_, _05350_, _23824_);
  and (_17147_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  or (_07818_, _17147_, _17146_);
  and (_17148_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  and (_17149_, _01967_, _23747_);
  or (_07820_, _17149_, _17148_);
  and (_17150_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and (_17151_, _16299_, _23824_);
  or (_07823_, _17151_, _17150_);
  or (_17152_, _12671_, _24043_);
  and (_17153_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_17154_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_17155_, _17154_, _17153_);
  or (_17156_, _17155_, _02077_);
  and (_17157_, _17156_, _12675_);
  and (_17158_, _17157_, _17152_);
  and (_17159_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_17160_, _17159_, _17158_);
  and (_07828_, _17160_, _22762_);
  or (_17161_, _12671_, _23939_);
  and (_17162_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_17163_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_17164_, _17163_, _17162_);
  or (_17165_, _17164_, _02077_);
  and (_17166_, _17165_, _12675_);
  and (_17167_, _17166_, _17161_);
  and (_17168_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_17169_, _17168_, _17167_);
  and (_07830_, _17169_, _22762_);
  or (_17170_, _12671_, _23642_);
  and (_17171_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_17172_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_17173_, _17172_, _17171_);
  or (_17174_, _17173_, _02077_);
  and (_17175_, _17174_, _12675_);
  and (_17176_, _17175_, _17170_);
  and (_17177_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_17178_, _17177_, _17176_);
  and (_07832_, _17178_, _22762_);
  or (_17179_, _12671_, _23738_);
  and (_17180_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_17181_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_17182_, _17181_, _17180_);
  or (_17183_, _17182_, _02077_);
  and (_17184_, _17183_, _12675_);
  and (_17185_, _17184_, _17179_);
  and (_17186_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_17187_, _17186_, _17185_);
  and (_07834_, _17187_, _22762_);
  or (_17188_, _12671_, _23816_);
  and (_17189_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_17190_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_17191_, _17190_, _17189_);
  or (_17192_, _17191_, _02077_);
  and (_17193_, _17192_, _12675_);
  and (_17194_, _17193_, _17188_);
  and (_17195_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_17196_, _17195_, _17194_);
  and (_07838_, _17196_, _22762_);
  and (_17197_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and (_17198_, _16299_, _23898_);
  or (_07851_, _17198_, _17197_);
  and (_17199_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  and (_17200_, _08351_, _23898_);
  or (_07854_, _17200_, _17199_);
  and (_17201_, _24331_, _23824_);
  and (_17202_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_08089_, _17202_, _17201_);
  and (_17203_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  and (_17204_, _15895_, _23747_);
  or (_08090_, _17204_, _17203_);
  and (_17205_, _06517_, _23649_);
  and (_17206_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_08092_, _17206_, _17205_);
  and (_17207_, _24275_, _23076_);
  and (_17208_, _17207_, _23824_);
  not (_17209_, _17207_);
  and (_17210_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_08094_, _17210_, _17208_);
  and (_17211_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and (_17212_, _16303_, _23824_);
  or (_08100_, _17212_, _17211_);
  and (_17213_, _06517_, _23747_);
  and (_17214_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_08103_, _17214_, _17213_);
  and (_17215_, _23903_, _23076_);
  and (_17216_, _17215_, _23946_);
  not (_17217_, _17215_);
  and (_17218_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  or (_08107_, _17218_, _17216_);
  and (_17219_, _25733_, _23707_);
  and (_17220_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_08110_, _17220_, _17219_);
  and (_17221_, _24085_, _23076_);
  and (_17222_, _17221_, _23649_);
  not (_17223_, _17221_);
  and (_17224_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_08115_, _17224_, _17222_);
  and (_17225_, _06517_, _23707_);
  and (_17226_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_08118_, _17226_, _17225_);
  and (_17227_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and (_17228_, _16780_, _23898_);
  or (_08162_, _17228_, _17227_);
  and (_17229_, _25078_, _23076_);
  and (_17230_, _17229_, _23707_);
  not (_17231_, _17229_);
  and (_17232_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_27207_, _17232_, _17230_);
  and (_17233_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and (_17234_, _16780_, _23824_);
  or (_08170_, _17234_, _17233_);
  and (_17235_, _16022_, _23707_);
  and (_17236_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_27195_, _17236_, _17235_);
  and (_17237_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and (_17238_, _16780_, _23649_);
  or (_08172_, _17238_, _17237_);
  and (_17239_, _05119_, _23898_);
  and (_17240_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  or (_08175_, _17240_, _17239_);
  and (_17241_, _02345_, _23649_);
  and (_17242_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_08179_, _17242_, _17241_);
  and (_17243_, _24699_, _23707_);
  and (_17244_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  or (_08181_, _17244_, _17243_);
  and (_17245_, _24283_, _23649_);
  and (_17246_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or (_08183_, _17246_, _17245_);
  and (_17247_, _25649_, _23824_);
  and (_17248_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_08188_, _17248_, _17247_);
  and (_17249_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  and (_17250_, _24222_, _23747_);
  or (_08190_, _17250_, _17249_);
  and (_17251_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  and (_17252_, _05193_, _24050_);
  or (_08195_, _17252_, _17251_);
  and (_17253_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and (_17254_, _16780_, _23946_);
  or (_26945_, _17254_, _17253_);
  and (_17255_, _23784_, _23076_);
  not (_17256_, _17255_);
  and (_17257_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and (_17258_, _17255_, _23778_);
  or (_08202_, _17258_, _17257_);
  and (_17259_, _24371_, _24050_);
  and (_17260_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_08203_, _17260_, _17259_);
  and (_17261_, _16022_, _23747_);
  and (_17262_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_08205_, _17262_, _17261_);
  and (_17263_, _24370_, _23986_);
  and (_17264_, _17263_, _23824_);
  not (_17265_, _17263_);
  and (_17266_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or (_08208_, _17266_, _17264_);
  and (_17268_, _25656_, _23778_);
  and (_17269_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_08210_, _17269_, _17268_);
  and (_17270_, _04922_, _23747_);
  and (_17271_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  or (_08215_, _17271_, _17270_);
  and (_17272_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  and (_17273_, _16303_, _23946_);
  or (_08421_, _17273_, _17272_);
  and (_17274_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  and (_17275_, _16303_, _23649_);
  or (_08424_, _17275_, _17274_);
  and (_17276_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  and (_17277_, _02298_, _23824_);
  or (_08427_, _17277_, _17276_);
  and (_17278_, _06517_, _24050_);
  and (_17279_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_08429_, _17279_, _17278_);
  and (_17280_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  and (_17281_, _15895_, _23649_);
  or (_08432_, _17281_, _17280_);
  and (_17282_, _17215_, _24050_);
  and (_17283_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or (_08435_, _17283_, _17282_);
  and (_17284_, _15850_, _23898_);
  and (_17285_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or (_08439_, _17285_, _17284_);
  and (_17286_, _05119_, _23824_);
  and (_17287_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  or (_08442_, _17287_, _17286_);
  and (_17288_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_17289_, _16307_, _23946_);
  or (_08449_, _17289_, _17288_);
  and (_17290_, _24283_, _23946_);
  and (_17291_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or (_08451_, _17291_, _17290_);
  and (_17292_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and (_17293_, _16307_, _23649_);
  or (_08454_, _17293_, _17292_);
  and (_17295_, _06524_, _23707_);
  and (_17296_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  or (_08458_, _17296_, _17295_);
  and (_17297_, _06524_, _24050_);
  and (_17298_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  or (_08463_, _17298_, _17297_);
  and (_17299_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  and (_17300_, _24222_, _23649_);
  or (_27246_, _17300_, _17299_);
  and (_17301_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  and (_17302_, _15895_, _23946_);
  or (_08476_, _17302_, _17301_);
  and (_17303_, _02374_, _23898_);
  and (_17304_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or (_08487_, _17304_, _17303_);
  or (_17305_, _06686_, _03323_);
  or (_17306_, _17305_, _06726_);
  or (_17307_, _04938_, _24608_);
  or (_17308_, _03274_, _26626_);
  or (_17309_, _17308_, _17307_);
  or (_17310_, _17309_, _04244_);
  or (_17311_, _17310_, _17306_);
  or (_17312_, _17311_, _03320_);
  and (_17313_, _17312_, _22768_);
  and (_17314_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_17315_, _17314_, _03336_);
  or (_17316_, _17315_, _17313_);
  and (_26873_, _17316_, _22762_);
  and (_17317_, _25618_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_17318_, _24613_, _24606_);
  or (_17319_, _17318_, _26635_);
  or (_17320_, _17319_, _06719_);
  or (_17321_, _05079_, _25633_);
  or (_17322_, _05065_, _05088_);
  or (_17323_, _17322_, _17321_);
  or (_17324_, _17323_, _17320_);
  and (_17325_, _17324_, _25644_);
  or (_26870_[1], _17325_, _17317_);
  and (_17326_, _25618_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_17327_, _03275_, _26641_);
  or (_17328_, _17327_, _12858_);
  or (_17329_, _17328_, _26653_);
  or (_17330_, _17329_, _02255_);
  or (_17331_, _04962_, _02263_);
  or (_17332_, _06686_, _06079_);
  or (_17333_, _17332_, _17331_);
  or (_17334_, _17333_, _06576_);
  or (_17335_, _17334_, _17330_);
  or (_17336_, _17335_, _06696_);
  and (_17337_, _17336_, _25644_);
  or (_26871_[3], _17337_, _17326_);
  and (_17338_, _02370_, _23747_);
  and (_17339_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_08522_, _17339_, _17338_);
  or (_17340_, _03331_, _26572_);
  or (_17341_, _03330_, _25636_);
  and (_17342_, _17341_, _22766_);
  and (_17343_, _17342_, _17340_);
  and (_17344_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_17345_, _17344_, _05003_);
  or (_17346_, _17345_, _17343_);
  and (_26869_[2], _17346_, _22762_);
  or (_17347_, _06870_, _04945_);
  and (_17348_, _17347_, _22768_);
  and (_17349_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_17350_, _17349_, _24570_);
  or (_17351_, _17350_, _17348_);
  and (_26872_[1], _17351_, _22762_);
  and (_17352_, _02370_, _23649_);
  and (_17353_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_08526_, _17353_, _17352_);
  and (_17354_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  and (_17355_, _07492_, _23898_);
  or (_08538_, _17355_, _17354_);
  and (_17356_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and (_17357_, _07492_, _23824_);
  or (_27240_, _17357_, _17356_);
  and (_17358_, _17263_, _23778_);
  and (_17359_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or (_27193_, _17359_, _17358_);
  and (_17360_, _05281_, _23707_);
  and (_17361_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_08740_, _17361_, _17360_);
  and (_17362_, _25656_, _24050_);
  and (_17363_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_08749_, _17363_, _17362_);
  and (_17364_, _25656_, _23707_);
  and (_17365_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_08765_, _17365_, _17364_);
  and (_17366_, _02370_, _23778_);
  and (_17367_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_08771_, _17367_, _17366_);
  and (_17368_, _05281_, _24050_);
  and (_17369_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_08773_, _17369_, _17368_);
  and (_17370_, _25739_, _23778_);
  and (_17371_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or (_27068_, _17371_, _17370_);
  and (_17372_, _25739_, _23898_);
  and (_17373_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  or (_08826_, _17373_, _17372_);
  and (_17374_, _25739_, _23824_);
  and (_17375_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  or (_08828_, _17375_, _17374_);
  and (_17376_, _06524_, _23946_);
  and (_17377_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  or (_08882_, _17377_, _17376_);
  and (_17378_, _23991_, _23789_);
  and (_17379_, _17378_, _23778_);
  not (_17380_, _17378_);
  and (_17381_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or (_27289_, _17381_, _17379_);
  and (_17382_, _17263_, _23747_);
  and (_17383_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or (_08909_, _17383_, _17382_);
  and (_17384_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  and (_17385_, _07492_, _23747_);
  or (_08931_, _17385_, _17384_);
  and (_17386_, _12782_, _24050_);
  and (_17387_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_08939_, _17387_, _17386_);
  and (_17388_, _23656_, _23076_);
  and (_17389_, _17388_, _24050_);
  not (_17390_, _17388_);
  and (_17391_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_08943_, _17391_, _17389_);
  and (_17392_, _04922_, _23946_);
  and (_17393_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or (_08947_, _17393_, _17392_);
  and (_17394_, _04922_, _23649_);
  and (_17395_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  or (_08951_, _17395_, _17394_);
  and (_17396_, _23903_, _23789_);
  and (_17397_, _17396_, _23649_);
  not (_17398_, _17396_);
  and (_17399_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or (_08959_, _17399_, _17397_);
  and (_17400_, _17396_, _23898_);
  and (_17401_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  or (_08963_, _17401_, _17400_);
  and (_17402_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and (_17403_, _16780_, _23707_);
  or (_08965_, _17403_, _17402_);
  and (_17404_, _24005_, _23789_);
  and (_17405_, _17404_, _23649_);
  not (_17406_, _17404_);
  and (_17407_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_08969_, _17407_, _17405_);
  and (_17408_, _17404_, _23824_);
  and (_17409_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_08971_, _17409_, _17408_);
  and (_17410_, _23986_, _23789_);
  and (_17411_, _17410_, _23946_);
  not (_17412_, _17410_);
  and (_17413_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_08975_, _17413_, _17411_);
  and (_17414_, _17410_, _23747_);
  and (_17415_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_08977_, _17415_, _17414_);
  and (_17416_, _23789_, _23069_);
  and (_17418_, _17416_, _23946_);
  not (_17419_, _17416_);
  and (_17420_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or (_08981_, _17420_, _17418_);
  and (_17421_, _17416_, _23747_);
  and (_17422_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  or (_08983_, _17422_, _17421_);
  and (_17423_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and (_17424_, _16307_, _23707_);
  or (_26986_, _17424_, _17423_);
  and (_17425_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and (_17426_, _16307_, _24050_);
  or (_08988_, _17426_, _17425_);
  and (_17427_, _17388_, _23946_);
  and (_17428_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_08995_, _17428_, _17427_);
  and (_17429_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  and (_17430_, _15895_, _23898_);
  or (_09002_, _17430_, _17429_);
  and (_17431_, _01808_, _23789_);
  and (_17432_, _17431_, _24050_);
  not (_17433_, _17431_);
  and (_17434_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or (_09010_, _17434_, _17432_);
  and (_17435_, _17431_, _23649_);
  and (_17436_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  or (_09011_, _17436_, _17435_);
  and (_17437_, _17431_, _23898_);
  and (_17438_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  or (_09014_, _17438_, _17437_);
  and (_17439_, _24329_, _23789_);
  and (_17440_, _17439_, _23707_);
  not (_17441_, _17439_);
  and (_17442_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_09018_, _17442_, _17440_);
  and (_17443_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  and (_17444_, _15991_, _23778_);
  or (_09022_, _17444_, _17443_);
  and (_17445_, _17439_, _23747_);
  and (_17446_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_09025_, _17446_, _17445_);
  and (_17447_, _25078_, _23789_);
  and (_17448_, _17447_, _23707_);
  not (_17449_, _17447_);
  and (_17450_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_09035_, _17450_, _17448_);
  and (_17451_, _06517_, _23778_);
  and (_17452_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_09038_, _17452_, _17451_);
  and (_17453_, _06517_, _23898_);
  and (_17454_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_27150_, _17454_, _17453_);
  and (_17455_, _14956_, _24050_);
  and (_17456_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_09047_, _17456_, _17455_);
  and (_17457_, _14956_, _23946_);
  and (_17458_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_09049_, _17458_, _17457_);
  and (_17459_, _15850_, _23778_);
  and (_17460_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  or (_27209_, _17460_, _17459_);
  and (_17461_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  and (_17462_, _15895_, _23824_);
  or (_09059_, _17462_, _17461_);
  and (_17463_, _12733_, _23747_);
  and (_17464_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or (_09061_, _17464_, _17463_);
  and (_17465_, _17447_, _23778_);
  and (_17466_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_09071_, _17466_, _17465_);
  and (_17467_, _24282_, _23789_);
  and (_17468_, _17467_, _23707_);
  not (_17469_, _17467_);
  and (_17470_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  or (_09074_, _17470_, _17468_);
  and (_17471_, _17467_, _23946_);
  and (_17472_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or (_09075_, _17472_, _17471_);
  and (_17473_, _17467_, _23898_);
  and (_17474_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  or (_09079_, _17474_, _17473_);
  and (_17475_, _23789_, _23752_);
  and (_17476_, _17475_, _23946_);
  not (_17477_, _17475_);
  and (_17478_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or (_09086_, _17478_, _17476_);
  and (_17479_, _23789_, _23656_);
  and (_17480_, _17479_, _24050_);
  not (_17481_, _17479_);
  and (_17482_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_27273_, _17482_, _17480_);
  and (_17483_, _17378_, _23824_);
  and (_17484_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or (_09094_, _17484_, _17483_);
  and (_17485_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and (_17486_, _16307_, _23778_);
  or (_26985_, _17486_, _17485_);
  and (_17487_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and (_17488_, _16582_, _23707_);
  or (_09101_, _17488_, _17487_);
  and (_17489_, _17404_, _24050_);
  and (_17490_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_09110_, _17490_, _17489_);
  and (_17491_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  and (_17492_, _16048_, _23707_);
  or (_09112_, _17492_, _17491_);
  and (_17493_, _17410_, _23707_);
  and (_17494_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_09114_, _17494_, _17493_);
  and (_17495_, _17416_, _23707_);
  and (_17496_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or (_09118_, _17496_, _17495_);
  and (_17497_, _02370_, _24050_);
  and (_17498_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_09140_, _17498_, _17497_);
  and (_17499_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and (_17500_, _16772_, _23778_);
  or (_09167_, _17500_, _17499_);
  and (_17501_, _17479_, _23824_);
  and (_17502_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_09172_, _17502_, _17501_);
  and (_17503_, _17447_, _23649_);
  and (_17504_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_09174_, _17504_, _17503_);
  and (_17505_, _17475_, _23707_);
  and (_17506_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or (_09179_, _17506_, _17505_);
  and (_17507_, _17221_, _24050_);
  and (_17508_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_09184_, _17508_, _17507_);
  and (_17509_, _06524_, _23778_);
  and (_17510_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  or (_09191_, _17510_, _17509_);
  and (_17511_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and (_17512_, _16307_, _23824_);
  or (_09194_, _17512_, _17511_);
  and (_17513_, _10347_, _23898_);
  and (_17514_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or (_27125_, _17514_, _17513_);
  and (_17515_, _17396_, _23946_);
  and (_17516_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or (_09202_, _17516_, _17515_);
  and (_17517_, _17416_, _23778_);
  and (_17518_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  or (_09206_, _17518_, _17517_);
  and (_17519_, _17447_, _23898_);
  and (_17520_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_09215_, _17520_, _17519_);
  and (_17521_, _17475_, _23898_);
  and (_17522_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or (_09219_, _17522_, _17521_);
  and (_17523_, _06530_, _23707_);
  and (_17524_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  or (_09225_, _17524_, _17523_);
  and (_17525_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and (_17526_, _16307_, _23898_);
  or (_09228_, _17526_, _17525_);
  and (_17527_, _17388_, _23778_);
  and (_17528_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_09254_, _17528_, _17527_);
  and (_17529_, _12782_, _23898_);
  and (_17530_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_27076_, _17530_, _17529_);
  and (_17531_, _12782_, _23778_);
  and (_17532_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_09258_, _17532_, _17531_);
  and (_17533_, _17410_, _23778_);
  and (_17534_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_09270_, _17534_, _17533_);
  and (_17535_, _23906_, _23069_);
  and (_17536_, _17535_, _23946_);
  not (_17537_, _17535_);
  and (_17538_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_09274_, _17538_, _17536_);
  and (_17539_, _01808_, _23906_);
  and (_17540_, _17539_, _23707_);
  not (_17541_, _17539_);
  and (_17542_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_26933_, _17542_, _17540_);
  and (_17543_, _17539_, _23824_);
  and (_17544_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_09282_, _17544_, _17543_);
  and (_17545_, _06530_, _24050_);
  and (_17546_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  or (_27148_, _17546_, _17545_);
  and (_17547_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and (_17548_, _16772_, _23824_);
  or (_09291_, _17548_, _17547_);
  and (_17549_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and (_17550_, _16582_, _23824_);
  or (_09296_, _17550_, _17549_);
  and (_17551_, _23906_, _23752_);
  and (_17552_, _17551_, _23707_);
  not (_17553_, _17551_);
  and (_17554_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_09299_, _17554_, _17552_);
  and (_17555_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_17556_, _17555_, _26154_);
  and (_17557_, _17555_, _26154_);
  or (_17558_, _17557_, _17556_);
  and (_09302_, _17558_, _22762_);
  and (_17559_, _17551_, _23649_);
  and (_17560_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_09305_, _17560_, _17559_);
  and (_17561_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and (_17562_, _16582_, _23898_);
  or (_09309_, _17562_, _17561_);
  and (_09312_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _22762_);
  and (_09315_, _00845_, _22762_);
  and (_09317_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _22762_);
  or (_17563_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_17564_, _17555_, rst);
  and (_09321_, _17564_, _17563_);
  and (_17565_, _05042_, _23946_);
  and (_17566_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_09327_, _17566_, _17565_);
  and (_17567_, _12733_, _23824_);
  and (_17568_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  or (_09331_, _17568_, _17567_);
  and (_17569_, _23906_, _23656_);
  and (_17570_, _17569_, _23946_);
  not (_17571_, _17569_);
  and (_17572_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or (_09334_, _17572_, _17570_);
  and (_17573_, _17569_, _23778_);
  and (_17574_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or (_09340_, _17574_, _17573_);
  and (_17575_, _25078_, _23906_);
  and (_17576_, _17575_, _24050_);
  not (_17577_, _17575_);
  and (_17578_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  or (_09343_, _17578_, _17576_);
  and (_17579_, _17575_, _23898_);
  and (_17580_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or (_09347_, _17580_, _17579_);
  and (_17581_, _24282_, _23906_);
  and (_17582_, _17581_, _23707_);
  not (_17583_, _17581_);
  and (_17584_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_09350_, _17584_, _17582_);
  and (_17585_, _17581_, _23824_);
  and (_17586_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_09354_, _17586_, _17585_);
  and (_17587_, _24010_, _23906_);
  and (_17588_, _17587_, _23946_);
  not (_17589_, _17587_);
  and (_17590_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  or (_09357_, _17590_, _17588_);
  and (_17591_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  and (_17592_, _08477_, _23747_);
  or (_09359_, _17592_, _17591_);
  and (_17593_, _24085_, _23906_);
  and (_17594_, _17593_, _23946_);
  not (_17595_, _17593_);
  and (_17596_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or (_09366_, _17596_, _17594_);
  and (_17597_, _17593_, _23824_);
  and (_17598_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  or (_09368_, _17598_, _17597_);
  and (_17599_, _23906_, _23784_);
  and (_17601_, _17599_, _23707_);
  not (_17602_, _17599_);
  and (_17603_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_09370_, _17603_, _17601_);
  and (_17604_, _17599_, _23649_);
  and (_17605_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_09373_, _17605_, _17604_);
  and (_17606_, _17599_, _23778_);
  and (_17607_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_09375_, _17607_, _17606_);
  and (_17608_, _23911_, _23906_);
  and (_17609_, _17608_, _24050_);
  not (_17610_, _17608_);
  and (_17611_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_09379_, _17611_, _17609_);
  and (_17612_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and (_17613_, _16582_, _23778_);
  or (_09382_, _17613_, _17612_);
  and (_17614_, _17608_, _23649_);
  and (_17615_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_09384_, _17615_, _17614_);
  and (_17616_, _06524_, _23747_);
  and (_17617_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  or (_09387_, _17617_, _17616_);
  and (_17618_, _05350_, _24050_);
  and (_17619_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or (_09421_, _17619_, _17618_);
  and (_17620_, _05119_, _23707_);
  and (_17621_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or (_09523_, _17621_, _17620_);
  and (_17622_, _25618_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_17623_, _02256_, _02273_);
  or (_17624_, _17623_, _06686_);
  or (_17625_, _06697_, _03273_);
  or (_17626_, _17625_, _17624_);
  or (_17627_, _17626_, _06696_);
  and (_17628_, _17627_, _25644_);
  or (_26867_[1], _17628_, _17622_);
  and (_17629_, _17388_, _23747_);
  and (_17630_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_09600_, _17630_, _17629_);
  and (_17631_, _17388_, _23824_);
  and (_17632_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_09612_, _17632_, _17631_);
  and (_17633_, _14956_, _23898_);
  and (_17634_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_09626_, _17634_, _17633_);
  and (_17635_, _07536_, _23824_);
  and (_17636_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  or (_09638_, _17636_, _17635_);
  and (_17637_, _14956_, _23778_);
  and (_17638_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or (_09652_, _17638_, _17637_);
  and (_17639_, _17229_, _23747_);
  and (_17640_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_09668_, _17640_, _17639_);
  and (_17641_, _05281_, _23778_);
  and (_17642_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_09681_, _17642_, _17641_);
  and (_17643_, _17229_, _23824_);
  and (_17644_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_27206_, _17644_, _17643_);
  and (_17645_, _14956_, _23747_);
  and (_17646_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_09731_, _17646_, _17645_);
  and (_17647_, _17229_, _24050_);
  and (_17648_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_09733_, _17648_, _17647_);
  and (_17649_, _14956_, _23824_);
  and (_17650_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_09737_, _17650_, _17649_);
  and (_17651_, _17229_, _23946_);
  and (_17652_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_09753_, _17652_, _17651_);
  or (_17653_, _04891_, _24043_);
  or (_17654_, _05165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_17655_, _05166_, _26098_);
  and (_17656_, _17655_, _17654_);
  and (_17657_, _07418_, _24310_);
  or (_17658_, _17657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_17659_, _05144_, _04860_);
  and (_17660_, _17659_, _17658_);
  or (_17661_, _05151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_17662_, _05152_);
  and (_17663_, _17662_, _24302_);
  and (_17664_, _17663_, _17661_);
  and (_17665_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_17666_, _17665_, _17664_);
  or (_17667_, _17666_, _17660_);
  or (_17668_, _17667_, _17656_);
  or (_17669_, _17668_, _24299_);
  and (_17670_, _17669_, _24294_);
  and (_17671_, _17670_, _17653_);
  and (_17672_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_17673_, _17672_, _17671_);
  and (_09769_, _17673_, _22762_);
  and (_17674_, _12786_, _23747_);
  and (_17675_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or (_09818_, _17675_, _17674_);
  and (_17676_, _24283_, _23707_);
  and (_17677_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or (_09821_, _17677_, _17676_);
  and (_17678_, _09913_, _23778_);
  and (_17679_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_09823_, _17679_, _17678_);
  and (_17680_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  and (_17681_, _08477_, _23824_);
  or (_09837_, _17681_, _17680_);
  and (_17682_, _12786_, _23824_);
  and (_17683_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  or (_09839_, _17683_, _17682_);
  and (_17684_, _24283_, _24050_);
  and (_17685_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  or (_09854_, _17685_, _17684_);
  and (_17686_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and (_17687_, _01967_, _23824_);
  or (_09860_, _17687_, _17686_);
  and (_17688_, _12786_, _23898_);
  and (_17689_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  or (_27075_, _17689_, _17688_);
  and (_17690_, _25649_, _24050_);
  and (_17691_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_09887_, _17691_, _17690_);
  and (_17692_, _17207_, _23946_);
  and (_17693_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_09900_, _17693_, _17692_);
  and (_17694_, _17207_, _23649_);
  and (_17695_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_09906_, _17695_, _17694_);
  and (_17696_, _17207_, _23747_);
  and (_17697_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_09919_, _17697_, _17696_);
  and (_17698_, _24652_, _24064_);
  nand (_17699_, _17698_, _24118_);
  and (_17700_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_17701_, _25170_, _24117_);
  and (_17702_, _17701_, _24064_);
  and (_17703_, _17702_, _24068_);
  and (_17704_, _17703_, _22948_);
  and (_17705_, _17704_, _00708_);
  or (_17706_, _17705_, _17700_);
  or (_17707_, _17706_, _06343_);
  not (_17708_, _06343_);
  or (_17709_, _17708_, _01255_);
  and (_17710_, _17709_, _22762_);
  and (_09940_, _17710_, _17707_);
  and (_17711_, _17535_, _23824_);
  and (_17712_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_09945_, _17712_, _17711_);
  and (_17713_, _17539_, _23649_);
  and (_17714_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_09950_, _17714_, _17713_);
  and (_17715_, _06524_, _23824_);
  and (_17716_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  or (_09952_, _17716_, _17715_);
  and (_17717_, _17539_, _23778_);
  and (_17718_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_09954_, _17718_, _17717_);
  and (_17719_, _24329_, _23906_);
  and (_17720_, _17719_, _23747_);
  not (_17721_, _17719_);
  and (_17722_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or (_09956_, _17722_, _17720_);
  and (_17723_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_17724_, _17704_, _00875_);
  or (_17725_, _17724_, _17723_);
  or (_17726_, _17725_, _06343_);
  or (_17727_, _17708_, _04299_);
  and (_17728_, _17727_, _22762_);
  and (_09964_, _17728_, _17726_);
  and (_17729_, _17719_, _23778_);
  and (_17730_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  or (_09966_, _17730_, _17729_);
  and (_17731_, _06524_, _23898_);
  and (_17732_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  or (_27149_, _17732_, _17731_);
  and (_17733_, _17551_, _23898_);
  and (_17734_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_09974_, _17734_, _17733_);
  and (_17735_, _17698_, _24291_);
  nor (_17736_, _17735_, _06343_);
  or (_17737_, _17736_, _26565_);
  not (_17738_, _17736_);
  or (_17739_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_17740_, _17739_, _22762_);
  and (_09976_, _17740_, _17737_);
  and (_17741_, _17569_, _23824_);
  and (_17742_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or (_09988_, _17742_, _17741_);
  and (_17743_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and (_17744_, _16582_, _23946_);
  or (_09991_, _17744_, _17743_);
  and (_17745_, _17575_, _23747_);
  and (_17746_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  or (_26918_, _17746_, _17745_);
  or (_17747_, _17736_, _00545_);
  or (_17748_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_17749_, _17748_, _22762_);
  and (_10005_, _17749_, _17747_);
  and (_17750_, _17581_, _23649_);
  and (_17751_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_10007_, _17751_, _17750_);
  and (_17752_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  and (_17753_, _05199_, _23707_);
  or (_10013_, _17753_, _17752_);
  and (_17754_, _15012_, _23898_);
  and (_17755_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_10021_, _17755_, _17754_);
  and (_17756_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and (_17757_, _16582_, _23649_);
  or (_10036_, _17757_, _17756_);
  and (_17758_, _05838_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_17759_, _17758_, _05839_);
  and (_17760_, _17759_, _00276_);
  or (_17761_, _00277_, _00276_);
  nor (_17762_, _17761_, _23594_);
  and (_17763_, _00280_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_17764_, _17763_, _25773_);
  or (_17765_, _17764_, _17762_);
  or (_17766_, _17765_, _17760_);
  nand (_17767_, _25777_, _23702_);
  and (_17768_, _17767_, _22762_);
  and (_10039_, _17768_, _17766_);
  nand (_17769_, _17738_, _00793_);
  or (_17770_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_17771_, _17770_, _22762_);
  and (_10048_, _17771_, _17769_);
  or (_17772_, _17736_, _00451_);
  or (_17773_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_17774_, _17773_, _22762_);
  and (_10050_, _17774_, _17772_);
  and (_17775_, _01808_, _24201_);
  not (_17776_, _17775_);
  and (_17777_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  and (_17778_, _17775_, _23778_);
  or (_10055_, _17778_, _17777_);
  and (_17779_, _17535_, _24050_);
  and (_17780_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_26934_, _17780_, _17779_);
  and (_17781_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_17782_, _17704_, _00620_);
  or (_17783_, _17782_, _17781_);
  or (_17784_, _17783_, _06343_);
  or (_17785_, _17708_, _01192_);
  and (_17786_, _17785_, _22762_);
  and (_10074_, _17786_, _17784_);
  and (_17787_, _17551_, _23946_);
  and (_17788_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_10083_, _17788_, _17787_);
  and (_17789_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_17790_, _17704_, _00545_);
  or (_17791_, _17790_, _17789_);
  or (_17792_, _17791_, _06343_);
  nand (_17793_, _06343_, _01129_);
  and (_17794_, _17793_, _22762_);
  and (_10085_, _17794_, _17792_);
  and (_17795_, _17569_, _24050_);
  and (_17796_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or (_26921_, _17796_, _17795_);
  and (_17797_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and (_17798_, _16772_, _23747_);
  or (_10089_, _17798_, _17797_);
  and (_17799_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_17800_, _17704_, _00451_);
  or (_17801_, _17800_, _17799_);
  or (_17802_, _17801_, _06343_);
  nand (_17803_, _06343_, _01061_);
  and (_17804_, _17803_, _22762_);
  and (_10097_, _17804_, _17802_);
  and (_17805_, _17593_, _23747_);
  and (_17806_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  or (_10100_, _17806_, _17805_);
  and (_17807_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and (_17808_, _16582_, _23747_);
  or (_10104_, _17808_, _17807_);
  and (_17809_, _17581_, _23778_);
  and (_17810_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_10108_, _17810_, _17809_);
  and (_17811_, _17608_, _23898_);
  and (_17812_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_10110_, _17812_, _17811_);
  and (_17813_, _17575_, _23707_);
  and (_17814_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or (_10114_, _17814_, _17813_);
  and (_17815_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and (_17816_, _16772_, _24050_);
  or (_26949_, _17816_, _17815_);
  nand (_17817_, _17738_, _00372_);
  or (_17818_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_17819_, _17818_, _22762_);
  and (_10125_, _17819_, _17817_);
  or (_17820_, _17736_, _00708_);
  or (_17821_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_17822_, _17821_, _22762_);
  and (_10128_, _17822_, _17820_);
  or (_17823_, _17736_, _00620_);
  or (_17824_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_17825_, _17824_, _22762_);
  and (_10130_, _17825_, _17823_);
  nor (_17826_, _17699_, _00372_);
  and (_17827_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_17828_, _17827_, _06343_);
  or (_17829_, _17828_, _17826_);
  nand (_17830_, _06343_, _00993_);
  and (_17831_, _17830_, _22762_);
  and (_10132_, _17831_, _17829_);
  and (_17832_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_17833_, _17704_, _26565_);
  or (_17834_, _17833_, _17832_);
  or (_17835_, _17834_, _06343_);
  or (_17836_, _17708_, _00930_);
  and (_17837_, _17836_, _22762_);
  and (_10133_, _17837_, _17835_);
  or (_17838_, _17736_, _00875_);
  or (_17839_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_17840_, _17839_, _22762_);
  and (_10143_, _17840_, _17838_);
  and (_17841_, _06530_, _23824_);
  and (_17842_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  or (_10147_, _17842_, _17841_);
  and (_17843_, _17608_, _23778_);
  and (_17844_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_27300_, _17844_, _17843_);
  and (_17845_, _17475_, _23778_);
  and (_17846_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  or (_10157_, _17846_, _17845_);
  and (_17847_, _25649_, _23707_);
  and (_17848_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_10163_, _17848_, _17847_);
  and (_17849_, _25649_, _23946_);
  and (_17850_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_10165_, _17850_, _17849_);
  nor (_17851_, _17699_, _00793_);
  and (_17852_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_17853_, _17852_, _06343_);
  or (_17854_, _17853_, _17851_);
  nand (_17855_, _06343_, _01318_);
  and (_17856_, _17855_, _22762_);
  and (_10169_, _17856_, _17854_);
  and (_17857_, _17587_, _24050_);
  and (_17858_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  or (_10172_, _17858_, _17857_);
  and (_26861_[1], _26676_, _22762_);
  and (_17859_, _17221_, _23707_);
  and (_17860_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_27202_, _17860_, _17859_);
  and (_17861_, _06530_, _23747_);
  and (_17862_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  or (_27146_, _17862_, _17861_);
  and (_17863_, _17479_, _23946_);
  and (_17864_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_10179_, _17864_, _17863_);
  and (_17865_, _17221_, _23946_);
  and (_17866_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_10182_, _17866_, _17865_);
  and (_17867_, _17587_, _23707_);
  and (_17868_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or (_27299_, _17868_, _17867_);
  and (_17869_, _17479_, _23707_);
  and (_17870_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_27274_, _17870_, _17869_);
  and (_17871_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and (_17872_, _16772_, _23707_);
  or (_10188_, _17872_, _17871_);
  and (_17873_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and (_17874_, _16766_, _23778_);
  or (_10192_, _17874_, _17873_);
  and (_17875_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  and (_17876_, _10331_, _23649_);
  or (_10194_, _17876_, _17875_);
  and (_17877_, _25649_, _23778_);
  and (_17878_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_10196_, _17878_, _17877_);
  and (_17879_, _17608_, _23824_);
  and (_17880_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_10197_, _17880_, _17879_);
  and (_17881_, _17475_, _23824_);
  and (_17882_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or (_10201_, _17882_, _17881_);
  and (_17883_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  and (_17884_, _10331_, _23747_);
  or (_26983_, _17884_, _17883_);
  and (_17885_, _04922_, _23707_);
  and (_17886_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  or (_10206_, _17886_, _17885_);
  and (_17887_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and (_17888_, _16766_, _23898_);
  or (_26950_, _17888_, _17887_);
  and (_17889_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and (_17890_, _16766_, _23747_);
  or (_10221_, _17890_, _17889_);
  and (_17891_, _17475_, _23747_);
  and (_17892_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or (_10225_, _17892_, _17891_);
  and (_17893_, _24852_, _24050_);
  and (_17894_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or (_10227_, _17894_, _17893_);
  and (_17895_, _17608_, _23747_);
  and (_17896_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_10231_, _17896_, _17895_);
  and (_17897_, _24283_, _23778_);
  and (_17898_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  or (_10239_, _17898_, _17897_);
  and (_17899_, _17608_, _23946_);
  and (_17900_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_10240_, _17900_, _17899_);
  and (_17901_, _17475_, _23649_);
  and (_17902_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  or (_10253_, _17902_, _17901_);
  and (_17903_, _17608_, _23707_);
  and (_17904_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_10258_, _17904_, _17903_);
  and (_17905_, _17475_, _24050_);
  and (_17906_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  or (_10260_, _17906_, _17905_);
  and (_17907_, _24050_, _23912_);
  and (_17908_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or (_27268_, _17908_, _17907_);
  and (_17909_, _24699_, _23747_);
  and (_17910_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  or (_27190_, _17910_, _17909_);
  and (_17911_, _24699_, _23898_);
  and (_17912_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  or (_10280_, _17912_, _17911_);
  and (_17913_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  and (_17914_, _10331_, _23946_);
  or (_26984_, _17914_, _17913_);
  and (_17915_, _17599_, _23898_);
  and (_17916_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_10287_, _17916_, _17915_);
  and (_17917_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  and (_17918_, _10331_, _23707_);
  or (_10289_, _17918_, _17917_);
  and (_17919_, _23912_, _23707_);
  and (_17920_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or (_10293_, _17920_, _17919_);
  and (_17921_, _24699_, _23946_);
  and (_17922_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or (_10297_, _17922_, _17921_);
  and (_17923_, _17599_, _23824_);
  and (_17924_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_10301_, _17924_, _17923_);
  and (_17925_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  and (_17926_, _10331_, _24050_);
  or (_10304_, _17926_, _17925_);
  and (_17927_, _17467_, _23778_);
  and (_17928_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or (_10308_, _17928_, _17927_);
  and (_17929_, _02345_, _23898_);
  and (_17930_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_10310_, _17930_, _17929_);
  and (_17931_, _17467_, _23824_);
  and (_17932_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or (_10314_, _17932_, _17931_);
  and (_17933_, _00276_, _24296_);
  nand (_17934_, _17933_, _23594_);
  not (_17935_, _25777_);
  or (_17936_, _17933_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_17937_, _17936_, _17935_);
  and (_17938_, _17937_, _17934_);
  or (_17939_, _17938_, _25918_);
  and (_10317_, _17939_, _22762_);
  and (_17940_, _17599_, _23747_);
  and (_17941_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_27295_, _17941_, _17940_);
  and (_17942_, _06530_, _23649_);
  and (_17943_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  or (_27147_, _17943_, _17942_);
  and (_17944_, _00276_, _24118_);
  or (_17945_, _17944_, _25775_);
  nand (_17946_, _17944_, _23594_);
  and (_17947_, _17946_, _17945_);
  or (_17948_, _17947_, _25779_);
  and (_10329_, _17948_, _22762_);
  and (_17949_, _00276_, _24125_);
  nand (_17950_, _17949_, _23594_);
  or (_17951_, _17949_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_17952_, _17951_, _17935_);
  and (_17953_, _17952_, _17950_);
  and (_17954_, _25777_, _23939_);
  or (_17955_, _17954_, _17953_);
  and (_10330_, _17955_, _22762_);
  and (_17956_, _17599_, _23946_);
  and (_17957_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_27296_, _17957_, _17956_);
  and (_17958_, _17467_, _23747_);
  and (_17959_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or (_27269_, _17959_, _17958_);
  and (_17960_, _25656_, _23747_);
  and (_17961_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_10336_, _17961_, _17960_);
  or (_17962_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_17963_, _00334_, _26541_);
  or (_17964_, _17963_, _00428_);
  or (_17965_, _17964_, _00511_);
  or (_17966_, _17965_, _00600_);
  or (_17967_, _17966_, _00679_);
  and (_17968_, _17967_, _23596_);
  and (_17969_, _23471_, _23143_);
  not (_17970_, _23471_);
  and (_17971_, _23473_, _17970_);
  or (_17972_, _17971_, _17969_);
  and (_17973_, _17972_, _23087_);
  nand (_17974_, _23516_, _23482_);
  or (_17975_, _23516_, _23145_);
  and (_17976_, _17975_, _23480_);
  and (_17977_, _17976_, _17974_);
  and (_17978_, _23599_, _23214_);
  and (_17979_, _17978_, _23418_);
  and (_17980_, _01112_, _26152_);
  and (_17982_, _17980_, _01233_);
  nand (_17983_, _17982_, _17979_);
  nand (_17984_, _17983_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_17985_, _17984_, _17977_);
  nor (_17986_, _17985_, _17973_);
  nand (_17987_, _17986_, _00767_);
  or (_17988_, _17987_, _17968_);
  or (_17989_, _17988_, _00852_);
  and (_17990_, _17989_, _17962_);
  or (_17991_, _17990_, _00276_);
  and (_17992_, _04388_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_17993_, _17992_, _04389_);
  nand (_17994_, _17993_, _00276_);
  and (_17995_, _17994_, _17991_);
  or (_17996_, _17995_, _25777_);
  or (_17997_, _17935_, _23816_);
  and (_17998_, _17997_, _22762_);
  and (_10338_, _17998_, _17996_);
  and (_17999_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and (_18000_, _23501_, _23480_);
  and (_18001_, _23467_, _23087_);
  or (_18002_, _18001_, _18000_);
  and (_18003_, _18002_, _17999_);
  not (_18004_, _17999_);
  or (_18005_, _18004_, _23579_);
  and (_18006_, _18005_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_18007_, _18006_, _00276_);
  or (_18008_, _18007_, _18003_);
  or (_18009_, _24705_, _00527_);
  nand (_18010_, _18009_, _00276_);
  or (_18011_, _18010_, _05827_);
  and (_18012_, _18011_, _18008_);
  or (_18013_, _18012_, _25777_);
  or (_18014_, _17935_, _24043_);
  and (_18015_, _18014_, _22762_);
  and (_10341_, _18015_, _18013_);
  and (_18016_, _17263_, _23898_);
  and (_18017_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or (_10342_, _18017_, _18016_);
  and (_18018_, _17599_, _24050_);
  and (_18019_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_10345_, _18019_, _18018_);
  and (_18020_, _17467_, _23649_);
  and (_18021_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or (_10346_, _18021_, _18020_);
  and (_18022_, _17593_, _23778_);
  and (_18023_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or (_10349_, _18023_, _18022_);
  and (_10353_, _05850_, _22762_);
  and (_18024_, _17263_, _23946_);
  and (_18025_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or (_10355_, _18025_, _18024_);
  and (_26861_[0], _24632_, _22762_);
  and (_18026_, _17467_, _24050_);
  and (_18027_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  or (_27270_, _18027_, _18026_);
  and (_18028_, _17207_, _24050_);
  and (_18029_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_10360_, _18029_, _18028_);
  and (_18030_, _00276_, _24067_);
  nand (_18031_, _18030_, _23594_);
  or (_18032_, _18030_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_18033_, _18032_, _17935_);
  and (_18034_, _18033_, _18031_);
  and (_18035_, _25777_, _23892_);
  or (_18036_, _18035_, _18034_);
  and (_10364_, _18036_, _22762_);
  and (_18037_, _17263_, _23649_);
  and (_18038_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  or (_27194_, _18038_, _18037_);
  and (_18039_, _17593_, _23898_);
  and (_18040_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or (_10368_, _18040_, _18039_);
  and (_18041_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and (_18042_, _16311_, _23824_);
  or (_10370_, _18042_, _18041_);
  and (_18043_, _17447_, _23824_);
  and (_18044_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_10375_, _18044_, _18043_);
  and (_18045_, _05119_, _24050_);
  and (_18046_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  or (_10377_, _18046_, _18045_);
  and (_18047_, _17593_, _23649_);
  and (_18048_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or (_10379_, _18048_, _18047_);
  and (_18049_, _15856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  or (_18050_, _24315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_18051_, _18050_, _26118_);
  nor (_18052_, _18051_, _26097_);
  nor (_18053_, _18052_, _05168_);
  or (_18054_, _18053_, _18049_);
  and (_18055_, _18054_, _22762_);
  nor (_18056_, _24299_, _24293_);
  and (_10382_, _18056_, _18055_);
  or (_18057_, _12675_, _23939_);
  and (_18058_, _02079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_18059_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_18060_, _18059_, _18058_);
  or (_18061_, _18060_, _02073_);
  and (_18062_, _18061_, _22762_);
  and (_10384_, _18062_, _18057_);
  and (_18063_, _17593_, _24050_);
  and (_18064_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or (_27297_, _18064_, _18063_);
  and (_18065_, _16022_, _23824_);
  and (_18066_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_10390_, _18066_, _18065_);
  and (_18067_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and (_18068_, _16311_, _23898_);
  or (_26976_, _18068_, _18067_);
  and (_18069_, _17447_, _23747_);
  and (_18070_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_10395_, _18070_, _18069_);
  and (_18071_, _06544_, _24050_);
  and (_18072_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_10397_, _18072_, _18071_);
  and (_18073_, _16022_, _23778_);
  and (_18074_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_10399_, _18074_, _18073_);
  and (_18075_, _17447_, _23946_);
  and (_18076_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_10401_, _18076_, _18075_);
  and (_18077_, _17593_, _23707_);
  and (_18078_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or (_10403_, _18078_, _18077_);
  and (_18079_, _16022_, _23946_);
  and (_18080_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_10406_, _18080_, _18079_);
  and (_18081_, _24371_, _23946_);
  and (_18082_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_27198_, _18082_, _18081_);
  and (_18083_, _17587_, _23778_);
  and (_18084_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  or (_27298_, _18084_, _18083_);
  and (_18085_, _17447_, _24050_);
  and (_18086_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_10413_, _18086_, _18085_);
  and (_18087_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and (_18088_, _16311_, _23946_);
  or (_26977_, _18088_, _18087_);
  and (_18089_, _24371_, _23824_);
  and (_18090_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_10416_, _18090_, _18089_);
  nor (_10431_, _05836_, rst);
  and (_18091_, _17479_, _23778_);
  and (_18092_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_10436_, _18092_, _18091_);
  and (_18093_, _25142_, _23747_);
  and (_18094_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or (_10452_, _18094_, _18093_);
  and (_18095_, _17587_, _23898_);
  and (_18096_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  or (_10454_, _18096_, _18095_);
  and (_10471_, _05752_, _22762_);
  and (_10500_, _05764_, _22762_);
  and (_18097_, _17587_, _23824_);
  and (_18098_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or (_10511_, _18098_, _18097_);
  and (_10516_, _05820_, _22762_);
  and (_18099_, _17479_, _23898_);
  and (_18100_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_27271_, _18100_, _18099_);
  and (_10550_, _05808_, _22762_);
  and (_18101_, _17479_, _23747_);
  and (_18102_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_10559_, _18102_, _18101_);
  and (_18103_, _17587_, _23747_);
  and (_18104_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or (_10569_, _18104_, _18103_);
  and (_18105_, _04797_, _23707_);
  and (_18106_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_10574_, _18106_, _18105_);
  and (_18107_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and (_18108_, _16311_, _23649_);
  or (_10599_, _18108_, _18107_);
  and (_18109_, _17479_, _23649_);
  and (_18110_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_27272_, _18110_, _18109_);
  and (_18111_, _15012_, _23747_);
  and (_18112_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_10606_, _18112_, _18111_);
  and (_18113_, _06530_, _23778_);
  and (_18114_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  or (_10623_, _18114_, _18113_);
  and (_18115_, _17587_, _23649_);
  and (_18116_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  or (_10625_, _18116_, _18115_);
  nor (_10641_, _05791_, rst);
  and (_18117_, _17221_, _23778_);
  and (_18118_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_10646_, _18118_, _18117_);
  and (_18119_, _17439_, _23778_);
  and (_18120_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_27275_, _18120_, _18119_);
  and (_18121_, _17229_, _23898_);
  and (_18122_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_10650_, _18122_, _18121_);
  and (_10657_, _05778_, _22762_);
  and (_18123_, _17581_, _23898_);
  and (_18124_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_10660_, _18124_, _18123_);
  and (_18125_, _17581_, _23747_);
  and (_18126_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_10677_, _18126_, _18125_);
  and (_18127_, _17439_, _23898_);
  and (_18128_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_10679_, _18128_, _18127_);
  and (_18129_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  and (_18130_, _16371_, _23649_);
  or (_10701_, _18130_, _18129_);
  and (_18131_, _17229_, _23649_);
  and (_18132_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_10706_, _18132_, _18131_);
  and (_18133_, _17581_, _23946_);
  and (_18134_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_26916_, _18134_, _18133_);
  and (_18135_, _12786_, _24050_);
  and (_18136_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  or (_10710_, _18136_, _18135_);
  and (_18137_, _17388_, _23649_);
  and (_18138_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_27208_, _18138_, _18137_);
  and (_18139_, _17439_, _23824_);
  and (_18140_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_27276_, _18140_, _18139_);
  and (_18141_, _17388_, _23898_);
  and (_18142_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_10731_, _18142_, _18141_);
  and (_18143_, _17439_, _23649_);
  and (_18144_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_10735_, _18144_, _18143_);
  and (_18145_, _16022_, _23898_);
  and (_18146_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_10737_, _18146_, _18145_);
  and (_18147_, _17581_, _24050_);
  and (_18148_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_10742_, _18148_, _18147_);
  and (_18149_, _17388_, _23707_);
  and (_18150_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_10745_, _18150_, _18149_);
  and (_18151_, _17229_, _23778_);
  and (_18152_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_10748_, _18152_, _18151_);
  and (_18153_, _17439_, _23946_);
  and (_18154_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_10750_, _18154_, _18153_);
  and (_18155_, _15850_, _23707_);
  and (_18156_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or (_10755_, _18156_, _18155_);
  and (_18157_, _17575_, _23778_);
  and (_18158_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  or (_26917_, _18158_, _18157_);
  and (_18159_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  and (_18160_, _16371_, _23946_);
  or (_26974_, _18160_, _18159_);
  and (_18161_, _02345_, _23747_);
  and (_18162_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_10770_, _18162_, _18161_);
  and (_18163_, _17575_, _23824_);
  and (_18164_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  or (_10775_, _18164_, _18163_);
  and (_18165_, _08043_, _23946_);
  and (_18166_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_10780_, _18166_, _18165_);
  and (_18167_, _23991_, _23076_);
  and (_18168_, _18167_, _24050_);
  not (_18169_, _18167_);
  and (_18170_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  or (_10784_, _18170_, _18168_);
  nor (_18171_, _14782_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_18172_, _18171_, _26115_);
  and (_18173_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_18174_, _18173_, _26118_);
  nor (_18175_, _18174_, _18172_);
  nor (_18176_, _18175_, _24299_);
  and (_18177_, _24299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_18178_, _18177_, _18176_);
  and (_18179_, _18178_, _24294_);
  and (_18180_, _24293_, _23642_);
  or (_18181_, _18180_, _18179_);
  and (_10788_, _18181_, _22762_);
  and (_18182_, _17439_, _24050_);
  and (_18183_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_10791_, _18183_, _18182_);
  and (_18184_, _08043_, _23824_);
  and (_18185_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_10797_, _18185_, _18184_);
  and (_18186_, _18167_, _23707_);
  and (_18187_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or (_10799_, _18187_, _18186_);
  and (_18189_, _15012_, _23649_);
  and (_18190_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_27084_, _18190_, _18189_);
  and (_18191_, _17575_, _23649_);
  and (_18192_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or (_26919_, _18192_, _18191_);
  and (_18193_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and (_18194_, _16766_, _23946_);
  or (_10806_, _18194_, _18193_);
  and (_18195_, _12786_, _23946_);
  and (_18196_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or (_10810_, _18196_, _18195_);
  and (_18197_, _23778_, _23077_);
  and (_18198_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  or (_10813_, _18198_, _18197_);
  and (_18199_, _17575_, _23946_);
  and (_18200_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or (_10826_, _18200_, _18199_);
  and (_18201_, _17431_, _23778_);
  and (_18202_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or (_10830_, _18202_, _18201_);
  and (_18203_, _05410_, _23946_);
  and (_18204_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  or (_10832_, _18204_, _18203_);
  and (_18205_, _17431_, _23824_);
  and (_18206_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or (_10834_, _18206_, _18205_);
  and (_18207_, _25733_, _23778_);
  and (_18208_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_10838_, _18208_, _18207_);
  and (_18209_, _17569_, _23898_);
  and (_18210_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  or (_10844_, _18210_, _18209_);
  and (_18211_, _02326_, _23824_);
  and (_18212_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_10856_, _18212_, _18211_);
  and (_18213_, _17431_, _23747_);
  and (_18214_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or (_10864_, _18214_, _18213_);
  and (_18215_, _17569_, _23747_);
  and (_18216_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or (_26920_, _18216_, _18215_);
  and (_18217_, _24005_, _23076_);
  and (_18218_, _18217_, _24050_);
  not (_18219_, _18217_);
  and (_18220_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_27216_, _18220_, _18218_);
  and (_18221_, _17431_, _23946_);
  and (_18222_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or (_27277_, _18222_, _18221_);
  or (_18223_, _24294_, _24043_);
  and (_18224_, _26115_, _26098_);
  nand (_18225_, _18224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_18226_, _18225_, _24299_);
  and (_18227_, _18226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand (_18228_, _17665_, _26118_);
  or (_18229_, _18225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_18230_, _18229_, _18228_);
  nor (_18231_, _18230_, _24299_);
  or (_18232_, _18231_, _24293_);
  or (_18233_, _18232_, _18227_);
  and (_18234_, _18233_, _22762_);
  and (_10873_, _18234_, _18223_);
  and (_18235_, _17431_, _23707_);
  and (_18236_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  or (_10876_, _18236_, _18235_);
  and (_18237_, _17569_, _23649_);
  and (_18238_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  or (_10880_, _18238_, _18237_);
  and (_18239_, _17569_, _23707_);
  and (_18240_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  or (_10886_, _18240_, _18239_);
  and (_18241_, _24050_, _23755_);
  and (_18242_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or (_10888_, _18242_, _18241_);
  and (_18243_, _17416_, _23898_);
  and (_18244_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or (_10892_, _18244_, _18243_);
  and (_18245_, _17207_, _23898_);
  and (_18246_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_10895_, _18246_, _18245_);
  and (_18247_, _18167_, _23946_);
  and (_18248_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or (_10897_, _18248_, _18247_);
  and (_18249_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and (_18250_, _16766_, _23707_);
  or (_10902_, _18250_, _18249_);
  and (_18251_, _17551_, _23778_);
  and (_18252_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_26922_, _18252_, _18251_);
  and (_18253_, _17416_, _23824_);
  and (_18254_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  or (_10915_, _18254_, _18253_);
  and (_18255_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  and (_18256_, _16758_, _23778_);
  or (_26952_, _18256_, _18255_);
  and (_18257_, _17207_, _23778_);
  and (_18258_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_10920_, _18258_, _18257_);
  and (_18259_, _17551_, _23824_);
  and (_18260_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_10928_, _18260_, _18259_);
  and (_18261_, _15004_, _23946_);
  and (_18262_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or (_10930_, _18262_, _18261_);
  and (_18263_, _17207_, _23707_);
  and (_18264_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_10938_, _18264_, _18263_);
  and (_18265_, _25260_, _24654_);
  nand (_18266_, _18265_, _23594_);
  or (_18267_, _18265_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_18268_, _18267_, _24645_);
  and (_18269_, _18268_, _18266_);
  nand (_18270_, _25266_, _23702_);
  or (_18271_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_18272_, _18271_, _24069_);
  and (_18273_, _18272_, _18270_);
  and (_18274_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_18275_, _18274_, rst);
  or (_18276_, _18275_, _18273_);
  or (_10940_, _18276_, _18269_);
  and (_18277_, _17416_, _23649_);
  and (_18278_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or (_10945_, _18278_, _18277_);
  and (_18279_, _12786_, _23649_);
  and (_18280_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  or (_10947_, _18280_, _18279_);
  and (_18281_, _06544_, _23824_);
  and (_18282_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_10952_, _18282_, _18281_);
  and (_18283_, _17416_, _24050_);
  and (_18284_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  or (_10955_, _18284_, _18283_);
  and (_18285_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  and (_18286_, _16758_, _23824_);
  or (_10958_, _18286_, _18285_);
  and (_18287_, _17551_, _23747_);
  and (_18288_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_10960_, _18288_, _18287_);
  and (_18289_, _15004_, _23649_);
  and (_18290_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_27083_, _18290_, _18289_);
  and (_18291_, _07536_, _23649_);
  and (_18292_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  or (_10966_, _18292_, _18291_);
  and (_18293_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  and (_18294_, _16758_, _23649_);
  or (_10968_, _18294_, _18293_);
  and (_18295_, _17410_, _23898_);
  and (_18296_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_10973_, _18296_, _18295_);
  and (_18297_, _15004_, _23747_);
  and (_18298_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_10975_, _18298_, _18297_);
  and (_18299_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  and (_18300_, _12829_, _23747_);
  or (_10980_, _18300_, _18299_);
  and (_18301_, _06544_, _23898_);
  and (_18302_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_10982_, _18302_, _18301_);
  and (_18304_, _17551_, _24050_);
  and (_18305_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_26923_, _18305_, _18304_);
  and (_18306_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and (_18307_, _12829_, _23778_);
  or (_27223_, _18307_, _18306_);
  and (_18308_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  and (_18309_, _16758_, _24050_);
  or (_26953_, _18309_, _18308_);
  and (_18310_, _17410_, _23824_);
  and (_18311_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_27279_, _18311_, _18310_);
  and (_18312_, _17719_, _23898_);
  and (_18313_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  or (_26924_, _18313_, _18312_);
  and (_18314_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and (_18315_, _08351_, _23707_);
  or (_27226_, _18315_, _18314_);
  and (_18316_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  and (_18317_, _16758_, _23707_);
  or (_26954_, _18317_, _18316_);
  and (_18318_, _17410_, _23649_);
  and (_18319_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_27280_, _18319_, _18318_);
  and (_18320_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and (_18321_, _08351_, _23649_);
  or (_27225_, _18321_, _18320_);
  and (_18322_, _17410_, _24050_);
  and (_18323_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_27281_, _18323_, _18322_);
  and (_18324_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  and (_18325_, _05193_, _23946_);
  or (_27229_, _18325_, _18324_);
  and (_18326_, _17719_, _23824_);
  and (_18327_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or (_26925_, _18327_, _18326_);
  and (_18328_, _17215_, _23707_);
  and (_18329_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  or (_27218_, _18329_, _18328_);
  and (_18330_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  and (_18331_, _05193_, _23824_);
  or (_27227_, _18331_, _18330_);
  and (_18332_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  and (_18333_, _16371_, _23707_);
  or (_26975_, _18333_, _18332_);
  and (_18334_, _17719_, _23649_);
  and (_18335_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  or (_26926_, _18335_, _18334_);
  and (_18336_, _17404_, _23778_);
  and (_18337_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_27282_, _18337_, _18336_);
  and (_18338_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  and (_18339_, _05199_, _23946_);
  or (_27231_, _18339_, _18338_);
  and (_18340_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  and (_18341_, _16752_, _23824_);
  or (_26955_, _18341_, _18340_);
  and (_18342_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  and (_18343_, _16752_, _23649_);
  or (_26956_, _18343_, _18342_);
  and (_18344_, _18167_, _23898_);
  and (_18345_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  or (_27220_, _18345_, _18344_);
  and (_18346_, _17719_, _23946_);
  and (_18347_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or (_26927_, _18347_, _18346_);
  and (_18348_, _17404_, _23898_);
  and (_18349_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_27283_, _18349_, _18348_);
  and (_18350_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  and (_18351_, _16752_, _24050_);
  or (_26957_, _18351_, _18350_);
  and (_18352_, _17719_, _24050_);
  and (_18353_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  or (_26928_, _18353_, _18352_);
  and (_18354_, _17404_, _23747_);
  and (_18355_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_27284_, _18355_, _18354_);
  and (_18356_, _17404_, _23946_);
  and (_18357_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_27285_, _18357_, _18356_);
  and (_18358_, _17719_, _23707_);
  and (_18359_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or (_26929_, _18359_, _18358_);
  and (_18360_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  and (_18361_, _16752_, _23707_);
  or (_26958_, _18361_, _18360_);
  and (_18362_, _18167_, _23778_);
  and (_18363_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or (_27219_, _18363_, _18362_);
  and (_18364_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and (_18365_, _07492_, _23778_);
  or (_27239_, _18365_, _18364_);
  and (_18366_, _06544_, _23649_);
  and (_18367_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_27145_, _18367_, _18366_);
  and (_18368_, _17539_, _23898_);
  and (_18369_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_26930_, _18369_, _18368_);
  and (_18370_, _17404_, _23707_);
  and (_18371_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_27286_, _18371_, _18370_);
  and (_18372_, _25164_, _24654_);
  nand (_18373_, _18372_, _23594_);
  or (_18374_, _18372_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_18375_, _18374_, _24645_);
  and (_18376_, _18375_, _18373_);
  nand (_18377_, _25173_, _23702_);
  or (_18378_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_18379_, _18378_, _24069_);
  and (_18380_, _18379_, _18377_);
  and (_18381_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_18382_, _18381_, rst);
  or (_18383_, _18382_, _18380_);
  or (_11053_, _18383_, _18376_);
  and (_18384_, _17539_, _23747_);
  and (_18385_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_11057_, _18385_, _18384_);
  and (_18386_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and (_18387_, _16748_, _23898_);
  or (_11062_, _18387_, _18386_);
  and (_18388_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and (_18389_, _16748_, _23824_);
  or (_26959_, _18389_, _18388_);
  and (_18390_, _17396_, _23778_);
  and (_18391_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  or (_11071_, _18391_, _18390_);
  and (_18392_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and (_18393_, _07492_, _23649_);
  or (_11074_, _18393_, _18392_);
  and (_18394_, _17539_, _23946_);
  and (_18395_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_26931_, _18395_, _18394_);
  and (_18396_, _17396_, _23824_);
  and (_18397_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  or (_11077_, _18397_, _18396_);
  and (_18398_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  and (_18399_, _17775_, _23649_);
  or (_11080_, _18399_, _18398_);
  and (_18400_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and (_18401_, _16748_, _23747_);
  or (_11083_, _18401_, _18400_);
  or (_18402_, _24294_, _23939_);
  and (_18403_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_18404_, _18403_, _26118_);
  nand (_18405_, _18225_, _18224_);
  and (_18406_, _18405_, _18404_);
  nor (_18407_, _18406_, _24299_);
  and (_18408_, _18226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_18409_, _18408_, _18407_);
  or (_18410_, _18409_, _24293_);
  and (_18411_, _18410_, _22762_);
  and (_11085_, _18411_, _18402_);
  and (_18412_, _25350_, _24654_);
  nand (_18413_, _18412_, _23594_);
  or (_18414_, _18412_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_18415_, _18414_, _24645_);
  and (_18416_, _18415_, _18413_);
  nand (_18417_, _25358_, _23702_);
  or (_18418_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_18419_, _18418_, _24069_);
  and (_18420_, _18419_, _18417_);
  and (_18421_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_18422_, _18421_, rst);
  or (_18423_, _18422_, _18420_);
  or (_11086_, _18423_, _18416_);
  and (_18424_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and (_18425_, _17775_, _23898_);
  or (_11092_, _18425_, _18424_);
  and (_18426_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and (_18427_, _16748_, _23946_);
  or (_11094_, _18427_, _18426_);
  and (_18428_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  and (_18429_, _16319_, _23707_);
  or (_26971_, _18429_, _18428_);
  and (_18430_, _17539_, _24050_);
  and (_18431_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_26932_, _18431_, _18430_);
  and (_18432_, _17396_, _23747_);
  and (_18433_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  or (_27287_, _18433_, _18432_);
  and (_18434_, _15004_, _23707_);
  and (_18435_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_11100_, _18435_, _18434_);
  and (_18436_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  and (_18437_, _02306_, _23778_);
  or (_11102_, _18437_, _18436_);
  and (_18438_, _17535_, _23778_);
  and (_18439_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_11104_, _18439_, _18438_);
  and (_18440_, _17396_, _24050_);
  and (_18441_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  or (_11106_, _18441_, _18440_);
  and (_18442_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and (_18443_, _16748_, _23707_);
  or (_11109_, _18443_, _18442_);
  and (_18444_, _25439_, _24654_);
  nand (_18445_, _18444_, _23594_);
  or (_18446_, _18444_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_18447_, _18446_, _24645_);
  and (_18448_, _18447_, _18445_);
  nand (_18449_, _25446_, _23702_);
  or (_18450_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_18451_, _18450_, _24069_);
  and (_18452_, _18451_, _18449_);
  and (_18453_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_18454_, _18453_, rst);
  or (_18455_, _18454_, _18452_);
  or (_11111_, _18455_, _18448_);
  and (_18456_, _06602_, _23946_);
  and (_18457_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  or (_11117_, _18457_, _18456_);
  and (_18458_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  and (_18459_, _16742_, _23778_);
  or (_11119_, _18459_, _18458_);
  and (_18460_, _17396_, _23707_);
  and (_18461_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  or (_27288_, _18461_, _18460_);
  and (_18462_, _17535_, _23898_);
  and (_18463_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_11124_, _18463_, _18462_);
  and (_18464_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  and (_18465_, _16742_, _23898_);
  or (_26961_, _18465_, _18464_);
  and (_18466_, _17535_, _23747_);
  and (_18467_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_11127_, _18467_, _18466_);
  and (_18468_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and (_18469_, _13763_, _23824_);
  or (_11132_, _18469_, _18468_);
  and (_18470_, _17378_, _23898_);
  and (_18471_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or (_11134_, _18471_, _18470_);
  and (_18472_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  and (_18473_, _24222_, _23824_);
  or (_11136_, _18473_, _18472_);
  and (_18474_, _17535_, _23649_);
  and (_18475_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_11139_, _18475_, _18474_);
  and (_18476_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  and (_18477_, _16742_, _23824_);
  or (_11141_, _18477_, _18476_);
  and (_18478_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  and (_18479_, _16742_, _23649_);
  or (_11147_, _18479_, _18478_);
  and (_18480_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  and (_18481_, _16742_, _24050_);
  or (_11149_, _18481_, _18480_);
  and (_18482_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_18483_, _17255_, _23707_);
  or (_11153_, _18483_, _18482_);
  and (_18484_, _08198_, _23707_);
  and (_18485_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_11156_, _18485_, _18484_);
  and (_18486_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  and (_18487_, _16742_, _23707_);
  or (_11159_, _18487_, _18486_);
  and (_18488_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and (_18489_, _04761_, _23778_);
  or (_11161_, _18489_, _18488_);
  and (_18490_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  and (_18491_, _08477_, _23778_);
  or (_11164_, _18491_, _18490_);
  and (_18492_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_18493_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or (_18494_, _18493_, _18492_);
  and (_18495_, _18494_, _02393_);
  and (_18496_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_18497_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_18498_, _18497_, _18496_);
  and (_18499_, _18498_, _02445_);
  or (_18500_, _18499_, _18495_);
  and (_18501_, _18500_, _02421_);
  and (_18502_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_18503_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_18504_, _18503_, _18502_);
  and (_18505_, _18504_, _02393_);
  and (_18506_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_18507_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or (_18508_, _18507_, _18506_);
  and (_18509_, _18508_, _02445_);
  or (_18510_, _18509_, _18505_);
  and (_18511_, _18510_, _02459_);
  or (_18512_, _18511_, _18501_);
  and (_18513_, _18512_, _02458_);
  or (_18514_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_18515_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_18516_, _18515_, _18514_);
  and (_18517_, _18516_, _02393_);
  or (_18518_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_18520_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_18521_, _18520_, _18518_);
  and (_18522_, _18521_, _02445_);
  or (_18523_, _18522_, _18517_);
  and (_18524_, _18523_, _02421_);
  or (_18525_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or (_18526_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_18527_, _18526_, _18525_);
  and (_18528_, _18527_, _02393_);
  or (_18529_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_18530_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_18531_, _18530_, _18529_);
  and (_18532_, _18531_, _02445_);
  or (_18533_, _18532_, _18528_);
  and (_18534_, _18533_, _02459_);
  or (_18535_, _18534_, _18524_);
  and (_18536_, _18535_, _02414_);
  or (_18537_, _18536_, _18513_);
  and (_18538_, _18537_, _02398_);
  and (_18539_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and (_18540_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_18541_, _18540_, _18539_);
  and (_18542_, _18541_, _02393_);
  and (_18543_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and (_18544_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_18545_, _18544_, _18543_);
  and (_18546_, _18545_, _02445_);
  or (_18547_, _18546_, _18542_);
  and (_18548_, _18547_, _02421_);
  and (_18549_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and (_18550_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or (_18551_, _18550_, _18549_);
  and (_18552_, _18551_, _02393_);
  and (_18553_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and (_18554_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or (_18555_, _18554_, _18553_);
  and (_18556_, _18555_, _02445_);
  or (_18557_, _18556_, _18552_);
  and (_18558_, _18557_, _02459_);
  or (_18559_, _18558_, _18548_);
  and (_18560_, _18559_, _02458_);
  or (_18561_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or (_18562_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and (_18563_, _18562_, _02445_);
  and (_18564_, _18563_, _18561_);
  or (_18565_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or (_18566_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and (_18567_, _18566_, _02393_);
  and (_18568_, _18567_, _18565_);
  or (_18569_, _18568_, _18564_);
  and (_18570_, _18569_, _02421_);
  or (_18571_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or (_18572_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and (_18573_, _18572_, _02445_);
  and (_18574_, _18573_, _18571_);
  or (_18575_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or (_18576_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and (_18577_, _18576_, _02393_);
  and (_18578_, _18577_, _18575_);
  or (_18579_, _18578_, _18574_);
  and (_18580_, _18579_, _02459_);
  or (_18581_, _18580_, _18570_);
  and (_18582_, _18581_, _02414_);
  or (_18583_, _18582_, _18560_);
  and (_18584_, _18583_, _02496_);
  or (_18585_, _18584_, _18538_);
  and (_18586_, _18585_, _02400_);
  and (_18587_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_18588_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or (_18589_, _18588_, _18587_);
  and (_18590_, _18589_, _02393_);
  and (_18591_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_18592_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or (_18593_, _18592_, _18591_);
  and (_18594_, _18593_, _02445_);
  or (_18595_, _18594_, _18590_);
  or (_18596_, _18595_, _02459_);
  and (_18597_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_18598_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or (_18599_, _18598_, _18597_);
  and (_18601_, _18599_, _02393_);
  and (_18602_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_18603_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or (_18604_, _18603_, _18602_);
  and (_18605_, _18604_, _02445_);
  or (_18606_, _18605_, _18601_);
  or (_18607_, _18606_, _02421_);
  and (_18608_, _18607_, _02458_);
  and (_18609_, _18608_, _18596_);
  or (_18610_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or (_18611_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_18612_, _18611_, _02445_);
  and (_18613_, _18612_, _18610_);
  or (_18614_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or (_18615_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_18616_, _18615_, _02393_);
  and (_18617_, _18616_, _18614_);
  or (_18618_, _18617_, _18613_);
  or (_18619_, _18618_, _02459_);
  or (_18620_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or (_18621_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_18622_, _18621_, _02445_);
  and (_18623_, _18622_, _18620_);
  or (_18624_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or (_18625_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_18626_, _18625_, _02393_);
  and (_18627_, _18626_, _18624_);
  or (_18628_, _18627_, _18623_);
  or (_18629_, _18628_, _02421_);
  and (_18630_, _18629_, _02414_);
  and (_18631_, _18630_, _18619_);
  or (_18632_, _18631_, _18609_);
  and (_18633_, _18632_, _02496_);
  and (_18634_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and (_18635_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_18636_, _18635_, _18634_);
  and (_18637_, _18636_, _02393_);
  and (_18638_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and (_18639_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_18640_, _18639_, _18638_);
  and (_18641_, _18640_, _02445_);
  or (_18642_, _18641_, _18637_);
  or (_18643_, _18642_, _02459_);
  and (_18644_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and (_18645_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_18646_, _18645_, _18644_);
  and (_18647_, _18646_, _02393_);
  and (_18648_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and (_18649_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_18650_, _18649_, _18648_);
  and (_18651_, _18650_, _02445_);
  or (_18652_, _18651_, _18647_);
  or (_18653_, _18652_, _02421_);
  and (_18654_, _18653_, _02458_);
  and (_18655_, _18654_, _18643_);
  or (_18656_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_18657_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and (_18658_, _18657_, _18656_);
  and (_18659_, _18658_, _02393_);
  or (_18660_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_18661_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and (_18662_, _18661_, _18660_);
  and (_18663_, _18662_, _02445_);
  or (_18664_, _18663_, _18659_);
  or (_18665_, _18664_, _02459_);
  or (_18666_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_18667_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and (_18668_, _18667_, _18666_);
  and (_18669_, _18668_, _02393_);
  or (_18670_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_18671_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and (_18672_, _18671_, _18670_);
  and (_18673_, _18672_, _02445_);
  or (_18674_, _18673_, _18669_);
  or (_18675_, _18674_, _02421_);
  and (_18676_, _18675_, _02414_);
  and (_18677_, _18676_, _18665_);
  or (_18678_, _18677_, _18655_);
  and (_18679_, _18678_, _02398_);
  or (_18680_, _18679_, _18633_);
  and (_18681_, _18680_, _02546_);
  or (_18682_, _18681_, _18586_);
  and (_18683_, _18682_, _02646_);
  or (_18684_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_18685_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and (_18686_, _18685_, _02445_);
  and (_18687_, _18686_, _18684_);
  or (_18688_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_18689_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and (_18690_, _18689_, _02393_);
  and (_18691_, _18690_, _18688_);
  or (_18692_, _18691_, _18687_);
  and (_18693_, _18692_, _02459_);
  or (_18694_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_18695_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and (_18696_, _18695_, _02445_);
  and (_18697_, _18696_, _18694_);
  or (_18698_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_18699_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and (_18700_, _18699_, _02393_);
  and (_18701_, _18700_, _18698_);
  or (_18702_, _18701_, _18697_);
  and (_18703_, _18702_, _02421_);
  or (_18704_, _18703_, _18693_);
  and (_18705_, _18704_, _02414_);
  and (_18706_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and (_18707_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_18708_, _18707_, _18706_);
  and (_18709_, _18708_, _02393_);
  and (_18710_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and (_18711_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_18712_, _18711_, _18710_);
  and (_18713_, _18712_, _02445_);
  or (_18714_, _18713_, _18709_);
  and (_18715_, _18714_, _02459_);
  and (_18716_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and (_18717_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_18718_, _18717_, _18716_);
  and (_18719_, _18718_, _02393_);
  and (_18720_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and (_18721_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_18722_, _18721_, _18720_);
  and (_18723_, _18722_, _02445_);
  or (_18724_, _18723_, _18719_);
  and (_18725_, _18724_, _02421_);
  or (_18726_, _18725_, _18715_);
  and (_18727_, _18726_, _02458_);
  or (_18728_, _18727_, _18705_);
  and (_18729_, _18728_, _02496_);
  or (_18730_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_18731_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_18732_, _18731_, _18730_);
  and (_18733_, _18732_, _02393_);
  or (_18734_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_18735_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and (_18736_, _18735_, _18734_);
  and (_18737_, _18736_, _02445_);
  or (_18738_, _18737_, _18733_);
  and (_18739_, _18738_, _02459_);
  or (_18740_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_18741_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_18742_, _18741_, _18740_);
  and (_18743_, _18742_, _02393_);
  or (_18744_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or (_18745_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_18746_, _18745_, _18744_);
  and (_18747_, _18746_, _02445_);
  or (_18748_, _18747_, _18743_);
  and (_18749_, _18748_, _02421_);
  or (_18750_, _18749_, _18739_);
  and (_18751_, _18750_, _02414_);
  and (_18752_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and (_18753_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_18754_, _18753_, _18752_);
  and (_18755_, _18754_, _02393_);
  and (_18756_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_18757_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_18758_, _18757_, _18756_);
  and (_18759_, _18758_, _02445_);
  or (_18760_, _18759_, _18755_);
  and (_18761_, _18760_, _02459_);
  and (_18762_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_18763_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_18764_, _18763_, _18762_);
  and (_18765_, _18764_, _02393_);
  and (_18766_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_18767_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_18768_, _18767_, _18766_);
  and (_18769_, _18768_, _02445_);
  or (_18770_, _18769_, _18765_);
  and (_18771_, _18770_, _02421_);
  or (_18772_, _18771_, _18761_);
  and (_18773_, _18772_, _02458_);
  or (_18774_, _18773_, _18751_);
  and (_18775_, _18774_, _02398_);
  or (_18776_, _18775_, _18729_);
  and (_18777_, _18776_, _02400_);
  and (_18778_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and (_18779_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_18780_, _18779_, _18778_);
  and (_18781_, _18780_, _02393_);
  and (_18782_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and (_18783_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_18784_, _18783_, _18782_);
  and (_18785_, _18784_, _02445_);
  or (_18786_, _18785_, _18781_);
  or (_18787_, _18786_, _02459_);
  and (_18788_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and (_18789_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_18790_, _18789_, _18788_);
  and (_18791_, _18790_, _02393_);
  and (_18792_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and (_18793_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_18794_, _18793_, _18792_);
  and (_18795_, _18794_, _02445_);
  or (_18796_, _18795_, _18791_);
  or (_18797_, _18796_, _02421_);
  and (_18798_, _18797_, _02458_);
  and (_18799_, _18798_, _18787_);
  or (_18800_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_18801_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and (_18802_, _18801_, _18800_);
  and (_18803_, _18802_, _02393_);
  or (_18804_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_18805_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and (_18806_, _18805_, _18804_);
  and (_18807_, _18806_, _02445_);
  or (_18808_, _18807_, _18803_);
  or (_18809_, _18808_, _02459_);
  or (_18810_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_18811_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_18812_, _18811_, _18810_);
  and (_18813_, _18812_, _02393_);
  or (_18814_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_18815_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and (_18816_, _18815_, _18814_);
  and (_18817_, _18816_, _02445_);
  or (_18818_, _18817_, _18813_);
  or (_18819_, _18818_, _02421_);
  and (_18820_, _18819_, _02414_);
  and (_18821_, _18820_, _18809_);
  or (_18822_, _18821_, _18799_);
  and (_18823_, _18822_, _02398_);
  and (_18824_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and (_18825_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_18826_, _18825_, _18824_);
  and (_18827_, _18826_, _02393_);
  and (_18828_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and (_18829_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_18830_, _18829_, _18828_);
  and (_18831_, _18830_, _02445_);
  or (_18832_, _18831_, _18827_);
  or (_18833_, _18832_, _02459_);
  and (_18834_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and (_18835_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_18836_, _18835_, _18834_);
  and (_18837_, _18836_, _02393_);
  and (_18838_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and (_18839_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_18840_, _18839_, _18838_);
  and (_18841_, _18840_, _02445_);
  or (_18842_, _18841_, _18837_);
  or (_18843_, _18842_, _02421_);
  and (_18844_, _18843_, _02458_);
  and (_18845_, _18844_, _18833_);
  or (_18846_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_18847_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and (_18848_, _18847_, _02445_);
  and (_18849_, _18848_, _18846_);
  or (_18850_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_18851_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and (_18852_, _18851_, _02393_);
  and (_18853_, _18852_, _18850_);
  or (_18854_, _18853_, _18849_);
  or (_18855_, _18854_, _02459_);
  or (_18856_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_18857_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and (_18858_, _18857_, _02445_);
  and (_18859_, _18858_, _18856_);
  or (_18860_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_18861_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and (_18862_, _18861_, _02393_);
  and (_18863_, _18862_, _18860_);
  or (_18864_, _18863_, _18859_);
  or (_18865_, _18864_, _02421_);
  and (_18866_, _18865_, _02414_);
  and (_18867_, _18866_, _18855_);
  or (_18868_, _18867_, _18845_);
  and (_18869_, _18868_, _02496_);
  or (_18870_, _18869_, _18823_);
  and (_18871_, _18870_, _02546_);
  or (_18872_, _18871_, _18777_);
  and (_18873_, _18872_, _02405_);
  or (_18874_, _18873_, _18683_);
  and (_18875_, _18874_, _26777_);
  and (_18876_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and (_18877_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_18878_, _18877_, _18876_);
  and (_18879_, _18878_, _02393_);
  and (_18880_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and (_18881_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_18882_, _18881_, _18880_);
  and (_18883_, _18882_, _02445_);
  or (_18884_, _18883_, _18879_);
  and (_18885_, _18884_, _02421_);
  and (_18886_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and (_18887_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_18888_, _18887_, _18886_);
  and (_18889_, _18888_, _02393_);
  and (_18890_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and (_18891_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_18892_, _18891_, _18890_);
  and (_18893_, _18892_, _02445_);
  or (_18894_, _18893_, _18889_);
  and (_18895_, _18894_, _02459_);
  or (_18896_, _18895_, _18885_);
  and (_18897_, _18896_, _02458_);
  or (_18898_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_18899_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and (_18900_, _18899_, _18898_);
  and (_18901_, _18900_, _02393_);
  or (_18902_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_18903_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and (_18904_, _18903_, _18902_);
  and (_18905_, _18904_, _02445_);
  or (_18906_, _18905_, _18901_);
  and (_18907_, _18906_, _02421_);
  or (_18908_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_18909_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and (_18910_, _18909_, _18908_);
  and (_18911_, _18910_, _02393_);
  or (_18912_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_18913_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and (_18914_, _18913_, _18912_);
  and (_18915_, _18914_, _02445_);
  or (_18916_, _18915_, _18911_);
  and (_18917_, _18916_, _02459_);
  or (_18918_, _18917_, _18907_);
  and (_18919_, _18918_, _02414_);
  or (_18920_, _18919_, _18897_);
  and (_18921_, _18920_, _02398_);
  and (_18922_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_18923_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_18924_, _18923_, _18922_);
  and (_18925_, _18924_, _02393_);
  and (_18926_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_18927_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_18928_, _18927_, _18926_);
  and (_18929_, _18928_, _02445_);
  or (_18930_, _18929_, _18925_);
  and (_18931_, _18930_, _02421_);
  and (_18932_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_18933_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_18934_, _18933_, _18932_);
  and (_18935_, _18934_, _02393_);
  and (_18936_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_18937_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_18938_, _18937_, _18936_);
  and (_18939_, _18938_, _02445_);
  or (_18940_, _18939_, _18935_);
  and (_18941_, _18940_, _02459_);
  or (_18942_, _18941_, _18931_);
  and (_18943_, _18942_, _02458_);
  or (_18944_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_18945_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_18946_, _18945_, _02445_);
  and (_18947_, _18946_, _18944_);
  or (_18948_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_18949_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_18950_, _18949_, _02393_);
  and (_18951_, _18950_, _18948_);
  or (_18952_, _18951_, _18947_);
  and (_18953_, _18952_, _02421_);
  or (_18954_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_18955_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_18956_, _18955_, _02445_);
  and (_18957_, _18956_, _18954_);
  or (_18958_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_18959_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_18960_, _18959_, _02393_);
  and (_18961_, _18960_, _18958_);
  or (_18962_, _18961_, _18957_);
  and (_18963_, _18962_, _02459_);
  or (_18964_, _18963_, _18953_);
  and (_18965_, _18964_, _02414_);
  or (_18966_, _18965_, _18943_);
  and (_18967_, _18966_, _02496_);
  or (_18968_, _18967_, _18921_);
  and (_18969_, _18968_, _02400_);
  and (_18970_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and (_18971_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_18972_, _18971_, _18970_);
  and (_18973_, _18972_, _02393_);
  and (_18974_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and (_18975_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_18976_, _18975_, _18974_);
  and (_18977_, _18976_, _02445_);
  or (_18978_, _18977_, _18973_);
  or (_18979_, _18978_, _02459_);
  and (_18980_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and (_18981_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_18982_, _18981_, _18980_);
  and (_18983_, _18982_, _02393_);
  and (_18984_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and (_18985_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_18986_, _18985_, _18984_);
  and (_18987_, _18986_, _02445_);
  or (_18988_, _18987_, _18983_);
  or (_18989_, _18988_, _02421_);
  and (_18990_, _18989_, _02458_);
  and (_18991_, _18990_, _18979_);
  or (_18992_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_18993_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and (_18994_, _18993_, _02445_);
  and (_18995_, _18994_, _18992_);
  or (_18996_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_18997_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and (_18998_, _18997_, _02393_);
  and (_18999_, _18998_, _18996_);
  or (_19000_, _18999_, _18995_);
  or (_19001_, _19000_, _02459_);
  or (_19002_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_19003_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and (_19004_, _19003_, _02445_);
  and (_19005_, _19004_, _19002_);
  or (_19006_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_19007_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and (_19008_, _19007_, _02393_);
  and (_19009_, _19008_, _19006_);
  or (_19010_, _19009_, _19005_);
  or (_19011_, _19010_, _02421_);
  and (_19012_, _19011_, _02414_);
  and (_19013_, _19012_, _19001_);
  or (_19014_, _19013_, _18991_);
  and (_19015_, _19014_, _02496_);
  and (_19016_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_19017_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_19018_, _19017_, _19016_);
  and (_19019_, _19018_, _02393_);
  and (_19020_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and (_19021_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_19022_, _19021_, _19020_);
  and (_19023_, _19022_, _02445_);
  or (_19024_, _19023_, _19019_);
  or (_19025_, _19024_, _02459_);
  and (_19026_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and (_19027_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_19028_, _19027_, _19026_);
  and (_19029_, _19028_, _02393_);
  and (_19030_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and (_19031_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_19032_, _19031_, _19030_);
  and (_19033_, _19032_, _02445_);
  or (_19034_, _19033_, _19029_);
  or (_19035_, _19034_, _02421_);
  and (_19036_, _19035_, _02458_);
  and (_19037_, _19036_, _19025_);
  or (_19038_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_19039_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and (_19040_, _19039_, _19038_);
  and (_19041_, _19040_, _02393_);
  or (_19042_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_19043_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and (_19044_, _19043_, _19042_);
  and (_19045_, _19044_, _02445_);
  or (_19046_, _19045_, _19041_);
  or (_19047_, _19046_, _02459_);
  or (_19048_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_19049_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and (_19050_, _19049_, _19048_);
  and (_19051_, _19050_, _02393_);
  or (_19052_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_19053_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and (_19054_, _19053_, _19052_);
  and (_19055_, _19054_, _02445_);
  or (_19056_, _19055_, _19051_);
  or (_19057_, _19056_, _02421_);
  and (_19058_, _19057_, _02414_);
  and (_19059_, _19058_, _19047_);
  or (_19060_, _19059_, _19037_);
  and (_19061_, _19060_, _02398_);
  or (_19062_, _19061_, _19015_);
  and (_19063_, _19062_, _02546_);
  or (_19064_, _19063_, _18969_);
  and (_19065_, _19064_, _02646_);
  or (_19066_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_19067_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and (_19068_, _19067_, _02445_);
  and (_19069_, _19068_, _19066_);
  or (_19070_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_19071_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and (_19072_, _19071_, _02393_);
  and (_19073_, _19072_, _19070_);
  or (_19074_, _19073_, _19069_);
  and (_19075_, _19074_, _02459_);
  or (_19076_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_19077_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and (_19078_, _19077_, _02445_);
  and (_19079_, _19078_, _19076_);
  or (_19080_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_19081_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and (_19082_, _19081_, _02393_);
  and (_19083_, _19082_, _19080_);
  or (_19084_, _19083_, _19079_);
  and (_19085_, _19084_, _02421_);
  or (_19086_, _19085_, _19075_);
  and (_19087_, _19086_, _02414_);
  and (_19088_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and (_19089_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_19090_, _19089_, _19088_);
  and (_19091_, _19090_, _02393_);
  and (_19092_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and (_19093_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_19094_, _19093_, _19092_);
  and (_19095_, _19094_, _02445_);
  or (_19096_, _19095_, _19091_);
  and (_19097_, _19096_, _02459_);
  and (_19098_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and (_19099_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_19100_, _19099_, _19098_);
  and (_19101_, _19100_, _02393_);
  and (_19102_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and (_19103_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_19104_, _19103_, _19102_);
  and (_19105_, _19104_, _02445_);
  or (_19106_, _19105_, _19101_);
  and (_19107_, _19106_, _02421_);
  or (_19108_, _19107_, _19097_);
  and (_19109_, _19108_, _02458_);
  or (_19110_, _19109_, _19087_);
  and (_19111_, _19110_, _02496_);
  or (_19112_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_19113_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and (_19114_, _19113_, _19112_);
  and (_19115_, _19114_, _02393_);
  or (_19116_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_19117_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and (_19118_, _19117_, _19116_);
  and (_19119_, _19118_, _02445_);
  or (_19120_, _19119_, _19115_);
  and (_19121_, _19120_, _02459_);
  or (_19122_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_19123_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and (_19124_, _19123_, _19122_);
  and (_19125_, _19124_, _02393_);
  or (_19126_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_19127_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and (_19128_, _19127_, _19126_);
  and (_19129_, _19128_, _02445_);
  or (_19130_, _19129_, _19125_);
  and (_19131_, _19130_, _02421_);
  or (_19132_, _19131_, _19121_);
  and (_19133_, _19132_, _02414_);
  and (_19134_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and (_19135_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_19136_, _19135_, _19134_);
  and (_19137_, _19136_, _02393_);
  and (_19138_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and (_19139_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_19140_, _19139_, _19138_);
  and (_19141_, _19140_, _02445_);
  or (_19142_, _19141_, _19137_);
  and (_19143_, _19142_, _02459_);
  and (_19144_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and (_19145_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_19146_, _19145_, _19144_);
  and (_19147_, _19146_, _02393_);
  and (_19148_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and (_19149_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_19150_, _19149_, _19148_);
  and (_19151_, _19150_, _02445_);
  or (_19152_, _19151_, _19147_);
  and (_19153_, _19152_, _02421_);
  or (_19154_, _19153_, _19143_);
  and (_19155_, _19154_, _02458_);
  or (_19156_, _19155_, _19133_);
  and (_19157_, _19156_, _02398_);
  or (_19158_, _19157_, _19111_);
  and (_19159_, _19158_, _02400_);
  and (_19160_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and (_19161_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_19162_, _19161_, _19160_);
  and (_19163_, _19162_, _02393_);
  and (_19164_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and (_19165_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_19166_, _19165_, _19164_);
  and (_19167_, _19166_, _02445_);
  or (_19168_, _19167_, _19163_);
  or (_19169_, _19168_, _02459_);
  and (_19170_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and (_19171_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_19172_, _19171_, _19170_);
  and (_19173_, _19172_, _02393_);
  and (_19174_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and (_19175_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_19176_, _19175_, _19174_);
  and (_19177_, _19176_, _02445_);
  or (_19178_, _19177_, _19173_);
  or (_19179_, _19178_, _02421_);
  and (_19180_, _19179_, _02458_);
  and (_19181_, _19180_, _19169_);
  or (_19182_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_19183_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and (_19184_, _19183_, _19182_);
  and (_19185_, _19184_, _02393_);
  or (_19186_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_19187_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and (_19188_, _19187_, _19186_);
  and (_19189_, _19188_, _02445_);
  or (_19190_, _19189_, _19185_);
  or (_19191_, _19190_, _02459_);
  or (_19192_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_19193_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and (_19194_, _19193_, _19192_);
  and (_19195_, _19194_, _02393_);
  or (_19196_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_19197_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and (_19198_, _19197_, _19196_);
  and (_19199_, _19198_, _02445_);
  or (_19200_, _19199_, _19195_);
  or (_19201_, _19200_, _02421_);
  and (_19202_, _19201_, _02414_);
  and (_19203_, _19202_, _19191_);
  or (_19204_, _19203_, _19181_);
  and (_19205_, _19204_, _02398_);
  and (_19206_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and (_19207_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_19208_, _19207_, _19206_);
  and (_19209_, _19208_, _02393_);
  and (_19210_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and (_19211_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_19212_, _19211_, _19210_);
  and (_19213_, _19212_, _02445_);
  or (_19214_, _19213_, _19209_);
  or (_19215_, _19214_, _02459_);
  and (_19216_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and (_19217_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_19218_, _19217_, _19216_);
  and (_19219_, _19218_, _02393_);
  and (_19220_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and (_19221_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_19222_, _19221_, _19220_);
  and (_19223_, _19222_, _02445_);
  or (_19224_, _19223_, _19219_);
  or (_19225_, _19224_, _02421_);
  and (_19226_, _19225_, _02458_);
  and (_19227_, _19226_, _19215_);
  or (_19228_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_19229_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and (_19230_, _19229_, _02445_);
  and (_19231_, _19230_, _19228_);
  or (_19232_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_19233_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and (_19234_, _19233_, _02393_);
  and (_19235_, _19234_, _19232_);
  or (_19236_, _19235_, _19231_);
  or (_19237_, _19236_, _02459_);
  or (_19238_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_19239_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and (_19240_, _19239_, _02445_);
  and (_19241_, _19240_, _19238_);
  or (_19242_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_19243_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and (_19244_, _19243_, _02393_);
  and (_19245_, _19244_, _19242_);
  or (_19246_, _19245_, _19241_);
  or (_19247_, _19246_, _02421_);
  and (_19248_, _19247_, _02414_);
  and (_19249_, _19248_, _19237_);
  or (_19250_, _19249_, _19227_);
  and (_19251_, _19250_, _02496_);
  or (_19252_, _19251_, _19205_);
  and (_19253_, _19252_, _02546_);
  or (_19254_, _19253_, _19159_);
  and (_19255_, _19254_, _02405_);
  or (_19256_, _19255_, _19065_);
  and (_19257_, _19256_, _02444_);
  or (_19258_, _19257_, _18875_);
  or (_19259_, _19258_, _02443_);
  or (_19260_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_19261_, _19260_, _22762_);
  and (_11175_, _19261_, _19259_);
  and (_19262_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  and (_19263_, _24222_, _23898_);
  or (_11183_, _19263_, _19262_);
  and (_19264_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  and (_19265_, _24222_, _23778_);
  or (_11189_, _19265_, _19264_);
  and (_19266_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  and (_19267_, _17775_, _23747_);
  or (_11193_, _19267_, _19266_);
  and (_19268_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  and (_19269_, _16371_, _23778_);
  or (_11195_, _19269_, _19268_);
  and (_19270_, _18167_, _23649_);
  and (_19271_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or (_11200_, _19271_, _19270_);
  and (_19272_, _18167_, _23747_);
  and (_19273_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or (_11203_, _19273_, _19272_);
  and (_19274_, _18167_, _23824_);
  and (_19275_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or (_27221_, _19275_, _19274_);
  and (_19276_, _06552_, _24050_);
  and (_19277_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_11207_, _19277_, _19276_);
  and (_19278_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and (_19279_, _16371_, _23898_);
  or (_26972_, _19279_, _19278_);
  and (_19280_, _06552_, _23946_);
  and (_19281_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_11216_, _19281_, _19280_);
  and (_19282_, _18217_, _23707_);
  and (_19283_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_11222_, _19283_, _19282_);
  and (_19284_, _17215_, _23898_);
  and (_19285_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or (_11228_, _19285_, _19284_);
  and (_19286_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and (_19287_, _17255_, _24050_);
  or (_11230_, _19287_, _19286_);
  and (_19288_, _17215_, _23778_);
  and (_19289_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  or (_11236_, _19289_, _19288_);
  and (_19290_, _24006_, _23649_);
  and (_19291_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or (_11242_, _19291_, _19290_);
  and (_19292_, _23946_, _23790_);
  and (_19293_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or (_11244_, _19293_, _19292_);
  and (_19294_, _02241_, _23898_);
  and (_19295_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_11246_, _19295_, _19294_);
  and (_19296_, _24050_, _23987_);
  and (_19297_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or (_26937_, _19297_, _19296_);
  and (_19298_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and (_19299_, _13763_, _23898_);
  or (_27243_, _19299_, _19298_);
  and (_19300_, _23987_, _23649_);
  and (_19301_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  or (_11252_, _19301_, _19300_);
  and (_19302_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and (_19303_, _13763_, _23778_);
  or (_11255_, _19303_, _19302_);
  and (_19304_, _02241_, _23778_);
  and (_19305_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_11258_, _19305_, _19304_);
  and (_19306_, _23898_, _23790_);
  and (_19307_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or (_11262_, _19307_, _19306_);
  and (_19308_, _06552_, _23707_);
  and (_19309_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_11265_, _19309_, _19308_);
  and (_19310_, _02326_, _23747_);
  and (_19311_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_11267_, _19311_, _19310_);
  and (_19312_, _02241_, _23824_);
  and (_19313_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_27292_, _19313_, _19312_);
  and (_19314_, _07743_, _23946_);
  and (_19315_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or (_11270_, _19315_, _19314_);
  and (_19316_, _24086_, _23747_);
  and (_19317_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_11273_, _19317_, _19316_);
  and (_19318_, _23987_, _23946_);
  and (_19319_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  or (_26936_, _19319_, _19318_);
  and (_19320_, _01971_, _23707_);
  and (_19321_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or (_11280_, _19321_, _19320_);
  and (_19322_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  and (_19323_, _16319_, _23747_);
  or (_11286_, _19323_, _19322_);
  and (_19324_, _23907_, _23778_);
  and (_19325_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_11289_, _19325_, _19324_);
  and (_19326_, _23907_, _23824_);
  and (_19327_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_11296_, _19327_, _19326_);
  and (_19328_, _23912_, _23649_);
  and (_19329_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  or (_11299_, _19329_, _19328_);
  and (_19330_, _02241_, _23946_);
  and (_19331_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_11307_, _19331_, _19330_);
  and (_19332_, _02241_, _23707_);
  and (_19333_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_11312_, _19333_, _19332_);
  and (_19334_, _24006_, _23778_);
  and (_19335_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  or (_11315_, _19335_, _19334_);
  and (_19336_, _24006_, _23824_);
  and (_19337_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or (_11317_, _19337_, _19336_);
  and (_19338_, _23987_, _23707_);
  and (_19339_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  or (_11319_, _19339_, _19338_);
  and (_19340_, _24086_, _24050_);
  and (_19341_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_27256_, _19341_, _19340_);
  and (_19342_, _24011_, _23946_);
  and (_19343_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_11322_, _19343_, _19342_);
  and (_19344_, _02241_, _23649_);
  and (_19345_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_27294_, _19345_, _19344_);
  and (_19346_, _24006_, _23898_);
  and (_19347_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or (_11329_, _19347_, _19346_);
  and (_19348_, _02241_, _24050_);
  and (_19349_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_11331_, _19349_, _19348_);
  and (_19350_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and (_19351_, _07513_, _23747_);
  or (_11335_, _19351_, _19350_);
  and (_19352_, _23912_, _23778_);
  and (_19353_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  or (_11341_, _19353_, _19352_);
  and (_19354_, _24050_, _23907_);
  and (_19355_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_11346_, _19355_, _19354_);
  and (_19356_, _23992_, _23898_);
  and (_19357_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_11349_, _19357_, _19356_);
  and (_19358_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and (_19359_, _13763_, _23649_);
  or (_27244_, _19359_, _19358_);
  and (_19360_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and (_19361_, _24203_, _23898_);
  or (_11353_, _19361_, _19360_);
  and (_19362_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and (_19363_, _24276_, _24050_);
  or (_27251_, _19363_, _19362_);
  and (_19364_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and (_19365_, _24276_, _23778_);
  or (_11356_, _19365_, _19364_);
  and (_19366_, _01971_, _24050_);
  and (_19367_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  or (_11358_, _19367_, _19366_);
  and (_19368_, _17378_, _23649_);
  and (_19369_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  or (_27291_, _19369_, _19368_);
  and (_19370_, _17378_, _24050_);
  and (_19371_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or (_11364_, _19371_, _19370_);
  and (_19372_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  and (_19373_, _13763_, _23747_);
  or (_11368_, _19373_, _19372_);
  and (_19374_, _23987_, _23898_);
  and (_19375_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  or (_11374_, _19375_, _19374_);
  and (_19376_, _23987_, _23824_);
  and (_19377_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  or (_11376_, _19377_, _19376_);
  and (_19378_, _17378_, _23707_);
  and (_19379_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or (_11388_, _19379_, _19378_);
  and (_19380_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  and (_19381_, _24276_, _23747_);
  or (_11394_, _19381_, _19380_);
  and (_19382_, _01971_, _23946_);
  and (_19383_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or (_11396_, _19383_, _19382_);
  and (_19384_, _17535_, _23707_);
  and (_19385_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_26935_, _19385_, _19384_);
  and (_19386_, _07743_, _23649_);
  and (_19387_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  or (_11400_, _19387_, _19386_);
  and (_19388_, _17378_, _23747_);
  and (_19389_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or (_27290_, _19389_, _19388_);
  and (_19390_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  and (_19391_, _24222_, _24050_);
  or (_11404_, _19391_, _19390_);
  and (_19392_, _23987_, _23778_);
  and (_19393_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or (_11406_, _19393_, _19392_);
  and (_19394_, _17378_, _23946_);
  and (_19395_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or (_11408_, _19395_, _19394_);
  and (_19396_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  and (_19397_, _16018_, _24050_);
  or (_11410_, _19397_, _19396_);
  and (_19398_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  and (_19399_, _16319_, _23946_);
  or (_11414_, _19399_, _19398_);
  and (_19400_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  and (_19401_, _24203_, _23649_);
  or (_11418_, _19401_, _19400_);
  and (_19402_, _17221_, _23747_);
  and (_19403_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_11425_, _19403_, _19402_);
  and (_19404_, _06552_, _23747_);
  and (_19405_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_27144_, _19405_, _19404_);
  and (_19406_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  and (_19407_, _16018_, _23649_);
  or (_26965_, _19407_, _19406_);
  and (_19408_, _17215_, _23824_);
  and (_19409_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  or (_27217_, _19409_, _19408_);
  and (_19410_, _06552_, _23824_);
  and (_19411_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_11454_, _19411_, _19410_);
  and (_19412_, _25156_, _23946_);
  and (_19413_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_11456_, _19413_, _19412_);
  and (_19414_, _25156_, _23747_);
  and (_19415_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_11458_, _19415_, _19414_);
  and (_19416_, _25091_, _24050_);
  and (_19417_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  or (_11460_, _19417_, _19416_);
  and (_19418_, _25091_, _23649_);
  and (_19419_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  or (_11463_, _19419_, _19418_);
  and (_19420_, _17215_, _23649_);
  and (_19422_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  or (_11468_, _19422_, _19420_);
  and (_19423_, _25079_, _23747_);
  and (_19424_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or (_11471_, _19424_, _19423_);
  and (_19425_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and (_19426_, _17091_, _23747_);
  or (_11473_, _19426_, _19425_);
  and (_19427_, _24999_, _23649_);
  and (_19428_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_27184_, _19428_, _19427_);
  and (_19429_, _24932_, _23649_);
  and (_19430_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_11478_, _19430_, _19429_);
  and (_19431_, _24932_, _23778_);
  and (_19432_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_27179_, _19432_, _19431_);
  and (_19433_, _08198_, _24050_);
  and (_19434_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_11483_, _19434_, _19433_);
  and (_19435_, _24858_, _23946_);
  and (_19436_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or (_11485_, _19436_, _19435_);
  and (_19437_, _24858_, _23824_);
  and (_19438_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or (_11487_, _19438_, _19437_);
  and (_19439_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  and (_19440_, _17091_, _23824_);
  or (_11489_, _19440_, _19439_);
  and (_19441_, _24839_, _23707_);
  and (_19442_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  or (_11491_, _19442_, _19441_);
  and (_19443_, _24839_, _23747_);
  and (_19444_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  or (_11493_, _19444_, _19443_);
  and (_19445_, _17215_, _23747_);
  and (_19446_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  or (_11497_, _19446_, _19445_);
  and (_19447_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and (_19448_, _16375_, _23707_);
  or (_11499_, _19448_, _19447_);
  and (_19449_, _24789_, _23946_);
  and (_19450_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_11502_, _19450_, _19449_);
  and (_19451_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and (_19452_, _16375_, _24050_);
  or (_26970_, _19452_, _19451_);
  and (_19453_, _24789_, _23898_);
  and (_19454_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_11505_, _19454_, _19453_);
  and (_19455_, _24722_, _24050_);
  and (_19456_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  or (_11506_, _19456_, _19455_);
  and (_19457_, _24722_, _23824_);
  and (_19458_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  or (_11510_, _19458_, _19457_);
  and (_19459_, _24121_, _23816_);
  nor (_19460_, _14722_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_19461_, _19460_, _14723_);
  nand (_19462_, _19461_, _24174_);
  or (_19463_, _24174_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_19464_, _19463_, _19462_);
  nand (_19465_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_19466_, _19465_, _24127_);
  or (_19467_, _19466_, _19464_);
  and (_19468_, _19467_, _24166_);
  or (_11512_, _19468_, _19459_);
  and (_19469_, _07743_, _23747_);
  and (_19470_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  or (_11515_, _19470_, _19469_);
  and (_19471_, _24688_, _24050_);
  and (_19472_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or (_11519_, _19472_, _19471_);
  and (_19473_, _24688_, _23824_);
  and (_19474_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or (_11522_, _19474_, _19473_);
  and (_19475_, _24688_, _23778_);
  and (_19476_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  or (_11524_, _19476_, _19475_);
  and (_19477_, _17221_, _23824_);
  and (_19478_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_11526_, _19478_, _19477_);
  and (_19479_, _24639_, _23707_);
  and (_19480_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_11528_, _19480_, _19479_);
  and (_19481_, _24375_, _23649_);
  and (_19482_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_11532_, _19482_, _19481_);
  and (_19483_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and (_19484_, _17091_, _24050_);
  or (_11534_, _19484_, _19483_);
  and (_19485_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and (_19486_, _01967_, _23649_);
  or (_11538_, _19486_, _19485_);
  and (_19487_, _25091_, _23778_);
  and (_19488_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or (_11539_, _19488_, _19487_);
  and (_19489_, _25079_, _23946_);
  and (_19490_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  or (_11541_, _19490_, _19489_);
  and (_19491_, _25079_, _23898_);
  and (_19492_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or (_11543_, _19492_, _19491_);
  and (_19493_, _24999_, _24050_);
  and (_19494_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_11545_, _19494_, _19493_);
  and (_19495_, _24999_, _23898_);
  and (_19496_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_11548_, _19496_, _19495_);
  and (_19497_, _24932_, _24050_);
  and (_19498_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_27181_, _19498_, _19497_);
  and (_19499_, _24932_, _23824_);
  and (_19500_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_27180_, _19500_, _19499_);
  and (_19501_, _24858_, _23707_);
  and (_19502_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or (_11562_, _19502_, _19501_);
  and (_19503_, _24950_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_19504_, _24865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_19505_, _24865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_19506_, _19505_, _19504_);
  nor (_19507_, _19506_, _02137_);
  or (_19508_, _19507_, _24862_);
  or (_19509_, _19508_, _19503_);
  or (_19510_, _19506_, _24954_);
  and (_19511_, _19510_, _22762_);
  and (_11565_, _19511_, _19509_);
  and (_19512_, _15004_, _23778_);
  and (_19513_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or (_11568_, _19513_, _19512_);
  and (_19514_, _24839_, _23778_);
  and (_19515_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  or (_11569_, _19515_, _19514_);
  and (_19516_, _24645_, _24076_);
  and (_19517_, _19516_, _24064_);
  nand (_19518_, _19517_, _23711_);
  or (_19519_, _25039_, _24961_);
  and (_19520_, _19519_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_19521_, _19520_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and (_19522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _24865_);
  and (_19523_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_19524_, _19523_, _19522_);
  nor (_19525_, _19524_, _24864_);
  nor (_19526_, _02156_, _02121_);
  nor (_19527_, _19526_, _24864_);
  nor (_19528_, _19527_, _19525_);
  nand (_19529_, _19528_, _19521_);
  nand (_19530_, _19529_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_19531_, _19530_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_19532_, _19531_, _19517_);
  and (_19533_, _19532_, _19518_);
  nand (_19534_, _19533_, _24817_);
  or (_19535_, _24817_, _23892_);
  and (_19536_, _19535_, _22762_);
  and (_11577_, _19536_, _19534_);
  and (_19537_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and (_19538_, _17091_, _23946_);
  or (_11591_, _19538_, _19537_);
  and (_19539_, _06552_, _23649_);
  and (_19540_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_11595_, _19540_, _19539_);
  and (_11604_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _22762_);
  and (_19541_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and (_19542_, _17091_, _23649_);
  or (_27242_, _19542_, _19541_);
  and (_19543_, _24688_, _23649_);
  and (_19544_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or (_11609_, _19544_, _19543_);
  and (_19545_, _24375_, _23898_);
  and (_19546_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_11613_, _19546_, _19545_);
  and (_19547_, _25156_, _23707_);
  and (_19548_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_11615_, _19548_, _19547_);
  and (_19549_, _25156_, _23778_);
  and (_19550_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_11617_, _19550_, _19549_);
  and (_19551_, _24858_, _23747_);
  and (_19552_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or (_11621_, _19552_, _19551_);
  and (_19553_, _24839_, _23649_);
  and (_19554_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  or (_11622_, _19554_, _19553_);
  and (_19555_, _24789_, _23824_);
  and (_19556_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_11625_, _19556_, _19555_);
  and (_19557_, _24722_, _23747_);
  and (_19558_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or (_27174_, _19558_, _19557_);
  and (_19559_, _24375_, _23946_);
  and (_19560_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_11628_, _19560_, _19559_);
  and (_19561_, _25091_, _23898_);
  and (_19562_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  or (_27186_, _19562_, _19561_);
  and (_19563_, _24999_, _23824_);
  and (_19564_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_27182_, _19564_, _19563_);
  not (_19565_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_19566_, _19520_, _19565_);
  nand (_19567_, _19526_, _19525_);
  or (_19568_, _19567_, _19566_);
  and (_19569_, _19568_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_19570_, _19569_, _06778_);
  and (_19571_, _24813_, _24654_);
  or (_19572_, _19571_, _19570_);
  nand (_19573_, _19571_, _23594_);
  and (_19574_, _19573_, _19572_);
  or (_19575_, _19574_, _24816_);
  nand (_19576_, _24816_, _23702_);
  and (_19577_, _19576_, _22762_);
  and (_11637_, _19577_, _19575_);
  and (_11643_, _26274_, _22762_);
  and (_19578_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  and (_19579_, _16319_, _23778_);
  or (_11645_, _19579_, _19578_);
  nand (_19580_, _23018_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_19581_, _19580_, _24653_);
  or (_19582_, _19581_, _05827_);
  and (_19583_, _19582_, _24813_);
  nand (_19584_, _24813_, _23018_);
  and (_19585_, _19584_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_19586_, _19585_, _24816_);
  or (_19587_, _19586_, _19583_);
  or (_19588_, _24817_, _24043_);
  and (_19589_, _19588_, _22762_);
  and (_11651_, _19589_, _19587_);
  and (_19590_, _24892_, _24880_);
  nand (_19591_, _24895_, _19590_);
  nand (_19592_, _24905_, _24902_);
  and (_19593_, _19592_, _24896_);
  or (_19594_, _19593_, _24895_);
  and (_19595_, _19594_, _24938_);
  and (_19596_, _19595_, _19591_);
  or (_19597_, _19596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_19598_, _24938_);
  not (_19599_, _24918_);
  or (_19600_, _19599_, _24914_);
  or (_19601_, _24889_, _24870_);
  and (_19602_, _19601_, _19600_);
  or (_19603_, _19602_, _19598_);
  and (_19604_, _19603_, _22762_);
  and (_11656_, _19604_, _19597_);
  and (_19605_, _04922_, _23778_);
  and (_19606_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  or (_11659_, _19606_, _19605_);
  and (_11662_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _22762_);
  and (_19607_, _19594_, _24863_);
  and (_19608_, _19607_, _19591_);
  or (_19609_, _19608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  not (_19610_, _24863_);
  or (_19611_, _19602_, _19610_);
  and (_19612_, _19611_, _22762_);
  and (_11663_, _19612_, _19609_);
  and (_11665_, _26366_, _22762_);
  and (_19613_, _25142_, _23707_);
  and (_19614_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or (_27201_, _19614_, _19613_);
  not (_19615_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_19616_, _19615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not (_19617_, _19525_);
  and (_19618_, _19527_, _19617_);
  not (_19619_, _19618_);
  or (_19620_, _19619_, _19566_);
  and (_19621_, _19620_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_19622_, _19621_, _19616_);
  and (_19623_, _24813_, _24125_);
  or (_19624_, _19623_, _19622_);
  nand (_19625_, _19623_, _23594_);
  and (_19626_, _19625_, _19624_);
  or (_19627_, _19626_, _24816_);
  or (_19628_, _24817_, _23939_);
  and (_19629_, _19628_, _22762_);
  and (_11677_, _19629_, _19627_);
  nand (_19630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_19631_, _19618_, _19521_);
  nor (_19632_, _19631_, _19630_);
  and (_19633_, _24118_, _23003_);
  and (_19634_, _19633_, _24064_);
  nand (_19635_, _24645_, _19634_);
  nand (_19636_, _19635_, _19632_);
  or (_19637_, _19635_, _23594_);
  and (_19638_, _19637_, _19636_);
  nand (_19639_, _19638_, _24817_);
  or (_19640_, _24817_, _23738_);
  and (_19641_, _19640_, _22762_);
  and (_11683_, _19641_, _19639_);
  and (_19642_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  and (_19643_, _16018_, _23946_);
  or (_11684_, _19643_, _19642_);
  and (_19644_, _24654_, _24648_);
  nand (_19645_, _19644_, _23594_);
  or (_19646_, _19644_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_19647_, _19646_, _24659_);
  and (_19648_, _19647_, _19645_);
  nor (_19649_, _24659_, _23702_);
  or (_19650_, _19649_, _19648_);
  and (_11687_, _19650_, _22762_);
  nor (_19651_, _14721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_19652_, _19651_, _14722_);
  and (_19653_, _19652_, _24174_);
  and (_19654_, _14719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_19655_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_19656_, _19655_, _24127_);
  or (_19657_, _19656_, _19654_);
  or (_19658_, _19657_, _19653_);
  and (_19659_, _19658_, _24171_);
  and (_19660_, _24120_, _23892_);
  or (_19661_, _19660_, _19659_);
  and (_11690_, _19661_, _22762_);
  and (_19662_, _17221_, _23898_);
  and (_19663_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_11694_, _19663_, _19662_);
  and (_19664_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  and (_19665_, _02306_, _24050_);
  or (_11696_, _19665_, _19664_);
  and (_19666_, _05119_, _23747_);
  and (_19667_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  or (_11698_, _19667_, _19666_);
  nand (_19668_, _24950_, _24864_);
  nand (_19669_, _19504_, _24862_);
  and (_19670_, _19669_, _22762_);
  and (_11704_, _19670_, _19668_);
  and (_19671_, _25754_, _23778_);
  and (_19672_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  or (_27033_, _19672_, _19671_);
  and (_19673_, _01759_, _23747_);
  and (_19674_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_11707_, _19674_, _19673_);
  and (_19675_, _24730_, _24654_);
  nand (_19676_, _19675_, _23594_);
  or (_19677_, _19675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_19678_, _19677_, _19676_);
  or (_19679_, _19678_, _24736_);
  nand (_19680_, _24736_, _23702_);
  and (_19681_, _19680_, _22762_);
  and (_11710_, _19681_, _19679_);
  and (_19682_, _02215_, _24050_);
  and (_19683_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_11711_, _19683_, _19682_);
  and (_19684_, _02350_, _23824_);
  and (_19685_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_11715_, _19685_, _19684_);
  and (_19686_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  and (_19687_, _02306_, _23946_);
  or (_11718_, _19687_, _19686_);
  and (_19688_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  and (_19689_, _02306_, _23649_);
  or (_11721_, _19689_, _19688_);
  and (_19690_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and (_19691_, _16375_, _23824_);
  or (_11723_, _19691_, _19690_);
  and (_19692_, _08642_, _23707_);
  and (_19693_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  or (_11724_, _19693_, _19692_);
  and (_19694_, _05298_, _23898_);
  and (_19695_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_11726_, _19695_, _19694_);
  and (_19696_, _05346_, _23649_);
  and (_19697_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_11728_, _19697_, _19696_);
  and (_19698_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and (_19699_, _16375_, _23747_);
  or (_26969_, _19699_, _19698_);
  and (_19700_, _08642_, _24050_);
  and (_19701_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  or (_11733_, _19701_, _19700_);
  and (_19702_, _05429_, _23898_);
  and (_19703_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_11734_, _19703_, _19702_);
  and (_19704_, _06615_, _23707_);
  and (_19705_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_11738_, _19705_, _19704_);
  or (_19706_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_11754_, _19706_, _05482_);
  and (_19707_, _15004_, _23898_);
  and (_19708_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_11755_, _19708_, _19707_);
  nor (_11758_, _00759_, rst);
  and (_11759_, _00341_, _22762_);
  and (_11762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _22762_);
  and (_19709_, _05119_, _23649_);
  and (_19710_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or (_11783_, _19710_, _19709_);
  and (_19711_, _25571_, _24050_);
  and (_19712_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_11787_, _19712_, _19711_);
  and (_19713_, _02087_, _23946_);
  and (_19714_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_27009_, _19714_, _19713_);
  and (_19715_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and (_19716_, _17091_, _23778_);
  or (_27241_, _19716_, _19715_);
  and (_19717_, _04656_, _23946_);
  and (_19718_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_11791_, _19718_, _19717_);
  and (_19719_, _04832_, _23898_);
  and (_19720_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_11793_, _19720_, _19719_);
  or (_19721_, _05223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_11795_, _19721_, _05224_);
  and (_19722_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_19723_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_19724_, _19723_, _19722_);
  and (_19725_, _19724_, _02393_);
  and (_19726_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_19727_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or (_19728_, _19727_, _19726_);
  and (_19729_, _19728_, _02445_);
  or (_19730_, _19729_, _19725_);
  and (_19731_, _19730_, _02421_);
  and (_19732_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and (_19733_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_19734_, _19733_, _19732_);
  and (_19735_, _19734_, _02393_);
  and (_19736_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_19737_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or (_19738_, _19737_, _19736_);
  and (_19739_, _19738_, _02445_);
  or (_19740_, _19739_, _19735_);
  and (_19741_, _19740_, _02459_);
  or (_19742_, _19741_, _19731_);
  and (_19743_, _19742_, _02458_);
  or (_19744_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or (_19745_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_19746_, _19745_, _19744_);
  and (_19747_, _19746_, _02393_);
  or (_19748_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or (_19749_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_19750_, _19749_, _19748_);
  and (_19751_, _19750_, _02445_);
  or (_19752_, _19751_, _19747_);
  and (_19753_, _19752_, _02421_);
  or (_19754_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_19755_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and (_19756_, _19755_, _19754_);
  and (_19757_, _19756_, _02393_);
  or (_19758_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or (_19759_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_19760_, _19759_, _19758_);
  and (_19761_, _19760_, _02445_);
  or (_19762_, _19761_, _19757_);
  and (_19763_, _19762_, _02459_);
  or (_19764_, _19763_, _19753_);
  and (_19765_, _19764_, _02414_);
  or (_19766_, _19765_, _19743_);
  and (_19767_, _19766_, _02398_);
  and (_19768_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and (_19769_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or (_19770_, _19769_, _19768_);
  and (_19771_, _19770_, _02393_);
  and (_19772_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and (_19773_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or (_19774_, _19773_, _19772_);
  and (_19775_, _19774_, _02445_);
  or (_19776_, _19775_, _19771_);
  and (_19777_, _19776_, _02421_);
  and (_19778_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and (_19779_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or (_19780_, _19779_, _19778_);
  and (_19781_, _19780_, _02393_);
  and (_19782_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and (_19783_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or (_19784_, _19783_, _19782_);
  and (_19785_, _19784_, _02445_);
  or (_19786_, _19785_, _19781_);
  and (_19787_, _19786_, _02459_);
  or (_19788_, _19787_, _19777_);
  and (_19789_, _19788_, _02458_);
  or (_19790_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or (_19791_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and (_19792_, _19791_, _02445_);
  and (_19793_, _19792_, _19790_);
  or (_19794_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or (_19795_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and (_19796_, _19795_, _02393_);
  and (_19797_, _19796_, _19794_);
  or (_19798_, _19797_, _19793_);
  and (_19799_, _19798_, _02421_);
  or (_19800_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or (_19801_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and (_19802_, _19801_, _02445_);
  and (_19803_, _19802_, _19800_);
  or (_19804_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or (_19805_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and (_19806_, _19805_, _02393_);
  and (_19807_, _19806_, _19804_);
  or (_19808_, _19807_, _19803_);
  and (_19809_, _19808_, _02459_);
  or (_19810_, _19809_, _19799_);
  and (_19811_, _19810_, _02414_);
  or (_19812_, _19811_, _19789_);
  and (_19813_, _19812_, _02496_);
  or (_19814_, _19813_, _19767_);
  and (_19815_, _19814_, _02400_);
  and (_19816_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_19817_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or (_19818_, _19817_, _19816_);
  and (_19819_, _19818_, _02393_);
  and (_19820_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_19821_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or (_19822_, _19821_, _19820_);
  and (_19823_, _19822_, _02445_);
  or (_19824_, _19823_, _19819_);
  or (_19825_, _19824_, _02459_);
  and (_19826_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_19827_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or (_19828_, _19827_, _19826_);
  and (_19829_, _19828_, _02393_);
  and (_19830_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_19831_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or (_19832_, _19831_, _19830_);
  and (_19833_, _19832_, _02445_);
  or (_19834_, _19833_, _19829_);
  or (_19835_, _19834_, _02421_);
  and (_19836_, _19835_, _02458_);
  and (_19837_, _19836_, _19825_);
  or (_19838_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or (_19839_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_19840_, _19839_, _02445_);
  and (_19841_, _19840_, _19838_);
  or (_19842_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or (_19843_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_19844_, _19843_, _02393_);
  and (_19845_, _19844_, _19842_);
  or (_19846_, _19845_, _19841_);
  or (_19847_, _19846_, _02459_);
  or (_19848_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or (_19849_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_19850_, _19849_, _02445_);
  and (_19851_, _19850_, _19848_);
  or (_19852_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or (_19853_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_19854_, _19853_, _02393_);
  and (_19855_, _19854_, _19852_);
  or (_19856_, _19855_, _19851_);
  or (_19857_, _19856_, _02421_);
  and (_19858_, _19857_, _02414_);
  and (_19859_, _19858_, _19847_);
  or (_19860_, _19859_, _19837_);
  and (_19861_, _19860_, _02496_);
  and (_19862_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and (_19863_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_19864_, _19863_, _19862_);
  and (_19865_, _19864_, _02393_);
  and (_19866_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and (_19867_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_19868_, _19867_, _19866_);
  and (_19869_, _19868_, _02445_);
  or (_19870_, _19869_, _19865_);
  or (_19871_, _19870_, _02459_);
  and (_19872_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and (_19873_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_19874_, _19873_, _19872_);
  and (_19875_, _19874_, _02393_);
  and (_19876_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and (_19877_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_19878_, _19877_, _19876_);
  and (_19879_, _19878_, _02445_);
  or (_19880_, _19879_, _19875_);
  or (_19881_, _19880_, _02421_);
  and (_19882_, _19881_, _02458_);
  and (_19883_, _19882_, _19871_);
  or (_19884_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_19885_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and (_19886_, _19885_, _19884_);
  and (_19887_, _19886_, _02393_);
  or (_19888_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_19889_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and (_19890_, _19889_, _19888_);
  and (_19891_, _19890_, _02445_);
  or (_19892_, _19891_, _19887_);
  or (_19893_, _19892_, _02459_);
  or (_19894_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_19895_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and (_19896_, _19895_, _19894_);
  and (_19897_, _19896_, _02393_);
  or (_19898_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_19899_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and (_19900_, _19899_, _19898_);
  and (_19901_, _19900_, _02445_);
  or (_19902_, _19901_, _19897_);
  or (_19903_, _19902_, _02421_);
  and (_19904_, _19903_, _02414_);
  and (_19905_, _19904_, _19893_);
  or (_19906_, _19905_, _19883_);
  and (_19907_, _19906_, _02398_);
  or (_19908_, _19907_, _19861_);
  and (_19909_, _19908_, _02546_);
  or (_19910_, _19909_, _19815_);
  and (_19911_, _19910_, _02646_);
  or (_19912_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_19913_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and (_19914_, _19913_, _02445_);
  and (_19915_, _19914_, _19912_);
  or (_19916_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_19917_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and (_19918_, _19917_, _02393_);
  and (_19919_, _19918_, _19916_);
  or (_19921_, _19919_, _19915_);
  and (_19922_, _19921_, _02459_);
  or (_19923_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_19924_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and (_19925_, _19924_, _02445_);
  and (_19926_, _19925_, _19923_);
  or (_19927_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_19928_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and (_19929_, _19928_, _02393_);
  and (_19930_, _19929_, _19927_);
  or (_19931_, _19930_, _19926_);
  and (_19932_, _19931_, _02421_);
  or (_19933_, _19932_, _19922_);
  and (_19934_, _19933_, _02414_);
  and (_19935_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and (_19936_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_19937_, _19936_, _19935_);
  and (_19938_, _19937_, _02393_);
  and (_19939_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and (_19940_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_19942_, _19940_, _19939_);
  and (_19943_, _19942_, _02445_);
  or (_19944_, _19943_, _19938_);
  and (_19945_, _19944_, _02459_);
  and (_19946_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and (_19947_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_19948_, _19947_, _19946_);
  and (_19949_, _19948_, _02393_);
  and (_19950_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and (_19951_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_19952_, _19951_, _19950_);
  and (_19953_, _19952_, _02445_);
  or (_19954_, _19953_, _19949_);
  and (_19955_, _19954_, _02421_);
  or (_19956_, _19955_, _19945_);
  and (_19957_, _19956_, _02458_);
  or (_19958_, _19957_, _19934_);
  and (_19959_, _19958_, _02496_);
  or (_19960_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or (_19961_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_19962_, _19961_, _19960_);
  and (_19963_, _19962_, _02393_);
  or (_19964_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or (_19965_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_19966_, _19965_, _19964_);
  and (_19967_, _19966_, _02445_);
  or (_19968_, _19967_, _19963_);
  and (_19969_, _19968_, _02459_);
  or (_19970_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or (_19971_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_19973_, _19971_, _19970_);
  and (_19974_, _19973_, _02393_);
  or (_19975_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_19976_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and (_19977_, _19976_, _19975_);
  and (_19978_, _19977_, _02445_);
  or (_19979_, _19978_, _19974_);
  and (_19980_, _19979_, _02421_);
  or (_19981_, _19980_, _19969_);
  and (_19982_, _19981_, _02414_);
  and (_19983_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_19984_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_19985_, _19984_, _19983_);
  and (_19986_, _19985_, _02393_);
  and (_19987_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and (_19988_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or (_19989_, _19988_, _19987_);
  and (_19990_, _19989_, _02445_);
  or (_19991_, _19990_, _19986_);
  and (_19992_, _19991_, _02459_);
  and (_19993_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_19994_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_19995_, _19994_, _19993_);
  and (_19996_, _19995_, _02393_);
  and (_19997_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and (_19998_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or (_19999_, _19998_, _19997_);
  and (_20000_, _19999_, _02445_);
  or (_20001_, _20000_, _19996_);
  and (_20002_, _20001_, _02421_);
  or (_20003_, _20002_, _19992_);
  and (_20004_, _20003_, _02458_);
  or (_20005_, _20004_, _19982_);
  and (_20006_, _20005_, _02398_);
  or (_20007_, _20006_, _19959_);
  and (_20008_, _20007_, _02400_);
  and (_20009_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and (_20010_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_20011_, _20010_, _20009_);
  and (_20012_, _20011_, _02393_);
  and (_20013_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and (_20014_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_20015_, _20014_, _20013_);
  and (_20016_, _20015_, _02445_);
  or (_20017_, _20016_, _20012_);
  or (_20018_, _20017_, _02459_);
  and (_20019_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and (_20020_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_20021_, _20020_, _20019_);
  and (_20022_, _20021_, _02393_);
  and (_20023_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and (_20024_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_20025_, _20024_, _20023_);
  and (_20026_, _20025_, _02445_);
  or (_20027_, _20026_, _20022_);
  or (_20028_, _20027_, _02421_);
  and (_20029_, _20028_, _02458_);
  and (_20030_, _20029_, _20018_);
  or (_20031_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_20032_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and (_20033_, _20032_, _20031_);
  and (_20034_, _20033_, _02393_);
  or (_20035_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_20036_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and (_20037_, _20036_, _20035_);
  and (_20038_, _20037_, _02445_);
  or (_20039_, _20038_, _20034_);
  or (_20040_, _20039_, _02459_);
  or (_20041_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_20042_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and (_20044_, _20042_, _20041_);
  and (_20045_, _20044_, _02393_);
  or (_20046_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_20047_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and (_20048_, _20047_, _20046_);
  and (_20049_, _20048_, _02445_);
  or (_20050_, _20049_, _20045_);
  or (_20051_, _20050_, _02421_);
  and (_20052_, _20051_, _02414_);
  and (_20053_, _20052_, _20040_);
  or (_20054_, _20053_, _20030_);
  and (_20055_, _20054_, _02398_);
  and (_20056_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and (_20057_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_20058_, _20057_, _20056_);
  and (_20059_, _20058_, _02393_);
  and (_20060_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and (_20061_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_20062_, _20061_, _20060_);
  and (_20063_, _20062_, _02445_);
  or (_20064_, _20063_, _20059_);
  or (_20065_, _20064_, _02459_);
  and (_20066_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and (_20067_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_20068_, _20067_, _20066_);
  and (_20069_, _20068_, _02393_);
  and (_20070_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and (_20071_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_20072_, _20071_, _20070_);
  and (_20073_, _20072_, _02445_);
  or (_20074_, _20073_, _20069_);
  or (_20075_, _20074_, _02421_);
  and (_20076_, _20075_, _02458_);
  and (_20077_, _20076_, _20065_);
  or (_20078_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_20079_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and (_20080_, _20079_, _02445_);
  and (_20081_, _20080_, _20078_);
  or (_20082_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_20083_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and (_20084_, _20083_, _02393_);
  and (_20085_, _20084_, _20082_);
  or (_20086_, _20085_, _20081_);
  or (_20087_, _20086_, _02459_);
  or (_20088_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_20089_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and (_20090_, _20089_, _02445_);
  and (_20091_, _20090_, _20088_);
  or (_20092_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_20093_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and (_20094_, _20093_, _02393_);
  and (_20095_, _20094_, _20092_);
  or (_20096_, _20095_, _20091_);
  or (_20097_, _20096_, _02421_);
  and (_20098_, _20097_, _02414_);
  and (_20099_, _20098_, _20087_);
  or (_20100_, _20099_, _20077_);
  and (_20101_, _20100_, _02496_);
  or (_20102_, _20101_, _20055_);
  and (_20103_, _20102_, _02546_);
  or (_20104_, _20103_, _20008_);
  and (_20105_, _20104_, _02405_);
  or (_20106_, _20105_, _19911_);
  and (_20107_, _20106_, _26777_);
  and (_20108_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and (_20109_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_20110_, _20109_, _20108_);
  and (_20111_, _20110_, _02393_);
  and (_20112_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and (_20113_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_20114_, _20113_, _20112_);
  and (_20115_, _20114_, _02445_);
  or (_20116_, _20115_, _20111_);
  and (_20117_, _20116_, _02421_);
  and (_20118_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and (_20119_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_20120_, _20119_, _20118_);
  and (_20121_, _20120_, _02393_);
  and (_20122_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and (_20123_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_20124_, _20123_, _20122_);
  and (_20125_, _20124_, _02445_);
  or (_20126_, _20125_, _20121_);
  and (_20127_, _20126_, _02459_);
  or (_20128_, _20127_, _20117_);
  and (_20129_, _20128_, _02458_);
  or (_20130_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_20131_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and (_20132_, _20131_, _20130_);
  and (_20133_, _20132_, _02393_);
  or (_20134_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_20135_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and (_20136_, _20135_, _20134_);
  and (_20137_, _20136_, _02445_);
  or (_20138_, _20137_, _20133_);
  and (_20139_, _20138_, _02421_);
  or (_20140_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_20141_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and (_20142_, _20141_, _20140_);
  and (_20143_, _20142_, _02393_);
  or (_20144_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_20145_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and (_20146_, _20145_, _20144_);
  and (_20147_, _20146_, _02445_);
  or (_20148_, _20147_, _20143_);
  and (_20149_, _20148_, _02459_);
  or (_20150_, _20149_, _20139_);
  and (_20151_, _20150_, _02414_);
  or (_20152_, _20151_, _20129_);
  and (_20153_, _20152_, _02398_);
  and (_20154_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_20155_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_20156_, _20155_, _20154_);
  and (_20157_, _20156_, _02393_);
  and (_20158_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_20159_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_20160_, _20159_, _20158_);
  and (_20161_, _20160_, _02445_);
  or (_20162_, _20161_, _20157_);
  and (_20163_, _20162_, _02421_);
  and (_20164_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_20165_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_20166_, _20165_, _20164_);
  and (_20167_, _20166_, _02393_);
  and (_20168_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and (_20169_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_20170_, _20169_, _20168_);
  and (_20171_, _20170_, _02445_);
  or (_20172_, _20171_, _20167_);
  and (_20173_, _20172_, _02459_);
  or (_20174_, _20173_, _20163_);
  and (_20175_, _20174_, _02458_);
  or (_20176_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_20177_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_20178_, _20177_, _02445_);
  and (_20179_, _20178_, _20176_);
  or (_20180_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_20181_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_20182_, _20181_, _02393_);
  and (_20183_, _20182_, _20180_);
  or (_20184_, _20183_, _20179_);
  and (_20185_, _20184_, _02421_);
  or (_20186_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_20187_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_20188_, _20187_, _02445_);
  and (_20189_, _20188_, _20186_);
  or (_20190_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_20191_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_20192_, _20191_, _02393_);
  and (_20193_, _20192_, _20190_);
  or (_20194_, _20193_, _20189_);
  and (_20195_, _20194_, _02459_);
  or (_20196_, _20195_, _20185_);
  and (_20197_, _20196_, _02414_);
  or (_20198_, _20197_, _20175_);
  and (_20199_, _20198_, _02496_);
  or (_20200_, _20199_, _20153_);
  and (_20201_, _20200_, _02400_);
  and (_20202_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and (_20203_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_20204_, _20203_, _20202_);
  and (_20205_, _20204_, _02393_);
  and (_20206_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and (_20207_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_20208_, _20207_, _20206_);
  and (_20209_, _20208_, _02445_);
  or (_20210_, _20209_, _20205_);
  or (_20211_, _20210_, _02459_);
  and (_20212_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and (_20213_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_20214_, _20213_, _20212_);
  and (_20215_, _20214_, _02393_);
  and (_20216_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and (_20217_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_20218_, _20217_, _20216_);
  and (_20219_, _20218_, _02445_);
  or (_20220_, _20219_, _20215_);
  or (_20221_, _20220_, _02421_);
  and (_20222_, _20221_, _02458_);
  and (_20223_, _20222_, _20211_);
  or (_20224_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_20225_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and (_20226_, _20225_, _02445_);
  and (_20227_, _20226_, _20224_);
  or (_20228_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_20229_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and (_20230_, _20229_, _02393_);
  and (_20231_, _20230_, _20228_);
  or (_20232_, _20231_, _20227_);
  or (_20233_, _20232_, _02459_);
  or (_20234_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_20235_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and (_20236_, _20235_, _02445_);
  and (_20237_, _20236_, _20234_);
  or (_20238_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_20239_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and (_20240_, _20239_, _02393_);
  and (_20241_, _20240_, _20238_);
  or (_20242_, _20241_, _20237_);
  or (_20243_, _20242_, _02421_);
  and (_20244_, _20243_, _02414_);
  and (_20245_, _20244_, _20233_);
  or (_20246_, _20245_, _20223_);
  and (_20247_, _20246_, _02496_);
  and (_20248_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and (_20249_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_20250_, _20249_, _20248_);
  and (_20251_, _20250_, _02393_);
  and (_20252_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and (_20253_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_20254_, _20253_, _20252_);
  and (_20255_, _20254_, _02445_);
  or (_20256_, _20255_, _20251_);
  or (_20257_, _20256_, _02459_);
  and (_20258_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and (_20259_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_20260_, _20259_, _20258_);
  and (_20261_, _20260_, _02393_);
  and (_20262_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and (_20263_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_20264_, _20263_, _20262_);
  and (_20265_, _20264_, _02445_);
  or (_20266_, _20265_, _20261_);
  or (_20267_, _20266_, _02421_);
  and (_20268_, _20267_, _02458_);
  and (_20269_, _20268_, _20257_);
  or (_20270_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_20271_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and (_20272_, _20271_, _20270_);
  and (_20273_, _20272_, _02393_);
  or (_20274_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_20275_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and (_20276_, _20275_, _20274_);
  and (_20277_, _20276_, _02445_);
  or (_20278_, _20277_, _20273_);
  or (_20279_, _20278_, _02459_);
  or (_20280_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_20281_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and (_20282_, _20281_, _20280_);
  and (_20283_, _20282_, _02393_);
  or (_20284_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_20285_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and (_20286_, _20285_, _20284_);
  and (_20287_, _20286_, _02445_);
  or (_20288_, _20287_, _20283_);
  or (_20289_, _20288_, _02421_);
  and (_20290_, _20289_, _02414_);
  and (_20291_, _20290_, _20279_);
  or (_20292_, _20291_, _20269_);
  and (_20293_, _20292_, _02398_);
  or (_20294_, _20293_, _20247_);
  and (_20295_, _20294_, _02546_);
  or (_20296_, _20295_, _20201_);
  and (_20297_, _20296_, _02646_);
  or (_20298_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or (_20299_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and (_20300_, _20299_, _02445_);
  and (_20301_, _20300_, _20298_);
  or (_20302_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_20303_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and (_20304_, _20303_, _02393_);
  and (_20305_, _20304_, _20302_);
  or (_20306_, _20305_, _20301_);
  and (_20307_, _20306_, _02459_);
  or (_20308_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_20309_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  and (_20310_, _20309_, _02445_);
  and (_20311_, _20310_, _20308_);
  or (_20312_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or (_20313_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and (_20314_, _20313_, _02393_);
  and (_20315_, _20314_, _20312_);
  or (_20316_, _20315_, _20311_);
  and (_20317_, _20316_, _02421_);
  or (_20318_, _20317_, _20307_);
  and (_20319_, _20318_, _02414_);
  and (_20320_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and (_20321_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_20322_, _20321_, _20320_);
  and (_20323_, _20322_, _02393_);
  and (_20324_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  and (_20325_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_20326_, _20325_, _20324_);
  and (_20327_, _20326_, _02445_);
  or (_20328_, _20327_, _20323_);
  and (_20329_, _20328_, _02459_);
  and (_20330_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  and (_20331_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or (_20332_, _20331_, _20330_);
  and (_20333_, _20332_, _02393_);
  and (_20334_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and (_20335_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or (_20336_, _20335_, _20334_);
  and (_20337_, _20336_, _02445_);
  or (_20338_, _20337_, _20333_);
  and (_20339_, _20338_, _02421_);
  or (_20340_, _20339_, _20329_);
  and (_20341_, _20340_, _02458_);
  or (_20342_, _20341_, _20319_);
  and (_20343_, _20342_, _02496_);
  or (_20344_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_20345_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and (_20346_, _20345_, _20344_);
  and (_20347_, _20346_, _02393_);
  or (_20348_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_20349_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and (_20350_, _20349_, _20348_);
  and (_20351_, _20350_, _02445_);
  or (_20352_, _20351_, _20347_);
  and (_20353_, _20352_, _02459_);
  or (_20354_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_20355_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and (_20356_, _20355_, _20354_);
  and (_20357_, _20356_, _02393_);
  or (_20358_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_20359_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and (_20360_, _20359_, _20358_);
  and (_20361_, _20360_, _02445_);
  or (_20362_, _20361_, _20357_);
  and (_20363_, _20362_, _02421_);
  or (_20364_, _20363_, _20353_);
  and (_20365_, _20364_, _02414_);
  and (_20366_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and (_20367_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_20368_, _20367_, _20366_);
  and (_20369_, _20368_, _02393_);
  and (_20370_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and (_20371_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_20372_, _20371_, _20370_);
  and (_20373_, _20372_, _02445_);
  or (_20374_, _20373_, _20369_);
  and (_20375_, _20374_, _02459_);
  and (_20376_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and (_20377_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_20378_, _20377_, _20376_);
  and (_20379_, _20378_, _02393_);
  and (_20380_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and (_20381_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_20382_, _20381_, _20380_);
  and (_20383_, _20382_, _02445_);
  or (_20384_, _20383_, _20379_);
  and (_20385_, _20384_, _02421_);
  or (_20386_, _20385_, _20375_);
  and (_20387_, _20386_, _02458_);
  or (_20388_, _20387_, _20365_);
  and (_20389_, _20388_, _02398_);
  or (_20390_, _20389_, _20343_);
  and (_20391_, _20390_, _02400_);
  and (_20392_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and (_20393_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_20394_, _20393_, _20392_);
  and (_20395_, _20394_, _02393_);
  and (_20396_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and (_20397_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_20398_, _20397_, _20396_);
  and (_20399_, _20398_, _02445_);
  or (_20400_, _20399_, _20395_);
  or (_20401_, _20400_, _02459_);
  and (_20402_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and (_20403_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_20404_, _20403_, _20402_);
  and (_20405_, _20404_, _02393_);
  and (_20406_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and (_20407_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_20408_, _20407_, _20406_);
  and (_20409_, _20408_, _02445_);
  or (_20410_, _20409_, _20405_);
  or (_20411_, _20410_, _02421_);
  and (_20412_, _20411_, _02458_);
  and (_20413_, _20412_, _20401_);
  or (_20414_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_20415_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and (_20416_, _20415_, _20414_);
  and (_20417_, _20416_, _02393_);
  or (_20418_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_20419_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and (_20420_, _20419_, _20418_);
  and (_20421_, _20420_, _02445_);
  or (_20422_, _20421_, _20417_);
  or (_20423_, _20422_, _02459_);
  or (_20424_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_20425_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and (_20426_, _20425_, _20424_);
  and (_20427_, _20426_, _02393_);
  or (_20428_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_20429_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and (_20430_, _20429_, _20428_);
  and (_20431_, _20430_, _02445_);
  or (_20432_, _20431_, _20427_);
  or (_20433_, _20432_, _02421_);
  and (_20434_, _20433_, _02414_);
  and (_20435_, _20434_, _20423_);
  or (_20436_, _20435_, _20413_);
  and (_20437_, _20436_, _02398_);
  and (_20438_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and (_20439_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_20440_, _20439_, _20438_);
  and (_20441_, _20440_, _02393_);
  and (_20442_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and (_20443_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_20444_, _20443_, _20442_);
  and (_20445_, _20444_, _02445_);
  or (_20446_, _20445_, _20441_);
  or (_20447_, _20446_, _02459_);
  and (_20448_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and (_20449_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_20450_, _20449_, _20448_);
  and (_20451_, _20450_, _02393_);
  and (_20452_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and (_20453_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_20454_, _20453_, _20452_);
  and (_20455_, _20454_, _02445_);
  or (_20456_, _20455_, _20451_);
  or (_20457_, _20456_, _02421_);
  and (_20458_, _20457_, _02458_);
  and (_20459_, _20458_, _20447_);
  or (_20460_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_20461_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and (_20462_, _20461_, _02445_);
  and (_20463_, _20462_, _20460_);
  or (_20464_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_20465_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and (_20466_, _20465_, _02393_);
  and (_20467_, _20466_, _20464_);
  or (_20468_, _20467_, _20463_);
  or (_20469_, _20468_, _02459_);
  or (_20470_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_20471_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and (_20472_, _20471_, _02445_);
  and (_20473_, _20472_, _20470_);
  or (_20474_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_20475_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and (_20476_, _20475_, _02393_);
  and (_20477_, _20476_, _20474_);
  or (_20478_, _20477_, _20473_);
  or (_20479_, _20478_, _02421_);
  and (_20480_, _20479_, _02414_);
  and (_20481_, _20480_, _20469_);
  or (_20482_, _20481_, _20459_);
  and (_20483_, _20482_, _02496_);
  or (_20484_, _20483_, _20437_);
  and (_20485_, _20484_, _02546_);
  or (_20486_, _20485_, _20391_);
  and (_20487_, _20486_, _02405_);
  or (_20488_, _20487_, _20297_);
  and (_20489_, _20488_, _02444_);
  or (_20490_, _20489_, _20107_);
  or (_20491_, _20490_, _02443_);
  or (_20492_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_20493_, _20492_, _22762_);
  and (_11797_, _20493_, _20491_);
  and (_20494_, _06615_, _23824_);
  and (_20495_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_11803_, _20495_, _20494_);
  and (_11817_, _00520_, _22762_);
  and (_11828_, _03305_, _24862_);
  and (_11830_, _00422_, _22762_);
  and (_20496_, _06651_, _23707_);
  and (_20497_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  or (_11834_, _20497_, _20496_);
  and (_20498_, _05346_, _23946_);
  and (_20499_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_11849_, _20499_, _20498_);
  and (_20500_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  and (_20501_, _02306_, _23707_);
  or (_11853_, _20501_, _20500_);
  and (_20502_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and (_20503_, _16375_, _23649_);
  or (_11855_, _20503_, _20502_);
  and (_11857_, _00673_, _22762_);
  and (_11859_, _26370_, _22762_);
  and (_20504_, _06552_, _23778_);
  and (_20505_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_11863_, _20505_, _20504_);
  and (_20506_, _02087_, _24050_);
  and (_20507_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_11867_, _20507_, _20506_);
  or (_20508_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand (_20509_, _22770_, _14710_);
  and (_20510_, _20509_, _22762_);
  and (_26883_[15], _20510_, _20508_);
  and (_11872_, _00595_, _22762_);
  and (_20511_, _18217_, _23824_);
  and (_20512_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_11882_, _20512_, _20511_);
  and (_20513_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and (_20514_, _06507_, _23747_);
  or (_11884_, _20514_, _20513_);
  and (_20515_, _07743_, _24050_);
  and (_20516_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or (_27073_, _20516_, _20515_);
  nand (_20517_, _02077_, _23702_);
  and (_20518_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_20519_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_20520_, _20519_, _20518_);
  or (_20521_, _20520_, _02077_);
  and (_20522_, _20521_, _12675_);
  and (_20523_, _20522_, _20517_);
  and (_20524_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_20525_, _20524_, _20523_);
  and (_11891_, _20525_, _22762_);
  and (_20526_, _07743_, _23707_);
  and (_20527_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or (_27074_, _20527_, _20526_);
  and (_20528_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and (_20529_, _17255_, _23824_);
  or (_11911_, _20529_, _20528_);
  and (_20530_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_20531_, _17255_, _23898_);
  or (_11924_, _20531_, _20530_);
  and (_20532_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and (_20533_, _16325_, _24050_);
  or (_11962_, _20533_, _20532_);
  and (_20534_, _08642_, _23898_);
  and (_20535_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  or (_11964_, _20535_, _20534_);
  and (_20536_, _03339_, _23707_);
  and (_20537_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_11998_, _20537_, _20536_);
  and (_20538_, _08642_, _23824_);
  and (_20539_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  or (_12002_, _20539_, _20538_);
  and (_20540_, _24086_, _23824_);
  and (_20541_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_12009_, _20541_, _20540_);
  and (_20542_, _05459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_26914_, _20542_, _05461_);
  and (_20543_, _08642_, _23778_);
  and (_20544_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  or (_27141_, _20544_, _20543_);
  nor (_20545_, _23596_, _26375_);
  and (_20546_, _23596_, _26375_);
  or (_20547_, _20546_, _20545_);
  and (_12022_, _20547_, _22762_);
  or (_20548_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_12024_, _20548_, _05470_);
  and (_12026_, _01169_, _22762_);
  and (_20549_, _06615_, _23898_);
  and (_20550_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_12028_, _20550_, _20549_);
  and (_12035_, _00919_, _22762_);
  and (_12037_, _00428_, _22762_);
  and (_12040_, _01048_, _22762_);
  and (_12042_, _01231_, _22762_);
  and (_12044_, _00334_, _22762_);
  and (_12048_, _01290_, _22762_);
  and (_12050_, _26541_, _22762_);
  and (_12052_, _01107_, _22762_);
  and (_12054_, _04279_, _22762_);
  and (_12056_, _00600_, _22762_);
  and (_12060_, _00511_, _22762_);
  and (_20551_, _05454_, _23747_);
  and (_20552_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_12063_, _20552_, _20551_);
  and (_20553_, _05454_, _23707_);
  and (_20554_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_12066_, _20554_, _20553_);
  and (_20555_, _05429_, _23707_);
  and (_20556_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_12068_, _20556_, _20555_);
  and (_20557_, _05429_, _23946_);
  and (_20558_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_12070_, _20558_, _20557_);
  and (_20559_, _05379_, _23649_);
  and (_20560_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_12072_, _20560_, _20559_);
  and (_12086_, _00679_, _22762_);
  and (_20561_, _08642_, _23649_);
  and (_20562_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  or (_27142_, _20562_, _20561_);
  and (_20563_, _17263_, _24050_);
  and (_20564_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or (_12101_, _20564_, _20563_);
  and (_20565_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  and (_20566_, _05199_, _24050_);
  or (_27232_, _20566_, _20565_);
  and (_20567_, _05319_, _23824_);
  and (_20568_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_12105_, _20568_, _20567_);
  and (_20569_, _05346_, _23707_);
  and (_20571_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_12107_, _20571_, _20569_);
  and (_20572_, _05319_, _24050_);
  and (_20573_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_12109_, _20573_, _20572_);
  and (_20574_, _05298_, _23946_);
  and (_20575_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_12111_, _20575_, _20574_);
  and (_20576_, _02107_, _23898_);
  and (_20577_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  or (_12113_, _20577_, _20576_);
  and (_20578_, _05223_, _24050_);
  and (_20579_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_12116_, _20579_, _20578_);
  and (_20580_, _07536_, _24050_);
  and (_20581_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or (_27114_, _20581_, _20580_);
  and (_20582_, _05119_, _23778_);
  and (_20583_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  or (_12185_, _20583_, _20582_);
  and (_20584_, _05102_, _23649_);
  and (_20585_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_27301_, _20585_, _20584_);
  and (_20586_, _05102_, _23824_);
  and (_20587_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_12224_, _20587_, _20586_);
  and (_20588_, _04832_, _23778_);
  and (_20589_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_12226_, _20589_, _20588_);
  and (_20590_, _04832_, _24050_);
  and (_20591_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_12228_, _20591_, _20590_);
  and (_20592_, _08642_, _23747_);
  and (_20593_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  or (_12230_, _20593_, _20592_);
  and (_20594_, _04832_, _23649_);
  and (_20595_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_12232_, _20595_, _20594_);
  and (_20596_, _04656_, _23649_);
  and (_20597_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_12234_, _20597_, _20596_);
  and (_20598_, _04656_, _23898_);
  and (_20599_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_12237_, _20599_, _20598_);
  and (_20600_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  and (_20601_, _17775_, _23707_);
  or (_12239_, _20601_, _20600_);
  and (_20602_, _02087_, _23649_);
  and (_20603_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_12241_, _20603_, _20602_);
  and (_20604_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  and (_20605_, _17775_, _24050_);
  or (_12243_, _20605_, _20604_);
  and (_20606_, _01759_, _24050_);
  and (_20607_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_12245_, _20607_, _20606_);
  and (_20608_, _25754_, _23707_);
  and (_20609_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or (_12247_, _20609_, _20608_);
  and (_20610_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and (_20611_, _07513_, _23946_);
  or (_12249_, _20611_, _20610_);
  and (_20612_, _25571_, _23946_);
  and (_20613_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_27058_, _20613_, _20612_);
  and (_20614_, _25571_, _23824_);
  and (_20615_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_12252_, _20615_, _20614_);
  and (_20616_, _25488_, _23649_);
  and (_20617_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_12254_, _20617_, _20616_);
  and (_20618_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  and (_20619_, _17775_, _23946_);
  or (_12256_, _20619_, _20618_);
  and (_20620_, _25340_, _23898_);
  and (_20621_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or (_12258_, _20621_, _20620_);
  and (_20622_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and (_20623_, _16325_, _23747_);
  or (_12260_, _20623_, _20622_);
  and (_20624_, _25340_, _23946_);
  and (_20625_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or (_12264_, _20625_, _20624_);
  and (_20626_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  and (_20627_, _17775_, _23824_);
  or (_12266_, _20627_, _20626_);
  and (_20628_, _24358_, _23946_);
  and (_20629_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or (_12268_, _20629_, _20628_);
  and (_20630_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and (_20631_, _16325_, _23824_);
  or (_26967_, _20631_, _20630_);
  and (_20632_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_20633_, _17255_, _23747_);
  or (_12273_, _20633_, _20632_);
  and (_20634_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and (_20635_, _17255_, _23946_);
  or (_12277_, _20635_, _20634_);
  and (_20636_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and (_20637_, _16325_, _23649_);
  or (_12280_, _20637_, _20636_);
  and (_20638_, _08548_, _23649_);
  and (_20639_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or (_12282_, _20639_, _20638_);
  and (_20640_, _06602_, _23824_);
  and (_20641_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  or (_12284_, _20641_, _20640_);
  and (_20642_, _18217_, _23898_);
  and (_20643_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_12288_, _20643_, _20642_);
  and (_12290_, _00984_, _22762_);
  and (_20644_, _17263_, _23707_);
  and (_20645_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  or (_12292_, _20645_, _20644_);
  and (_20646_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and (_20647_, _17255_, _23649_);
  or (_12294_, _20647_, _20646_);
  and (_20648_, _18217_, _23778_);
  and (_20649_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_12477_, _20649_, _20648_);
  and (_20650_, _08548_, _24050_);
  and (_20651_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or (_27137_, _20651_, _20650_);
  and (_20652_, _25739_, _23649_);
  and (_20653_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or (_12509_, _20653_, _20652_);
  and (_20654_, _07743_, _23778_);
  and (_20655_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or (_27071_, _20655_, _20654_);
  and (_20656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_20657_, _20656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_20658_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_20659_, _20658_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_20660_, _20659_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_20661_, _20660_, _20657_);
  and (_20662_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_20663_, _20662_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_20664_, _20663_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_20665_, _20664_, _20661_);
  and (_20666_, _20665_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_20667_, _20666_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_20668_, _20667_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_20669_, _20667_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_20670_, _20669_, _20668_);
  nor (_20671_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20672_, _20671_);
  and (_20673_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _22841_);
  and (_20674_, _20656_, _22854_);
  nor (_20675_, _20656_, _22854_);
  nor (_20676_, _20675_, _20674_);
  nor (_20677_, _20676_, _22841_);
  nor (_20678_, _20677_, _20673_);
  not (_20679_, _20678_);
  nor (_20680_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20681_, _22849_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_20682_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _22845_);
  nor (_20683_, _20682_, _20681_);
  and (_20684_, _20683_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20685_, _20684_, _20680_);
  nor (_20686_, _20685_, _08039_);
  and (_20687_, _20685_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_20688_, _20687_, _20686_);
  nor (_20689_, _20688_, _20679_);
  nor (_20690_, _20685_, _07621_);
  and (_20691_, _20685_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_20692_, _20691_, _20690_);
  nor (_20693_, _20692_, _20678_);
  nor (_20694_, _20693_, _20689_);
  nor (_20695_, _20694_, _20672_);
  and (_20696_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _22841_);
  not (_20697_, _20696_);
  nor (_20698_, _20685_, _07600_);
  and (_20699_, _20685_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_20700_, _20699_, _20698_);
  nor (_20701_, _20700_, _20679_);
  not (_20702_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_20703_, _20685_, _20702_);
  and (_20704_, _20685_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_20705_, _20704_, _20703_);
  nor (_20706_, _20705_, _20678_);
  nor (_20707_, _20706_, _20701_);
  nor (_20708_, _20707_, _20697_);
  nor (_20709_, _20708_, _20695_);
  and (_20710_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20711_, _20710_);
  not (_20712_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_20713_, _20685_, _20712_);
  and (_20714_, _20685_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_20715_, _20714_, _20713_);
  nor (_20716_, _20715_, _20679_);
  nor (_20717_, _20685_, _07665_);
  and (_20718_, _20685_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_20719_, _20718_, _20717_);
  nor (_20720_, _20719_, _20678_);
  nor (_20721_, _20720_, _20716_);
  nor (_20722_, _20721_, _20711_);
  and (_20723_, _22845_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20724_, _20723_);
  nor (_20725_, _20685_, _07657_);
  and (_20726_, _20685_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_20727_, _20726_, _20725_);
  nor (_20728_, _20727_, _20679_);
  nor (_20729_, _20685_, _08225_);
  and (_20730_, _20685_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_20731_, _20730_, _20729_);
  nor (_20732_, _20731_, _20678_);
  nor (_20733_, _20732_, _20728_);
  nor (_20734_, _20733_, _20724_);
  nor (_20735_, _20734_, _20722_);
  and (_20736_, _20735_, _20709_);
  not (_20737_, _20685_);
  and (_20738_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_20739_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_20740_, _20739_, _20738_);
  and (_20741_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_20742_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_20743_, _20742_, _20741_);
  and (_20744_, _20743_, _20740_);
  and (_20745_, _20744_, _20737_);
  and (_20746_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_20747_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_20748_, _20747_, _20746_);
  and (_20749_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_20750_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_20751_, _20750_, _20749_);
  and (_20752_, _20751_, _20748_);
  and (_20753_, _20752_, _20685_);
  or (_20754_, _20753_, _20679_);
  nor (_20755_, _20754_, _20745_);
  and (_20756_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_20757_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_20758_, _20757_, _20756_);
  and (_20759_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_20760_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_20761_, _20760_, _20759_);
  and (_20762_, _20761_, _20758_);
  nor (_20763_, _20762_, _20685_);
  and (_20764_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_20765_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_20766_, _20765_, _20764_);
  and (_20767_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_20768_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_20769_, _20768_, _20767_);
  and (_20770_, _20769_, _20766_);
  nor (_20771_, _20770_, _20737_);
  or (_20772_, _20771_, _20763_);
  and (_20773_, _20772_, _20679_);
  nor (_20774_, _20773_, _20755_);
  nor (_20775_, _20774_, _20736_);
  and (_20776_, _20775_, _20670_);
  nor (_20777_, _20666_, _22897_);
  and (_20778_, _20663_, _20661_);
  and (_20779_, _20778_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_20780_, _20779_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_20781_, _20780_, _22897_);
  nor (_20782_, _20781_, _20777_);
  not (_20783_, _20782_);
  and (_20784_, _20783_, _20775_);
  nor (_20785_, _20665_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_20786_, _20785_, _20666_);
  and (_20787_, _20786_, _20775_);
  nor (_20788_, _20783_, _20775_);
  nor (_20789_, _20788_, _20784_);
  nor (_20790_, _20778_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_20791_, _20790_, _20779_);
  and (_20792_, _20791_, _20775_);
  nor (_20793_, _20791_, _20775_);
  and (_20794_, _20662_, _20661_);
  nor (_20795_, _20794_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_20796_, _20795_, _20778_);
  and (_20797_, _20796_, _20775_);
  nor (_20798_, _20796_, _20775_);
  nor (_20799_, _20798_, _20797_);
  and (_20800_, _20661_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_20801_, _20800_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_20802_, _20801_, _20794_);
  and (_20803_, _20802_, _20775_);
  nor (_20804_, _20802_, _20775_);
  nor (_20805_, _20661_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_20806_, _20805_, _20800_);
  and (_20807_, _20806_, _20775_);
  and (_20808_, _20659_, _20657_);
  nor (_20809_, _20808_, _22874_);
  and (_20810_, _20808_, _22874_);
  nor (_20811_, _20810_, _20809_);
  not (_20812_, _20811_);
  and (_20813_, _20812_, _20775_);
  nor (_20814_, _20812_, _20775_);
  and (_20815_, _20658_, _20657_);
  nor (_20816_, _20815_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_20817_, _20816_, _20808_);
  and (_20818_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_20819_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_20820_, _20819_, _20818_);
  and (_20821_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_20822_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_20823_, _20822_, _20821_);
  and (_20824_, _20823_, _20820_);
  and (_20825_, _20824_, _20685_);
  and (_20826_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_20827_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_20828_, _20827_, _20826_);
  and (_20829_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_20830_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_20831_, _20830_, _20829_);
  and (_20832_, _20831_, _20828_);
  and (_20833_, _20832_, _20737_);
  or (_20834_, _20833_, _20679_);
  nor (_20835_, _20834_, _20825_);
  and (_20836_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_20837_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_20838_, _20837_, _20836_);
  and (_20839_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_20840_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_20841_, _20840_, _20839_);
  and (_20842_, _20841_, _20838_);
  nor (_20843_, _20842_, _20685_);
  and (_20844_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_20845_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_20846_, _20845_, _20844_);
  and (_20847_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_20848_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_20849_, _20848_, _20847_);
  and (_20850_, _20849_, _20846_);
  nor (_20851_, _20850_, _20737_);
  or (_20852_, _20851_, _20843_);
  and (_20853_, _20852_, _20679_);
  nor (_20854_, _20853_, _20835_);
  nor (_20855_, _20854_, _20736_);
  and (_20856_, _20855_, _20817_);
  nor (_20857_, _20855_, _20817_);
  nor (_20858_, _20857_, _20856_);
  not (_20859_, _20858_);
  and (_20860_, _20657_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_20861_, _20860_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_20862_, _20861_, _20815_);
  and (_20863_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_20864_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_20865_, _20864_, _20863_);
  and (_20866_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_20867_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_20868_, _20867_, _20866_);
  and (_20869_, _20868_, _20865_);
  and (_20870_, _20869_, _20737_);
  and (_20871_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_20872_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_20873_, _20872_, _20871_);
  and (_20874_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_20875_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_20876_, _20875_, _20874_);
  and (_20877_, _20876_, _20873_);
  and (_20878_, _20877_, _20685_);
  or (_20879_, _20878_, _20679_);
  nor (_20880_, _20879_, _20870_);
  and (_20881_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_20882_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_20883_, _20882_, _20881_);
  and (_20884_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_20885_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_20886_, _20885_, _20884_);
  and (_20887_, _20886_, _20883_);
  and (_20888_, _20887_, _20737_);
  and (_20889_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_20890_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_20891_, _20890_, _20889_);
  and (_20892_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_20893_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_20894_, _20893_, _20892_);
  and (_20895_, _20894_, _20891_);
  and (_20896_, _20895_, _20685_);
  nor (_20897_, _20896_, _20888_);
  and (_20898_, _20897_, _20679_);
  nor (_20899_, _20898_, _20880_);
  nor (_20900_, _20899_, _20736_);
  and (_20901_, _20900_, _20862_);
  nor (_20902_, _20900_, _20862_);
  nor (_20903_, _20902_, _20901_);
  not (_20904_, _20903_);
  and (_20905_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_20906_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_20907_, _20906_, _20905_);
  and (_20908_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_20909_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_20910_, _20909_, _20908_);
  and (_20911_, _20910_, _20907_);
  and (_20912_, _20911_, _20737_);
  and (_20913_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_20914_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_20915_, _20914_, _20913_);
  and (_20916_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_20917_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_20918_, _20917_, _20916_);
  and (_20919_, _20918_, _20915_);
  and (_20920_, _20919_, _20685_);
  or (_20921_, _20920_, _20679_);
  nor (_20922_, _20921_, _20912_);
  and (_20923_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_20924_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_20925_, _20924_, _20923_);
  and (_20926_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_20927_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_20928_, _20927_, _20926_);
  and (_20929_, _20928_, _20925_);
  nor (_20930_, _20929_, _20685_);
  and (_20931_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_20932_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_20933_, _20932_, _20931_);
  and (_20934_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_20935_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_20936_, _20935_, _20934_);
  and (_20937_, _20936_, _20933_);
  nor (_20938_, _20937_, _20737_);
  or (_20939_, _20938_, _20930_);
  and (_20940_, _20939_, _20679_);
  nor (_20941_, _20940_, _20922_);
  nor (_20942_, _20941_, _20736_);
  nor (_20943_, _20657_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_20944_, _20943_, _20860_);
  and (_20945_, _20944_, _20942_);
  not (_20946_, _20676_);
  and (_20947_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_20948_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_20949_, _20948_, _20947_);
  and (_20950_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_20951_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_20952_, _20951_, _20950_);
  and (_20953_, _20952_, _20949_);
  and (_20954_, _20953_, _20737_);
  and (_20955_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_20956_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_20957_, _20956_, _20955_);
  and (_20958_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_20959_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_20960_, _20959_, _20958_);
  and (_20961_, _20960_, _20957_);
  and (_20962_, _20961_, _20685_);
  or (_20963_, _20962_, _20679_);
  nor (_20964_, _20963_, _20954_);
  and (_20965_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_20966_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_20967_, _20966_, _20965_);
  and (_20968_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_20969_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_20970_, _20969_, _20968_);
  and (_20971_, _20970_, _20967_);
  nor (_20972_, _20971_, _20685_);
  and (_20973_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_20974_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_20975_, _20974_, _20973_);
  and (_20976_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_20977_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_20978_, _20977_, _20976_);
  and (_20979_, _20978_, _20975_);
  nor (_20980_, _20979_, _20737_);
  or (_20981_, _20980_, _20972_);
  and (_20982_, _20981_, _20679_);
  nor (_20983_, _20982_, _20964_);
  nor (_20984_, _20983_, _20736_);
  and (_20985_, _20984_, _20946_);
  nor (_20986_, _20984_, _20946_);
  nor (_20987_, _20986_, _20985_);
  not (_20988_, _20987_);
  not (_20989_, _20683_);
  and (_20990_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_20991_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_20992_, _20991_, _20990_);
  and (_20993_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_20994_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_20995_, _20994_, _20993_);
  and (_20996_, _20995_, _20992_);
  and (_20997_, _20996_, _20737_);
  and (_20998_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_20999_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_21000_, _20999_, _20998_);
  and (_21001_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_21002_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_21003_, _21002_, _21001_);
  and (_21004_, _21003_, _21000_);
  and (_21005_, _21004_, _20685_);
  or (_21006_, _21005_, _20679_);
  nor (_21007_, _21006_, _20997_);
  and (_21008_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_21009_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_21010_, _21009_, _21008_);
  and (_21011_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_21012_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_21013_, _21012_, _21011_);
  and (_21014_, _21013_, _21010_);
  and (_21015_, _21014_, _20737_);
  and (_21016_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_21017_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_21018_, _21017_, _21016_);
  and (_21019_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_21020_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_21021_, _21020_, _21019_);
  and (_21022_, _21021_, _21018_);
  and (_21023_, _21022_, _20685_);
  nor (_21024_, _21023_, _21015_);
  and (_21025_, _21024_, _20679_);
  nor (_21026_, _21025_, _21007_);
  nor (_21027_, _21026_, _20736_);
  and (_21028_, _21027_, _20989_);
  and (_21029_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_21030_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_21031_, _21030_, _21029_);
  and (_21032_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_21033_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_21034_, _21033_, _21032_);
  and (_21035_, _21034_, _21031_);
  and (_21036_, _21035_, _20737_);
  and (_21037_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_21038_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_21039_, _21038_, _21037_);
  and (_21040_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_21041_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_21042_, _21041_, _21040_);
  and (_21043_, _21042_, _21039_);
  and (_21044_, _21043_, _20685_);
  or (_21045_, _21044_, _20679_);
  nor (_21046_, _21045_, _21036_);
  and (_21047_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_21048_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_21049_, _21048_, _21047_);
  and (_21050_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_21051_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_21052_, _21051_, _21050_);
  and (_21053_, _21052_, _21049_);
  nor (_21054_, _21053_, _20685_);
  and (_21055_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_21056_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_21057_, _21056_, _21055_);
  and (_21058_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_21059_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_21060_, _21059_, _21058_);
  and (_21061_, _21060_, _21057_);
  nor (_21062_, _21061_, _20737_);
  or (_21063_, _21062_, _21054_);
  and (_21064_, _21063_, _20679_);
  nor (_21065_, _21064_, _21046_);
  nor (_21066_, _21065_, _20736_);
  and (_21067_, _21066_, _22845_);
  and (_21068_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_21069_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_21070_, _21069_, _21068_);
  and (_21071_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_21072_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_21073_, _21072_, _21071_);
  and (_21074_, _21073_, _21070_);
  and (_21075_, _21074_, _20737_);
  and (_21076_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_21077_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_21078_, _21077_, _21076_);
  and (_21079_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_21080_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_21081_, _21080_, _21079_);
  and (_21082_, _21081_, _21078_);
  and (_21083_, _21082_, _20685_);
  or (_21084_, _21083_, _20679_);
  nor (_21085_, _21084_, _21075_);
  and (_21086_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_21087_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_21088_, _21087_, _21086_);
  and (_21089_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_21090_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_21091_, _21090_, _21089_);
  and (_21092_, _21091_, _21088_);
  and (_21093_, _21092_, _20737_);
  and (_21094_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_21095_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_21096_, _21095_, _21094_);
  and (_21097_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_21098_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_21099_, _21098_, _21097_);
  and (_21100_, _21099_, _21096_);
  and (_21101_, _21100_, _20685_);
  nor (_21102_, _21101_, _21093_);
  and (_21103_, _21102_, _20679_);
  nor (_21104_, _21103_, _21085_);
  nor (_21105_, _21104_, _20736_);
  and (_21106_, _21105_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21107_, _21066_, _22845_);
  nor (_21108_, _21107_, _21067_);
  and (_21109_, _21108_, _21106_);
  nor (_21110_, _21109_, _21067_);
  nor (_21111_, _21027_, _20989_);
  nor (_21112_, _21111_, _21028_);
  not (_21113_, _21112_);
  nor (_21114_, _21113_, _21110_);
  nor (_21115_, _21114_, _21028_);
  nor (_21116_, _21115_, _20988_);
  nor (_21117_, _21116_, _20985_);
  nor (_21118_, _20944_, _20942_);
  nor (_21119_, _21118_, _20945_);
  not (_21120_, _21119_);
  nor (_21121_, _21120_, _21117_);
  nor (_21122_, _21121_, _20945_);
  nor (_21123_, _21122_, _20904_);
  nor (_21124_, _21123_, _20901_);
  nor (_21125_, _21124_, _20859_);
  nor (_21126_, _21125_, _20856_);
  nor (_21127_, _21126_, _20814_);
  or (_21128_, _21127_, _20813_);
  nor (_21129_, _20806_, _20775_);
  nor (_21130_, _21129_, _20807_);
  and (_21131_, _21130_, _21128_);
  nor (_21132_, _21131_, _20807_);
  nor (_21133_, _21132_, _20804_);
  or (_21134_, _21133_, _20803_);
  and (_21135_, _21134_, _20799_);
  nor (_21136_, _21135_, _20797_);
  nor (_21137_, _21136_, _20793_);
  or (_21138_, _21137_, _20792_);
  nor (_21139_, _20786_, _20775_);
  nor (_21140_, _21139_, _20787_);
  and (_21141_, _21140_, _21138_);
  and (_21142_, _21141_, _20789_);
  or (_21143_, _21142_, _20787_);
  nor (_21144_, _21143_, _20784_);
  nor (_21145_, _20775_, _20670_);
  nor (_21146_, _21145_, _20776_);
  not (_21147_, _21146_);
  nor (_21148_, _21147_, _21144_);
  nor (_21149_, _21148_, _20776_);
  nor (_21150_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_21151_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_21152_, _21151_, _21150_);
  not (_21153_, _21152_);
  nor (_21154_, _21153_, _20669_);
  and (_21155_, _21153_, _20669_);
  nor (_21156_, _21155_, _21154_);
  not (_21157_, _21156_);
  and (_21158_, _21157_, _20775_);
  nor (_21159_, _21157_, _20775_);
  nor (_21160_, _21159_, _21158_);
  not (_21161_, _21160_);
  nand (_21162_, _21161_, _21149_);
  or (_21163_, _21161_, _21149_);
  and (_21164_, _21163_, _21162_);
  and (_21165_, _21147_, _21144_);
  nor (_21166_, _21165_, _21148_);
  nor (_21167_, _21166_, _22837_);
  and (_21168_, _21166_, _22837_);
  nor (_21169_, _21141_, _20787_);
  and (_21170_, _20789_, _22832_);
  nor (_21171_, _20789_, _22832_);
  nor (_21172_, _21171_, _21170_);
  nand (_21173_, _21172_, _21169_);
  or (_21174_, _21172_, _21169_);
  and (_21175_, _21174_, _21173_);
  nor (_21176_, _21140_, _21138_);
  nor (_21177_, _21176_, _21141_);
  nor (_21178_, _21177_, _22827_);
  and (_21179_, _21177_, _22827_);
  nor (_21180_, _20791_, _22823_);
  and (_21181_, _20791_, _22823_);
  or (_21182_, _21181_, _21180_);
  nand (_21183_, _21182_, _20775_);
  or (_21184_, _21182_, _20775_);
  and (_21185_, _21184_, _21183_);
  not (_21186_, _21185_);
  nand (_21187_, _21186_, _21136_);
  or (_21188_, _21186_, _21136_);
  and (_21189_, _21188_, _21187_);
  nor (_21190_, _21134_, _20799_);
  nor (_21191_, _21190_, _21135_);
  nor (_21192_, _21191_, _22819_);
  and (_21193_, _21191_, _22819_);
  not (_21194_, _20775_);
  nor (_21195_, _20802_, _22814_);
  and (_21196_, _20802_, _22814_);
  or (_21197_, _21196_, _21195_);
  nand (_21198_, _21197_, _21194_);
  or (_21199_, _21197_, _21194_);
  and (_21200_, _21199_, _21198_);
  or (_21201_, _21200_, _21132_);
  nand (_21202_, _21200_, _21132_);
  and (_21203_, _21202_, _21201_);
  nor (_21204_, _20813_, _20814_);
  nor (_21205_, _21204_, _21126_);
  and (_21206_, _21204_, _21126_);
  or (_21207_, _21206_, _21205_);
  nor (_21208_, _21207_, _22806_);
  and (_21209_, _21207_, _22806_);
  and (_21210_, _21124_, _20859_);
  nor (_21211_, _21210_, _21125_);
  and (_21212_, _21211_, _22802_);
  nor (_21213_, _21211_, _22802_);
  and (_21214_, _21122_, _20904_);
  nor (_21215_, _21214_, _21123_);
  nor (_21216_, _21215_, _22798_);
  and (_21217_, _21215_, _22798_);
  and (_21218_, _21120_, _21117_);
  nor (_21219_, _21218_, _21121_);
  and (_21220_, _21219_, _22794_);
  and (_21221_, _21115_, _20988_);
  nor (_21222_, _21221_, _21116_);
  and (_21223_, _21222_, _22788_);
  nor (_21224_, _21222_, _22788_);
  and (_21225_, _21113_, _21110_);
  nor (_21226_, _21225_, _21114_);
  nor (_21227_, _21226_, _22783_);
  nor (_21228_, _21108_, _21106_);
  nor (_21229_, _21228_, _21109_);
  nor (_21230_, _21229_, _22778_);
  and (_21231_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21232_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_21233_, _21232_, _21231_);
  and (_21234_, _21233_, _21105_);
  nor (_21235_, _21233_, _21105_);
  or (_21236_, _21235_, _21234_);
  and (_21237_, _21229_, _22778_);
  or (_21238_, _21237_, _21236_);
  or (_21239_, _21238_, _21230_);
  and (_21240_, _21226_, _22783_);
  or (_21241_, _21240_, _21239_);
  or (_21242_, _21241_, _21227_);
  or (_21243_, _21242_, _21224_);
  or (_21244_, _21243_, _21223_);
  nor (_21245_, _21219_, _22794_);
  or (_21246_, _21245_, _21244_);
  or (_21248_, _21246_, _21220_);
  or (_21249_, _21248_, _21217_);
  or (_21250_, _21249_, _21216_);
  or (_21251_, _21250_, _21213_);
  or (_21252_, _21251_, _21212_);
  or (_21253_, _21252_, _21209_);
  or (_21254_, _21253_, _21208_);
  nor (_21255_, _21130_, _21128_);
  nor (_21256_, _21255_, _21131_);
  nor (_21257_, _21256_, _22810_);
  and (_21258_, _21256_, _22810_);
  or (_21259_, _21258_, _21257_);
  or (_21260_, _21259_, _21254_);
  or (_21261_, _21260_, _21203_);
  or (_21262_, _21261_, _21193_);
  or (_21263_, _21262_, _21192_);
  or (_21264_, _21263_, _21189_);
  or (_21265_, _21264_, _21179_);
  or (_21266_, _21265_, _21178_);
  or (_21267_, _21266_, _21175_);
  or (_21268_, _21267_, _21168_);
  or (_21269_, _21268_, _21167_);
  or (_21270_, _21269_, _21164_);
  and (_21271_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21272_, _21271_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_21273_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21274_, _21273_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_21275_, _21274_, _21272_);
  not (_21276_, _21275_);
  nor (_21277_, _21272_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21278_, _21272_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21279_, _21278_, _21277_);
  nand (_21280_, _21279_, _20702_);
  or (_21281_, _21279_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_21282_, _21281_, _21280_);
  and (_21283_, _21282_, _21276_);
  nand (_21284_, _21279_, _07612_);
  or (_21285_, _21279_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_21286_, _21285_, _21275_);
  and (_21287_, _21286_, _21284_);
  or (_21288_, _21287_, _21283_);
  or (_21289_, _21288_, _22778_);
  and (_21290_, _22783_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21291_, \oc8051_symbolic_cxrom1.regvalid [5], _22788_);
  and (_21292_, \oc8051_symbolic_cxrom1.regvalid [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21293_, _21292_, _21291_);
  and (_21294_, _21293_, _21290_);
  or (_21295_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21296_, \oc8051_symbolic_cxrom1.regvalid [1], _22788_);
  and (_21297_, _21296_, _21271_);
  and (_21298_, _21297_, _21295_);
  or (_21299_, _21298_, _21294_);
  nor (_21300_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21301_, _21300_, _22783_);
  nor (_21302_, _21301_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21303_, _21301_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21304_, _21303_, _21302_);
  and (_21305_, _21304_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_21306_, _21300_, _22783_);
  nor (_21307_, _21306_, _21301_);
  or (_21308_, _08145_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_21309_, _21308_, _21307_);
  or (_21310_, _21309_, _21305_);
  and (_21311_, _21310_, _22778_);
  nor (_21312_, _21304_, _07600_);
  and (_21313_, _21304_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_21314_, _21313_, _21312_);
  or (_21315_, _21314_, _21307_);
  and (_21316_, _21315_, _21311_);
  or (_21317_, _21316_, _21299_);
  and (_21318_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21319_, \oc8051_symbolic_cxrom1.regvalid [0], _22788_);
  or (_21320_, _21319_, _21318_);
  and (_21321_, _21320_, _22783_);
  and (_21322_, \oc8051_symbolic_cxrom1.regvalid [4], _22788_);
  and (_21323_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21324_, _21323_, _21322_);
  and (_21325_, _21324_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_21326_, _21325_, _21321_);
  or (_21327_, _21326_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21328_, _21290_, _21324_);
  or (_21329_, \oc8051_symbolic_cxrom1.regvalid [0], _22788_);
  or (_21330_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21331_, _21330_, _21271_);
  and (_21332_, _21331_, _21329_);
  or (_21333_, _21332_, _21328_);
  and (_21334_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21335_, \oc8051_symbolic_cxrom1.regvalid [6], _22788_);
  or (_21336_, _21335_, _22783_);
  or (_21337_, _21336_, _21334_);
  or (_21338_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21339_, \oc8051_symbolic_cxrom1.regvalid [10], _22788_);
  and (_21340_, _21339_, _21338_);
  or (_21341_, _21340_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21342_, _21341_, _21337_);
  and (_21343_, _21342_, _22778_);
  or (_21344_, _21343_, _21333_);
  or (_21345_, _21342_, _22778_);
  and (_21346_, _21345_, _22772_);
  and (_21347_, _21346_, _21344_);
  and (_21349_, _21347_, _21327_);
  nand (_21350_, _21279_, _07621_);
  or (_21351_, _21279_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_21352_, _21351_, _21350_);
  and (_21353_, _21352_, _21276_);
  nand (_21354_, _21279_, _07572_);
  or (_21355_, _21279_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_21356_, _21355_, _21275_);
  and (_21357_, _21356_, _21354_);
  or (_21358_, _21357_, _21353_);
  or (_21359_, _21358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21360_, _21359_, _21349_);
  and (_21361_, _21360_, _21317_);
  and (_21362_, _21361_, _21289_);
  or (_21363_, \oc8051_symbolic_cxrom1.regvalid [10], _22778_);
  or (_21364_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_21365_, _21364_, _21363_);
  nand (_21366_, _21365_, _21304_);
  or (_21367_, \oc8051_symbolic_cxrom1.regvalid [2], _22778_);
  or (_21368_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21369_, _21368_, _21367_);
  or (_21370_, _21369_, _21304_);
  and (_21371_, _21370_, _21366_);
  or (_21372_, _21371_, _21307_);
  nor (_21373_, _21279_, _20712_);
  and (_21374_, _21279_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_21375_, _21374_, _21373_);
  and (_21376_, _21375_, _21276_);
  or (_21377_, _21279_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_21378_, \oc8051_symbolic_cxrom1.regvalid [12], _22788_);
  and (_21379_, _21378_, _21275_);
  and (_21380_, _21379_, _21377_);
  or (_21381_, _21380_, _22778_);
  or (_21382_, _21381_, _21376_);
  nand (_21383_, \oc8051_symbolic_cxrom1.regvalid [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_21384_, _21383_, _21308_);
  or (_21385_, _21384_, _22783_);
  or (_21386_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21387_, \oc8051_symbolic_cxrom1.regvalid [11], _22788_);
  and (_21388_, _21387_, _21386_);
  or (_21389_, _21388_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21390_, _21389_, _21385_);
  and (_21391_, _21390_, _21273_);
  and (_21392_, _22778_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_21393_, _21293_, _22783_);
  or (_21394_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21395_, \oc8051_symbolic_cxrom1.regvalid [9], _22788_);
  and (_21396_, _21395_, _21394_);
  or (_21397_, _21396_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21398_, _21397_, _21393_);
  and (_21399_, _21398_, _21392_);
  or (_21400_, _21399_, _21391_);
  and (_21401_, _21390_, _22778_);
  or (_21402_, _21401_, _21299_);
  and (_21403_, _21402_, _21400_);
  and (_21404_, _21403_, _21382_);
  and (_21405_, _21404_, _21372_);
  or (_21406_, _21279_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_21407_, \oc8051_symbolic_cxrom1.regvalid [14], _22788_);
  and (_21408_, _21407_, _21406_);
  or (_21409_, _21408_, _21276_);
  nand (_21410_, _21279_, _08225_);
  or (_21411_, _21279_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_21412_, _21411_, _21410_);
  or (_21413_, _21412_, _21275_);
  and (_21414_, _21413_, _21409_);
  or (_21415_, _21414_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21416_, _21304_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_21417_, _21335_, _22778_);
  or (_21418_, _21417_, _21416_);
  and (_21420_, _21304_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_21421_, _21322_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_21422_, _21421_, _21420_);
  nand (_21423_, _21422_, _21418_);
  nand (_21424_, _21423_, _21307_);
  and (_21425_, _21424_, _21415_);
  and (_21426_, _21425_, _21405_);
  or (_21427_, _21426_, _21362_);
  nor (_21428_, _20671_, _22849_);
  and (_21429_, _20680_, _22845_);
  nor (_21430_, _21429_, _21428_);
  not (_21431_, _21430_);
  and (_21432_, _21428_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21433_, _21428_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21434_, _21433_, _21432_);
  and (_21435_, _21434_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_21436_, _21434_, _07600_);
  or (_21437_, _21436_, _21435_);
  and (_21438_, _21437_, _21431_);
  nand (_21439_, _21434_, _07612_);
  nor (_21440_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21441_, _21440_, _21431_);
  and (_21442_, _21441_, _21439_);
  or (_21443_, _21442_, _21438_);
  and (_21444_, _21443_, _20671_);
  and (_21445_, _21434_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_21446_, _21434_, _20712_);
  or (_21447_, _21446_, _21445_);
  and (_21448_, _21447_, _21431_);
  or (_21449_, _21434_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_21450_, \oc8051_symbolic_cxrom1.regvalid [12], _22854_);
  nor (_21451_, _21450_, _21431_);
  and (_21452_, _21451_, _21449_);
  or (_21453_, _21452_, _21448_);
  and (_21454_, _21453_, _20723_);
  or (_21455_, _21454_, _21444_);
  and (_21456_, _21434_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_21457_, _21434_, _07657_);
  or (_21458_, _21457_, _21456_);
  and (_21459_, _21458_, _21431_);
  or (_21460_, _21434_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_21461_, _07637_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21462_, _21461_, _21431_);
  and (_21463_, _21462_, _21460_);
  or (_21464_, _21463_, _21459_);
  and (_21465_, _21464_, _20710_);
  and (_21466_, _21434_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_21467_, _21434_, _08039_);
  or (_21468_, _21467_, _21466_);
  and (_21469_, _21468_, _21431_);
  nand (_21470_, _21434_, _07572_);
  nor (_21471_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21472_, _21471_, _21431_);
  and (_21473_, _21472_, _21470_);
  or (_21474_, _21473_, _21469_);
  and (_21475_, _21474_, _20696_);
  or (_21476_, _21475_, _21465_);
  or (_21477_, _21476_, _21455_);
  and (_21478_, _07612_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21479_, _21478_);
  nor (_21480_, _21440_, _22849_);
  and (_21481_, _21480_, _21479_);
  and (_21482_, _20702_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21483_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21484_, _21483_, _21482_);
  and (_21485_, _21484_, _22849_);
  nor (_21486_, _21485_, _21481_);
  nor (_21487_, _21486_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_21488_, _07572_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21489_, _21488_, _21471_);
  and (_21490_, _21489_, _20681_);
  and (_21491_, _08039_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21492_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21493_, _21492_, _22849_);
  nor (_21494_, _21493_, _21491_);
  and (_21495_, _21494_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_21496_, _21495_, _21490_);
  not (_21497_, _21496_);
  nor (_21498_, _21497_, _21487_);
  nor (_21499_, _21498_, _22841_);
  not (_21500_, _21499_);
  nor (_21501_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21502_, _21501_);
  nor (_21503_, _21461_, _22849_);
  and (_21504_, _21503_, _21502_);
  and (_21505_, _08225_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21506_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21507_, _21506_, _21505_);
  and (_21508_, _21507_, _22849_);
  nor (_21509_, _21508_, _21504_);
  nor (_21510_, _21509_, _20672_);
  and (_21511_, _20696_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_21512_, _20712_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21513_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21514_, _21513_, _21512_);
  and (_21515_, _21514_, _21511_);
  nor (_21516_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21517_, _21516_, _21450_);
  and (_21518_, _20681_, _22841_);
  and (_21519_, _21518_, _21517_);
  nor (_21520_, _21519_, _21515_);
  not (_21521_, _21520_);
  nor (_21522_, _21521_, _21510_);
  and (_21523_, _21522_, _21500_);
  and (_21524_, _21489_, _20682_);
  nor (_21525_, _21524_, _22841_);
  nor (_21526_, _21486_, _22845_);
  nor (_21527_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_21528_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_21529_, _07621_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21530_, _21529_, _21528_);
  and (_21531_, _21530_, _21527_);
  nor (_21532_, _21531_, _21526_);
  and (_21533_, _21532_, _21525_);
  nor (_21534_, _21509_, _22845_);
  nor (_21535_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_21536_, _07665_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21537_, _21536_, _21535_);
  and (_21538_, _21537_, _21527_);
  and (_21539_, _21517_, _20682_);
  or (_21540_, _21539_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_21541_, _21540_, _21538_);
  nor (_21542_, _21541_, _21534_);
  nor (_21543_, _21542_, _21533_);
  not (_21544_, _22770_);
  nor (_21545_, _21544_, first_instr);
  nand (_21546_, _21545_, _21543_);
  nor (_21547_, _21546_, _21523_);
  nand (_21548_, _21547_, _21477_);
  nor (_21549_, _21548_, _20736_);
  and (_21550_, _21549_, _21427_);
  nor (_21551_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21552_, _08575_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21553_, _21552_, _21551_);
  and (_21554_, _21553_, _21527_);
  nor (_21555_, _21554_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21556_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21557_, _09098_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21558_, _21557_, _21556_);
  and (_21559_, _21558_, _20682_);
  not (_21560_, _21559_);
  nor (_21561_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21562_, _08830_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21563_, _21562_, _21561_);
  and (_21564_, _21563_, _20681_);
  nor (_21565_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21566_, _09352_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21567_, _21566_, _21565_);
  and (_21568_, _21567_, _20656_);
  nor (_21569_, _21568_, _21564_);
  and (_21570_, _21569_, _21560_);
  and (_21571_, _21570_, _21555_);
  nor (_21572_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21573_, _09586_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21574_, _21573_, _21572_);
  and (_21575_, _21574_, _21527_);
  nor (_21576_, _21575_, _22854_);
  nor (_21577_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21578_, _10084_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21579_, _21578_, _21577_);
  and (_21580_, _21579_, _20682_);
  not (_21581_, _21580_);
  nor (_21582_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21583_, _09819_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21584_, _21583_, _21582_);
  and (_21585_, _21584_, _20681_);
  nor (_21586_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21587_, _10388_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21588_, _21587_, _21586_);
  and (_21589_, _21588_, _20656_);
  nor (_21590_, _21589_, _21585_);
  and (_21591_, _21590_, _21581_);
  and (_21592_, _21591_, _21576_);
  nor (_21593_, _21592_, _21571_);
  and (_21594_, _21593_, _21543_);
  nor (_21595_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21596_, _09333_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21597_, _21596_, _21595_);
  and (_21598_, _21597_, _20656_);
  nor (_21599_, _21598_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21600_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21601_, _08809_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21602_, _21601_, _21600_);
  and (_21603_, _21602_, _20681_);
  not (_21604_, _21603_);
  nor (_21605_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21606_, _09080_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21607_, _21606_, _21605_);
  and (_21608_, _21607_, _20682_);
  nor (_21609_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21610_, _08556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21611_, _21610_, _21609_);
  and (_21612_, _21611_, _21527_);
  nor (_21613_, _21612_, _21608_);
  and (_21614_, _21613_, _21604_);
  and (_21615_, _21614_, _21599_);
  nor (_21616_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21617_, _10369_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21618_, _21617_, _21616_);
  and (_21619_, _21618_, _20656_);
  nor (_21620_, _21619_, _22854_);
  nor (_21621_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21622_, _09802_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21623_, _21622_, _21621_);
  and (_21624_, _21623_, _20681_);
  not (_21625_, _21624_);
  nor (_21626_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21627_, _10069_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21628_, _21627_, _21626_);
  and (_21629_, _21628_, _20682_);
  nor (_21630_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21631_, _09570_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21632_, _21631_, _21630_);
  and (_21633_, _21632_, _21527_);
  nor (_21634_, _21633_, _21629_);
  and (_21635_, _21634_, _21625_);
  and (_21636_, _21635_, _21620_);
  nor (_21637_, _21636_, _21615_);
  and (_21638_, _21637_, _21543_);
  nor (_21639_, _21638_, _21594_);
  nor (_21640_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21641_, _08857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21642_, _21641_, _21640_);
  and (_21643_, _21642_, _20681_);
  nor (_21644_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21645_, _09128_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21646_, _21645_, _21644_);
  and (_21647_, _21646_, _20682_);
  nor (_21648_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21649_, _08602_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21650_, _21649_, _21648_);
  and (_21651_, _21650_, _21527_);
  nor (_21652_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21653_, _09389_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21654_, _21653_, _21652_);
  and (_21655_, _21654_, _20656_);
  or (_21656_, _21655_, _21651_);
  or (_21657_, _21656_, _21647_);
  or (_21658_, _21657_, _21643_);
  and (_21659_, _21658_, _22854_);
  nor (_21660_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21661_, _09849_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21662_, _21661_, _21660_);
  and (_21663_, _21662_, _20681_);
  nor (_21664_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21665_, _10118_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21666_, _21665_, _21664_);
  and (_21667_, _21666_, _20682_);
  nor (_21668_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21669_, _09613_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21670_, _21669_, _21668_);
  and (_21671_, _21670_, _21527_);
  nor (_21672_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21673_, _10426_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21674_, _21673_, _21672_);
  and (_21675_, _21674_, _20656_);
  or (_21676_, _21675_, _21671_);
  or (_21677_, _21676_, _21667_);
  or (_21678_, _21677_, _21663_);
  and (_21679_, _21678_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21680_, _21679_, _21659_);
  and (_21681_, _21680_, _21543_);
  nor (_21682_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21683_, _08844_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21684_, _21683_, _21682_);
  and (_21685_, _21684_, _20681_);
  nor (_21686_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21687_, _09113_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21688_, _21687_, _21686_);
  and (_21689_, _21688_, _20682_);
  nor (_21690_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21691_, _08589_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21692_, _21691_, _21690_);
  and (_21693_, _21692_, _21527_);
  nor (_21694_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21695_, _09371_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21696_, _21695_, _21694_);
  and (_21697_, _21696_, _20656_);
  or (_21698_, _21697_, _21693_);
  or (_21699_, _21698_, _21689_);
  or (_21700_, _21699_, _21685_);
  and (_21701_, _21700_, _22854_);
  nor (_21702_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21703_, _09834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21704_, _21703_, _21702_);
  and (_21705_, _21704_, _20681_);
  nor (_21706_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21707_, _10102_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21708_, _21707_, _21706_);
  and (_21709_, _21708_, _20682_);
  nor (_21710_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21711_, _09598_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21712_, _21711_, _21710_);
  and (_21713_, _21712_, _21527_);
  nor (_21714_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21715_, _10410_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21716_, _21715_, _21714_);
  and (_21717_, _21716_, _20656_);
  or (_21718_, _21717_, _21713_);
  or (_21719_, _21718_, _21709_);
  or (_21720_, _21719_, _21705_);
  and (_21721_, _21720_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21722_, _21721_, _21701_);
  and (_21723_, _21722_, _21543_);
  nor (_21724_, _21723_, _21681_);
  and (_21725_, _21724_, _21639_);
  nor (_21726_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21727_, _08883_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21728_, _21727_, _21726_);
  and (_21729_, _21728_, _20681_);
  nor (_21730_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21731_, _09153_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21732_, _21731_, _21730_);
  and (_21733_, _21732_, _20682_);
  nor (_21734_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21735_, _08630_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21736_, _21735_, _21734_);
  and (_21737_, _21736_, _21527_);
  nor (_21738_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21739_, _09415_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21740_, _21739_, _21738_);
  and (_21741_, _21740_, _20656_);
  or (_21742_, _21741_, _21737_);
  or (_21743_, _21742_, _21733_);
  or (_21744_, _21743_, _21729_);
  and (_21745_, _21744_, _22854_);
  nor (_21746_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21747_, _09875_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21748_, _21747_, _21746_);
  and (_21749_, _21748_, _20681_);
  nor (_21750_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21751_, _10150_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21752_, _21751_, _21750_);
  and (_21753_, _21752_, _20682_);
  nor (_21754_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21755_, _09641_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21756_, _21755_, _21754_);
  and (_21757_, _21756_, _21527_);
  nor (_21758_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21759_, _10453_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21760_, _21759_, _21758_);
  and (_21761_, _21760_, _20656_);
  or (_21762_, _21761_, _21757_);
  or (_21763_, _21762_, _21753_);
  or (_21764_, _21763_, _21749_);
  and (_21765_, _21764_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21766_, _21765_, _21745_);
  and (_21767_, _21766_, _21543_);
  nor (_21768_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21769_, _08617_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21770_, _21769_, _21768_);
  and (_21771_, _21770_, _21527_);
  nor (_21772_, _21771_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21773_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21774_, _09141_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21775_, _21774_, _21773_);
  and (_21776_, _21775_, _20682_);
  not (_21777_, _21776_);
  nor (_21778_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21779_, _08870_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21780_, _21779_, _21778_);
  and (_21781_, _21780_, _20681_);
  nor (_21782_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21783_, _09402_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21784_, _21783_, _21782_);
  and (_21785_, _21784_, _20656_);
  nor (_21786_, _21785_, _21781_);
  and (_21787_, _21786_, _21777_);
  and (_21788_, _21787_, _21772_);
  nor (_21789_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21790_, _09627_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21791_, _21790_, _21789_);
  and (_21792_, _21791_, _21527_);
  nor (_21793_, _21792_, _22854_);
  nor (_21794_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21795_, _10135_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21796_, _21795_, _21794_);
  and (_21797_, _21796_, _20682_);
  not (_21798_, _21797_);
  nor (_21799_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21800_, _09863_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21801_, _21800_, _21799_);
  and (_21802_, _21801_, _20681_);
  nor (_21803_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21804_, _10441_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21805_, _21804_, _21803_);
  and (_21806_, _21805_, _20656_);
  nor (_21807_, _21806_, _21802_);
  and (_21808_, _21807_, _21798_);
  and (_21809_, _21808_, _21793_);
  nor (_21810_, _21809_, _21788_);
  and (_21811_, _21810_, _21543_);
  nor (_21812_, _21811_, _21767_);
  nor (_21813_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21814_, _07675_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21815_, _21814_, _21813_);
  and (_21816_, _21815_, _21527_);
  nor (_21817_, _21816_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21818_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21819_, _07689_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21821_, _21819_, _21818_);
  and (_21822_, _21821_, _20682_);
  not (_21823_, _21822_);
  nor (_21824_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21825_, _07696_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21826_, _21825_, _21824_);
  and (_21827_, _21826_, _20681_);
  nor (_21828_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21829_, _07682_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21830_, _21829_, _21828_);
  and (_21831_, _21830_, _20656_);
  nor (_21832_, _21831_, _21827_);
  and (_21833_, _21832_, _21823_);
  and (_21834_, _21833_, _21817_);
  nor (_21835_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21836_, _07709_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21837_, _21836_, _21835_);
  and (_21838_, _21837_, _21527_);
  nor (_21839_, _21838_, _22854_);
  nor (_21840_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21841_, _07717_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21842_, _21841_, _21840_);
  and (_21843_, _21842_, _20682_);
  not (_21844_, _21843_);
  nor (_21845_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21846_, _07731_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21847_, _21846_, _21845_);
  and (_21848_, _21847_, _20681_);
  nor (_21849_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21850_, _07723_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21851_, _21850_, _21849_);
  and (_21852_, _21851_, _20656_);
  nor (_21853_, _21852_, _21848_);
  and (_21854_, _21853_, _21844_);
  and (_21855_, _21854_, _21839_);
  nor (_21856_, _21855_, _21834_);
  and (_21857_, _21856_, _21543_);
  nor (_21858_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21859_, _08646_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21860_, _21859_, _21858_);
  and (_21861_, _21860_, _21527_);
  nor (_21862_, _21861_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21863_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21864_, _09166_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21865_, _21864_, _21863_);
  and (_21866_, _21865_, _20682_);
  not (_21867_, _21866_);
  nor (_21868_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21869_, _08898_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21870_, _21869_, _21868_);
  and (_21871_, _21870_, _20681_);
  nor (_21872_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21873_, _09428_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21874_, _21873_, _21872_);
  and (_21875_, _21874_, _20656_);
  nor (_21876_, _21875_, _21871_);
  and (_21877_, _21876_, _21867_);
  and (_21878_, _21877_, _21862_);
  nor (_21879_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21880_, _09654_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21881_, _21880_, _21879_);
  and (_21882_, _21881_, _21527_);
  nor (_21883_, _21882_, _22854_);
  nor (_21884_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21885_, _10166_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21886_, _21885_, _21884_);
  and (_21887_, _21886_, _20682_);
  not (_21888_, _21887_);
  nor (_21889_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21890_, _09888_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21891_, _21890_, _21889_);
  and (_21892_, _21891_, _20681_);
  nor (_21893_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21894_, _10467_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21895_, _21894_, _21893_);
  and (_21896_, _21895_, _20656_);
  nor (_21897_, _21896_, _21892_);
  and (_21898_, _21897_, _21888_);
  and (_21899_, _21898_, _21883_);
  nor (_21900_, _21899_, _21878_);
  not (_21901_, _21900_);
  and (_21902_, _21901_, _21857_);
  and (_21903_, _21902_, _21812_);
  and (_21904_, _21903_, _21725_);
  and (_21905_, _21904_, _21550_);
  and (_21906_, _21905_, _21270_);
  not (_21907_, _21857_);
  and (_21908_, _21900_, _21543_);
  nand (_21909_, _21811_, _21766_);
  and (_21910_, _21723_, _21594_);
  nor (_21911_, _21910_, _21680_);
  nor (_21912_, _21911_, _21909_);
  not (_21913_, _21638_);
  and (_21914_, _21724_, _21913_);
  and (_21915_, _21914_, _21594_);
  not (_21916_, _21637_);
  not (_21917_, _21593_);
  not (_21918_, _21680_);
  and (_21919_, _21723_, _21918_);
  and (_21920_, _21919_, _21917_);
  and (_21921_, _21920_, _21916_);
  or (_21922_, _21921_, _21915_);
  or (_21923_, _21922_, _21912_);
  and (_21924_, _21923_, _21908_);
  and (_21925_, _21901_, _21767_);
  and (_21926_, _21925_, _21920_);
  not (_21927_, _21767_);
  and (_21928_, _21920_, _21638_);
  and (_21929_, _21928_, _21927_);
  or (_21930_, _21929_, _21926_);
  or (_21931_, _21930_, _21924_);
  and (_21932_, _21931_, _21907_);
  and (_21933_, _21915_, _21927_);
  not (_21934_, _21908_);
  nor (_21935_, _21934_, _21766_);
  and (_21936_, _21935_, _21914_);
  and (_21937_, _21908_, _21766_);
  and (_21938_, _21937_, _21928_);
  or (_21939_, _21938_, _21936_);
  or (_21940_, _21939_, _21933_);
  and (_21941_, _21940_, _21857_);
  not (_21942_, _21810_);
  and (_21943_, _21908_, _21942_);
  and (_21944_, _21943_, _21928_);
  and (_21945_, _21811_, _21927_);
  and (_21946_, _21945_, _21920_);
  and (_21947_, _21767_, _21914_);
  and (_21948_, _21942_, _21681_);
  not (_21949_, _21811_);
  and (_21950_, _21910_, _21949_);
  or (_21951_, _21950_, _21948_);
  or (_21952_, _21951_, _21947_);
  or (_21953_, _21952_, _21946_);
  and (_21954_, _21953_, _21902_);
  or (_21955_, _21954_, _21944_);
  or (_21956_, _21955_, _21941_);
  or (_21957_, _21956_, _21932_);
  nor (_21958_, _20782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_21959_, _20782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_21960_, _21959_, _21958_);
  nor (_21961_, _20786_, _22827_);
  and (_21962_, _20786_, _22827_);
  or (_21963_, _21962_, _21961_);
  or (_21964_, _21963_, _21960_);
  and (_21965_, _20670_, _22837_);
  nor (_21966_, _20670_, _22837_);
  or (_21967_, _21966_, _21965_);
  or (_21968_, _21967_, _21157_);
  or (_21969_, _21968_, _21964_);
  or (_21970_, _20796_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_21971_, _20796_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_21972_, _21971_, _21970_);
  or (_21973_, _21197_, _21182_);
  and (_21974_, _20817_, _22802_);
  nor (_21975_, _20683_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21976_, _20683_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_21977_, _21976_, _21975_);
  nor (_21978_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_21979_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_21980_, _21979_, _21978_);
  not (_21981_, _21980_);
  and (_21982_, _21981_, _20657_);
  or (_21983_, _21982_, _21977_);
  and (_21984_, _20676_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21985_, _20676_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21986_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_21987_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_21988_, _21987_, _21986_);
  nand (_21989_, _21988_, _21233_);
  nor (_21990_, _21981_, _20657_);
  or (_21991_, _21990_, _21989_);
  or (_21992_, _21991_, _21985_);
  or (_21993_, _21992_, _21984_);
  or (_21994_, _21993_, _21983_);
  nor (_21995_, _20817_, _22802_);
  or (_21996_, _21995_, _21994_);
  or (_21997_, _21996_, _21974_);
  or (_21998_, _20806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_21999_, _20806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_22000_, _21999_, _21998_);
  nor (_22001_, _20862_, _22798_);
  and (_22002_, _20862_, _22798_);
  or (_22003_, _22002_, _22001_);
  nor (_22004_, _20811_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_22005_, _20811_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_22006_, _22005_, _22004_);
  or (_22007_, _22006_, _22003_);
  or (_22008_, _22007_, _22000_);
  or (_22009_, _22008_, _21997_);
  or (_22010_, _22009_, _21973_);
  or (_22011_, _22010_, _21972_);
  or (_22012_, _22011_, _21969_);
  and (_22013_, _22012_, _21957_);
  and (_22014_, _21638_, _21594_);
  and (_22015_, _22014_, _21724_);
  and (_22016_, _21921_, _21812_);
  or (_22017_, _22016_, _22015_);
  nor (_22018_, _21766_, _21637_);
  nand (_22019_, _22018_, _21723_);
  nand (_22020_, _21812_, _21639_);
  and (_22021_, _22020_, _22019_);
  nor (_22022_, _22021_, _21857_);
  or (_22023_, _22022_, _22017_);
  and (_22024_, _22023_, _21934_);
  and (_22025_, _21926_, _21949_);
  or (_22026_, _21919_, _21767_);
  or (_22027_, _21680_, _21916_);
  and (_22028_, _22027_, _21908_);
  and (_22029_, _22028_, _22026_);
  or (_22030_, _22029_, _22025_);
  and (_22031_, _22030_, _21857_);
  nor (_22032_, _21856_, _21766_);
  not (_22033_, _21856_);
  or (_22034_, _21945_, _22033_);
  and (_22035_, _22034_, _21901_);
  or (_22036_, _22035_, _22032_);
  and (_22037_, _22036_, _21681_);
  nor (_22038_, _21908_, _21857_);
  or (_22039_, _21942_, _21767_);
  nor (_22040_, _22039_, _21681_);
  or (_22041_, _22040_, _22038_);
  and (_22042_, _22041_, _21910_);
  and (_22043_, _21948_, _21908_);
  nor (_22044_, _22027_, _22033_);
  and (_22045_, _22044_, _21594_);
  or (_22046_, _22045_, _21950_);
  and (_22047_, _22046_, _21908_);
  or (_22048_, _22047_, _22043_);
  or (_22049_, _22048_, _22042_);
  or (_22050_, _22049_, _22037_);
  or (_22051_, _22050_, _22031_);
  or (_22052_, _22051_, _22024_);
  and (_22053_, _20780_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_22054_, _22053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_22055_, _22054_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22056_, _22053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22057_, _22056_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or (_22058_, _22057_, _22055_);
  and (_22059_, _22058_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_22060_, _20791_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_22061_, _22890_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22062_, _22061_, _22060_);
  nor (_22063_, _22062_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_22064_, _22062_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not (_22065_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_22066_, _20657_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22067_, _22066_, _20660_);
  and (_22068_, _22067_, _20664_);
  and (_22069_, _22068_, _22065_);
  nor (_22070_, _22068_, _22065_);
  or (_22071_, _22070_, _22069_);
  and (_22072_, _22071_, _22827_);
  or (_22073_, _22072_, _22064_);
  or (_22074_, _22073_, _22063_);
  and (_22075_, _22067_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_22076_, _22075_, _22882_);
  nor (_22077_, _22075_, _22882_);
  nor (_22078_, _22077_, _22076_);
  and (_22079_, _22078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_22080_, _20678_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22081_, _20678_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22082_, _22081_, _22080_);
  and (_22083_, _20808_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22084_, _22083_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_22085_, _22084_, _22067_);
  nor (_22086_, _22085_, _22806_);
  and (_22087_, _22085_, _22806_);
  or (_22088_, _22087_, _22086_);
  or (_22089_, _22088_, _22082_);
  nor (_22090_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_22091_, _22090_, _22083_);
  nor (_22092_, _22091_, _20816_);
  and (_22093_, _22092_, _22802_);
  nor (_22094_, _20685_, _22783_);
  and (_22095_, _20685_, _22783_);
  or (_22096_, _22095_, _22094_);
  nand (_22097_, _21988_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_22098_, _21988_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22099_, _22098_, _22097_);
  nor (_22100_, _22066_, _21981_);
  and (_22101_, _22066_, _21981_);
  or (_22102_, _22101_, _21233_);
  or (_22103_, _22102_, _22100_);
  or (_22104_, _22103_, _22099_);
  or (_22105_, _22104_, _22096_);
  or (_22106_, _22105_, _22093_);
  or (_22107_, _22106_, _22089_);
  or (_22108_, _22864_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_22109_, _20862_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22110_, _22109_, _22108_);
  and (_22111_, _22110_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_22112_, _22110_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_22113_, _22112_, _22111_);
  or (_22114_, _22113_, _22107_);
  or (_22115_, _22114_, _22079_);
  nor (_22116_, _22071_, _22827_);
  nor (_22117_, _22078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or (_22118_, _22117_, _22116_);
  or (_22119_, _22118_, _22115_);
  or (_22120_, _22119_, _22074_);
  or (_22121_, _22120_, _22059_);
  nor (_22122_, _22057_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_22123_, _22122_, _21152_);
  nor (_22124_, _22123_, _22055_);
  or (_22125_, _20782_, _22841_);
  or (_22126_, _22897_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22127_, _22126_, _22125_);
  and (_22128_, _22127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22129_, _22067_, _20662_);
  and (_22130_, _22129_, _22886_);
  nor (_22131_, _22129_, _22886_);
  or (_22132_, _22131_, _22130_);
  nor (_22133_, _22132_, _22819_);
  and (_22134_, _22132_, _22819_);
  nor (_22135_, _22067_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_22136_, _22135_, _22075_);
  and (_22137_, _22136_, _22810_);
  nor (_22138_, _22136_, _22810_);
  nor (_22139_, _22092_, _22802_);
  or (_22140_, _22139_, _22138_);
  or (_22141_, _22140_, _22137_);
  or (_22142_, _22141_, _22134_);
  or (_22143_, _22142_, _22133_);
  or (_22144_, _22143_, _22128_);
  nor (_22145_, _22127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22146_, _22055_, _21153_);
  or (_22147_, _22146_, _22145_);
  or (_22148_, _22147_, _22144_);
  or (_22149_, _22148_, _22124_);
  or (_22150_, _22149_, _22121_);
  and (_22151_, _22150_, _22052_);
  and (_22152_, _21945_, _21725_);
  and (_22153_, _21929_, _21942_);
  or (_22154_, _22153_, _22152_);
  and (_22155_, _22154_, _21902_);
  and (_22156_, _21938_, _21811_);
  and (_22157_, _21909_, _21908_);
  and (_22158_, _22157_, _22015_);
  or (_22159_, _22158_, _22156_);
  and (_22160_, _22159_, _21907_);
  or (_22161_, _22160_, _22155_);
  and (_22162_, _21432_, _20660_);
  and (_22163_, _22162_, _20663_);
  and (_22164_, _22163_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_22165_, _22164_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_22166_, _22165_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_22167_, _22166_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_22168_, _22166_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_22169_, _22168_, _22167_);
  nor (_22170_, _22169_, _22837_);
  nor (_22171_, _22165_, _22897_);
  and (_22172_, _22165_, _22897_);
  nor (_22173_, _22172_, _22171_);
  nor (_22174_, _22173_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22175_, _22169_, _22837_);
  or (_22176_, _22175_, _22174_);
  or (_22177_, _22176_, _22170_);
  nor (_22178_, _22164_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_22179_, _22178_, _22165_);
  and (_22180_, _22179_, _22827_);
  nor (_22181_, _22179_, _22827_);
  or (_22182_, _22181_, _22180_);
  nor (_22183_, _22167_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_22184_, _22167_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_22185_, _22184_, _22183_);
  nor (_22186_, _22185_, _14710_);
  or (_22187_, _22186_, _22182_);
  and (_22188_, _22162_, _20662_);
  nor (_22189_, _22188_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_22190_, _22189_, _22163_);
  and (_22191_, _22190_, _22819_);
  and (_22192_, _22185_, _14710_);
  or (_22193_, _22192_, _22191_);
  and (_22194_, _22173_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22195_, _21432_, _20659_);
  and (_22196_, _21432_, _20658_);
  nor (_22197_, _22196_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_22198_, _22197_, _22195_);
  and (_22199_, _22198_, _22802_);
  nor (_22200_, _22163_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_22201_, _22200_, _22164_);
  nor (_22202_, _22201_, _22823_);
  and (_22203_, _22162_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_22204_, _22162_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_22205_, _22204_, _22203_);
  nor (_22206_, _22205_, _22810_);
  and (_22207_, _22205_, _22810_);
  or (_22208_, _22207_, _22206_);
  or (_22209_, _22208_, _22202_);
  or (_22210_, _22209_, _22199_);
  or (_22211_, _22210_, _22194_);
  and (_22212_, _22201_, _22823_);
  nor (_22213_, _22203_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_22214_, _22213_, _22188_);
  nor (_22215_, _22214_, _22814_);
  and (_22216_, _22214_, _22814_);
  or (_22217_, _22216_, _22215_);
  nor (_22218_, _22195_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_22219_, _22218_, _22162_);
  and (_22220_, _22219_, _22806_);
  nor (_22221_, _22190_, _22819_);
  or (_22222_, _22221_, _22220_);
  or (_22223_, _22222_, _22217_);
  or (_22224_, _21980_, _21432_);
  nand (_22225_, _21980_, _21432_);
  and (_22226_, _22225_, _22224_);
  nand (_22227_, _21430_, _22783_);
  nand (_22228_, _22227_, _22099_);
  or (_22229_, _22228_, _22226_);
  and (_22230_, _21432_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_22231_, _22230_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_22232_, _22231_, _22196_);
  and (_22233_, _22232_, _22798_);
  nor (_22234_, _22198_, _22802_);
  or (_22235_, _22234_, _22233_);
  nor (_22236_, _22232_, _22798_);
  nor (_22237_, _21430_, _22783_);
  or (_22238_, _22237_, _21233_);
  or (_22239_, _22238_, _22236_);
  or (_22240_, _22239_, _22235_);
  nor (_22241_, _22219_, _22806_);
  or (_22242_, _21434_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_22243_, _21434_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22244_, _22243_, _22242_);
  or (_22245_, _22244_, _22241_);
  or (_22246_, _22245_, _22240_);
  or (_22247_, _22246_, _22229_);
  or (_22248_, _22247_, _22223_);
  or (_22249_, _22248_, _22212_);
  or (_22250_, _22249_, _22211_);
  or (_22251_, _22250_, _22193_);
  or (_22252_, _22251_, _22187_);
  or (_22253_, _22252_, _22177_);
  and (_22254_, _22253_, _22161_);
  or (_22255_, _22254_, _22151_);
  or (_22256_, _22255_, _22013_);
  and (_22257_, _22256_, _21550_);
  or (_22258_, _20984_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_22259_, _20984_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22260_, _22259_, _22258_);
  or (_22261_, _20900_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_22262_, _20900_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_22263_, _22262_, _22261_);
  or (_22264_, _22263_, _22260_);
  or (_22265_, _21066_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_22266_, _21066_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_22267_, _22266_, _22265_);
  and (_22268_, _21105_, _22772_);
  nor (_22269_, _21027_, _22783_);
  or (_22270_, _22269_, _22268_);
  or (_22271_, _22270_, _22267_);
  and (_22272_, _21767_, _22810_);
  nor (_22273_, _21767_, _22810_);
  or (_22274_, _22273_, _22272_);
  nor (_22275_, _21908_, _22814_);
  and (_22276_, _21908_, _22814_);
  or (_22277_, _22276_, _22275_);
  or (_22278_, _22277_, _22274_);
  nor (_22279_, _21857_, _22819_);
  and (_22280_, _21857_, _22819_);
  or (_22281_, _22280_, _22279_);
  or (_22282_, _22281_, _21182_);
  or (_22283_, _22282_, _22278_);
  nor (_22284_, _21105_, _22772_);
  or (_22285_, _22284_, _21969_);
  or (_22286_, _22285_, _22283_);
  or (_22287_, _22286_, _22271_);
  or (_22288_, _20775_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_22289_, _20775_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_22290_, _22289_, _22288_);
  and (_22291_, _20855_, _22802_);
  or (_22292_, _22291_, _22290_);
  nor (_22293_, _20855_, _22802_);
  and (_22294_, _20942_, _22794_);
  or (_22295_, _22294_, _22293_);
  nor (_22296_, _20942_, _22794_);
  and (_22297_, _21027_, _22783_);
  or (_22298_, _22297_, _22296_);
  or (_22299_, _22298_, _22295_);
  or (_22300_, _22299_, _22292_);
  or (_22301_, _22300_, _22287_);
  or (_22302_, _22301_, _22264_);
  and (_22303_, _21638_, _21917_);
  and (_22304_, _22303_, _21724_);
  and (_22305_, _22304_, _22302_);
  and (_22306_, _21886_, _20681_);
  or (_22307_, _22306_, _20676_);
  and (_22308_, _21881_, _20656_);
  and (_22309_, _21891_, _21527_);
  and (_22310_, _21895_, _20682_);
  or (_22311_, _22310_, _22309_);
  or (_22312_, _22311_, _22308_);
  or (_22313_, _22312_, _22307_);
  and (_22314_, _21865_, _20681_);
  or (_22315_, _22314_, _20946_);
  and (_22316_, _21860_, _20656_);
  and (_22317_, _21870_, _21527_);
  and (_22318_, _21874_, _20682_);
  or (_22319_, _22318_, _22317_);
  or (_22320_, _22319_, _22316_);
  or (_22321_, _22320_, _22315_);
  nand (_22322_, _22321_, _22313_);
  nor (_22323_, _22322_, _21523_);
  nand (_22324_, _22323_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_22325_, _22323_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_22326_, _22325_, _22324_);
  not (_22327_, _21523_);
  and (_22328_, _21842_, _20681_);
  and (_22329_, _21851_, _20682_);
  nor (_22330_, _22329_, _22328_);
  and (_22331_, _21837_, _20656_);
  and (_22332_, _21847_, _21527_);
  nor (_22333_, _22332_, _22331_);
  and (_22334_, _22333_, _22330_);
  and (_22335_, _22334_, _20946_);
  and (_22336_, _21830_, _20682_);
  and (_22337_, _21815_, _20656_);
  and (_22338_, _21821_, _20681_);
  or (_22339_, _22338_, _22337_);
  nor (_22340_, _22339_, _22336_);
  and (_22341_, _21826_, _21527_);
  nor (_22342_, _22341_, _20946_);
  and (_22343_, _22342_, _22340_);
  nor (_22344_, _22343_, _22335_);
  and (_22345_, _22344_, _22327_);
  nor (_22346_, _22345_, _22806_);
  and (_22347_, _22345_, _22806_);
  or (_22348_, _22347_, _22346_);
  or (_22349_, _22348_, _22326_);
  and (_22350_, _21732_, _20681_);
  or (_22351_, _22350_, _20946_);
  and (_22352_, _21736_, _20656_);
  and (_22353_, _21728_, _21527_);
  and (_22354_, _21740_, _20682_);
  or (_22355_, _22354_, _22353_);
  or (_22356_, _22355_, _22352_);
  or (_22357_, _22356_, _22351_);
  and (_22358_, _21752_, _20681_);
  or (_22359_, _22358_, _20676_);
  and (_22360_, _21756_, _20656_);
  and (_22361_, _21748_, _21527_);
  and (_22362_, _21760_, _20682_);
  or (_22363_, _22362_, _22361_);
  or (_22364_, _22363_, _22360_);
  or (_22365_, _22364_, _22359_);
  nand (_22366_, _22365_, _22357_);
  nor (_22367_, _22366_, _21523_);
  nand (_22368_, _22367_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_22369_, _22367_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_22370_, _22369_, _22368_);
  and (_22371_, _21775_, _20681_);
  and (_22372_, _21784_, _20682_);
  and (_22373_, _21770_, _20656_);
  or (_22374_, _22373_, _22372_);
  or (_22375_, _22374_, _22371_);
  and (_22376_, _21780_, _21527_);
  or (_22377_, _22376_, _20946_);
  or (_22378_, _22377_, _22375_);
  and (_22379_, _21796_, _20681_);
  or (_22380_, _22379_, _20676_);
  and (_22381_, _21791_, _20656_);
  and (_22382_, _21801_, _21527_);
  and (_22383_, _21805_, _20682_);
  or (_22384_, _22383_, _22382_);
  or (_22385_, _22384_, _22381_);
  or (_22386_, _22385_, _22380_);
  nand (_22387_, _22386_, _22378_);
  nor (_22388_, _22387_, _21523_);
  nand (_22389_, _22388_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_22390_, _22388_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_22391_, _22390_, _22389_);
  or (_22392_, _22391_, _22370_);
  or (_22393_, _22392_, _22349_);
  and (_22394_, _21646_, _20681_);
  or (_22395_, _22394_, _20946_);
  and (_22396_, _21650_, _20656_);
  and (_22397_, _21642_, _21527_);
  and (_22398_, _21654_, _20682_);
  or (_22399_, _22398_, _22397_);
  or (_22400_, _22399_, _22396_);
  or (_22401_, _22400_, _22395_);
  and (_22402_, _21666_, _20681_);
  or (_22403_, _22402_, _20676_);
  and (_22404_, _21670_, _20656_);
  and (_22405_, _21662_, _21527_);
  and (_22406_, _21674_, _20682_);
  or (_22407_, _22406_, _22405_);
  or (_22408_, _22407_, _22404_);
  or (_22409_, _22408_, _22403_);
  nand (_22410_, _22409_, _22401_);
  nor (_22411_, _22410_, _21523_);
  nand (_22412_, _22411_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22413_, _22411_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22414_, _22413_, _22412_);
  and (_22415_, _21704_, _21527_);
  and (_22416_, _21716_, _20682_);
  and (_22417_, _21712_, _20656_);
  and (_22418_, _21708_, _20681_);
  or (_22419_, _22418_, _22417_);
  or (_22420_, _22419_, _22416_);
  or (_22421_, _22420_, _22415_);
  and (_22422_, _22421_, _20946_);
  and (_22423_, _21684_, _21527_);
  and (_22424_, _21696_, _20682_);
  and (_22425_, _21692_, _20656_);
  and (_22426_, _21688_, _20681_);
  or (_22427_, _22426_, _22425_);
  or (_22428_, _22427_, _22424_);
  or (_22429_, _22428_, _22423_);
  and (_22430_, _22429_, _20676_);
  or (_22431_, _22430_, _22422_);
  and (_22432_, _22431_, _22327_);
  and (_22433_, _22432_, _22783_);
  nor (_22434_, _22432_, _22783_);
  or (_22435_, _22434_, _22433_);
  or (_22436_, _22435_, _22414_);
  and (_22437_, _21588_, _20682_);
  and (_22438_, _21579_, _20681_);
  nor (_22439_, _22438_, _22437_);
  and (_22440_, _21584_, _21527_);
  and (_22441_, _21574_, _20656_);
  nor (_22442_, _22441_, _22440_);
  and (_22443_, _22442_, _22439_);
  nor (_22444_, _22443_, _20676_);
  and (_22445_, _21567_, _20682_);
  and (_22446_, _21558_, _20681_);
  nor (_22447_, _22446_, _22445_);
  and (_22448_, _21563_, _21527_);
  and (_22449_, _21553_, _20656_);
  nor (_22450_, _22449_, _22448_);
  and (_22451_, _22450_, _22447_);
  nor (_22452_, _22451_, _20946_);
  nor (_22453_, _22452_, _22444_);
  nor (_22454_, _22453_, _21523_);
  and (_22455_, _22454_, _22778_);
  nor (_22456_, _22454_, _22778_);
  or (_22457_, _22456_, _22455_);
  and (_22458_, _21607_, _20681_);
  or (_22459_, _22458_, _20946_);
  and (_22460_, _21611_, _20656_);
  and (_22461_, _21602_, _21527_);
  and (_22462_, _21597_, _20682_);
  or (_22463_, _22462_, _22461_);
  or (_22464_, _22463_, _22460_);
  or (_22465_, _22464_, _22459_);
  and (_22466_, _21628_, _20681_);
  or (_22467_, _22466_, _20676_);
  and (_22468_, _21632_, _20656_);
  and (_22469_, _21623_, _21527_);
  and (_22470_, _21618_, _20682_);
  or (_22471_, _22470_, _22469_);
  or (_22472_, _22471_, _22468_);
  or (_22473_, _22472_, _22467_);
  nand (_22474_, _22473_, _22465_);
  nor (_22475_, _22474_, _21523_);
  and (_22476_, _22475_, _22772_);
  nor (_22477_, _22475_, _22772_);
  or (_22478_, _22477_, _22476_);
  or (_22479_, _22478_, _22457_);
  or (_22480_, _22479_, _22436_);
  or (_22481_, _22480_, _22393_);
  or (_22482_, _21066_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_22483_, _21066_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_22484_, _22483_, _22482_);
  and (_22485_, _21105_, _22810_);
  nor (_22486_, _21105_, _22810_);
  or (_22487_, _22486_, _22485_);
  or (_22488_, _22487_, _22484_);
  or (_22489_, _20984_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_22490_, _20984_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_22491_, _22490_, _22489_);
  nor (_22492_, _21027_, _22819_);
  and (_22493_, _21027_, _22819_);
  or (_22494_, _22493_, _22492_);
  or (_22495_, _22494_, _22491_);
  or (_22496_, _22495_, _22488_);
  and (_22497_, _20942_, _22827_);
  nor (_22498_, _20942_, _22827_);
  or (_22499_, _22498_, _22497_);
  or (_22500_, _20900_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_22501_, _20900_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22502_, _22501_, _22500_);
  or (_22503_, _22502_, _22499_);
  and (_22504_, _20775_, _14710_);
  nor (_22505_, _20775_, _14710_);
  or (_22506_, _22505_, _22504_);
  and (_22507_, _20855_, _22837_);
  nor (_22508_, _20855_, _22837_);
  or (_22509_, _22508_, _22507_);
  or (_22510_, _22509_, _22506_);
  or (_22511_, _22510_, _22503_);
  or (_22512_, _22511_, _22496_);
  or (_22513_, _22512_, _22481_);
  and (_22514_, _22038_, _21933_);
  and (_22515_, _22514_, _22513_);
  or (_22516_, _22515_, _22305_);
  and (_22517_, _22516_, _21550_);
  or (_22518_, _22517_, _22257_);
  or (property_invalid, _22518_, _21906_);
  and (_22519_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not (_22520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_22521_, _25687_, _25024_);
  nor (_22522_, _22521_, _22520_);
  and (_22523_, _22521_, _22520_);
  nor (_22524_, _22523_, _22522_);
  nor (_22525_, _22524_, _24127_);
  and (_22526_, _24127_, _23642_);
  or (_22527_, _22526_, _22525_);
  and (_22528_, _22527_, _24166_);
  or (_12540_, _22528_, _22519_);
  and (_22529_, _03300_, _23707_);
  and (_22530_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_12543_, _22530_, _22529_);
  and (_22531_, _18217_, _23946_);
  and (_22532_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_12545_, _22532_, _22531_);
  and (_22533_, _21544_, first_instr);
  or (_00000_, _22533_, rst);
  and (_22534_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  and (_22535_, _16331_, _23707_);
  or (_12565_, _22535_, _22534_);
  and (_22536_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  and (_22537_, _16331_, _24050_);
  or (_12569_, _22537_, _22536_);
  and (_22538_, _18217_, _23649_);
  and (_22539_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_12586_, _22539_, _22538_);
  and (_22540_, _25739_, _24050_);
  and (_22541_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or (_12613_, _22541_, _22540_);
  and (_22543_, _03300_, _24050_);
  and (_22544_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_12615_, _22544_, _22543_);
  and (_22545_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and (_22546_, _16325_, _23778_);
  or (_12617_, _22546_, _22545_);
  and (_22547_, _18217_, _23747_);
  and (_22548_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_27215_, _22548_, _22547_);
  and (_22549_, _10347_, _23824_);
  and (_22550_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or (_12632_, _22550_, _22549_);
  and (_22551_, _08548_, _23778_);
  and (_22552_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or (_27136_, _22552_, _22551_);
  and (_22553_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and (_22554_, _06507_, _23649_);
  or (_12672_, _22554_, _22553_);
  and (_22555_, _03300_, _23946_);
  and (_22556_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_12674_, _22556_, _22555_);
  and (_22557_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  and (_22558_, _16331_, _23898_);
  or (_12679_, _22558_, _22557_);
  and (_22559_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  and (_22560_, _16331_, _23778_);
  or (_12681_, _22560_, _22559_);
  and (_22561_, _08548_, _23824_);
  and (_22562_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  or (_12704_, _22562_, _22561_);
  and (_22563_, _08548_, _23898_);
  and (_22564_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  or (_12706_, _22564_, _22563_);
  and (_22565_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  and (_22566_, _16331_, _23649_);
  or (_12711_, _22566_, _22565_);
  or (_22567_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_22568_, _22567_, _22762_);
  or (_22569_, _24079_, _23892_);
  and (_12717_, _22569_, _22568_);
  nand (_22570_, _24073_, _23772_);
  or (_22571_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_22572_, _22571_, _22762_);
  and (_12720_, _22572_, _22570_);
  and (_22573_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  and (_22574_, _16331_, _23747_);
  or (_26966_, _22574_, _22573_);
  and (_22575_, _25748_, _23707_);
  and (_22576_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_27070_, _22576_, _22575_);
  or (_22577_, _04891_, _23892_);
  and (_22578_, _26115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_22579_, _22578_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_22580_, _04880_, _26098_);
  and (_22581_, _22580_, _22579_);
  and (_22582_, _24300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_22583_, _22582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_22584_, _14815_);
  and (_22585_, _22584_, _24302_);
  and (_22586_, _22585_, _22583_);
  not (_22587_, _14810_);
  and (_22588_, _22587_, _04860_);
  or (_22589_, _22588_, _26100_);
  and (_22590_, _26110_, _26099_);
  and (_22591_, _22590_, _15862_);
  or (_22592_, _22591_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_22593_, _22592_, _22589_);
  or (_22594_, _22593_, _22586_);
  or (_22595_, _22594_, _22581_);
  or (_22596_, _22595_, _24299_);
  and (_22597_, _22596_, _24294_);
  and (_22598_, _22597_, _22577_);
  and (_22599_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_22600_, _22599_, _22598_);
  and (_12731_, _22600_, _22762_);
  not (_22601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_22602_, _26115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_22603_, _22602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_22604_, _22603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nand (_22605_, _22604_, _26099_);
  nand (_22606_, _22605_, _22601_);
  or (_22607_, _22605_, _22601_);
  and (_22608_, _22607_, _22606_);
  and (_22609_, _22608_, _04861_);
  or (_22610_, _24300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not (_22611_, _22582_);
  and (_22612_, _22611_, _24302_);
  and (_22613_, _22612_, _22610_);
  or (_22614_, _26115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_22615_, _22578_, _26098_);
  and (_22616_, _22615_, _22614_);
  or (_22617_, _22616_, _22613_);
  or (_22618_, _22617_, _22609_);
  or (_22619_, _22618_, _24299_);
  nand (_22620_, _24299_, _23772_);
  and (_22621_, _22620_, _24294_);
  and (_22622_, _22621_, _22619_);
  and (_22623_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_22624_, _22623_, _22622_);
  and (_12736_, _22624_, _22762_);
  and (_22625_, _05042_, _23649_);
  and (_22626_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_12741_, _22626_, _22625_);
  dff (first_instr, _00000_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _26843_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _26843_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _26843_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _26843_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _26843_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _26843_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _26843_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _26843_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _26859_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _26842_[1]);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _26842_[2]);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _26842_[3]);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _26842_[4]);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _26842_[5]);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _26842_[6]);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _26842_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _26842_[8]);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _26842_[9]);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _26842_[10]);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _26842_[11]);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _26842_[12]);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _26842_[13]);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _26842_[14]);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _26842_[15]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _26850_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _26850_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _26850_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _26850_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _26850_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _26850_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _26850_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _26850_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _26851_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _26851_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _26851_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _26851_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _26851_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _26851_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _26851_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _26851_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _26852_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _26852_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _26852_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _26852_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _26852_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _26852_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _26852_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _26852_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _26853_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _26853_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _26853_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _26853_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _26853_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _26853_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _26853_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _26853_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _26854_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _26854_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _26854_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _26854_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _26854_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _26854_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _26854_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _26854_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _26855_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _26855_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _26855_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _26855_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _26855_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _26855_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _26855_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _26855_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _26856_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _26856_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _26856_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _26856_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _26856_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _26856_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _26856_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _26856_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _26857_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _26857_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _26857_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _26857_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _26857_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _26857_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _26857_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _26857_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _26858_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _26858_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _26858_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _26858_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _26858_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _26858_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _26858_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _26858_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _26844_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _26844_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _26844_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _26844_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _26844_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _26844_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _26844_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _26844_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _26845_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _26845_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _26845_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _26845_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _26845_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _26845_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _26845_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _26845_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _26846_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _26846_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _26846_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _26846_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _26846_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _26846_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _26846_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _26846_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _26847_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _26847_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _26847_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _26847_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _26847_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _26847_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _26847_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _26847_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _26848_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _26848_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _26848_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _26848_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _26848_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _26848_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _26848_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _26848_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _26849_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _26849_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _26849_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _26849_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _26849_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _26849_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _26849_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _26849_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _11665_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _11643_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _09312_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _11604_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _11662_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _09317_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _09321_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _09302_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _11859_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _11759_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _11830_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _11817_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _11872_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _11857_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _11758_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _09315_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _12022_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22706_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _12035_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _12290_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _12040_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _12052_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _12026_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _12042_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _12048_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _12054_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _12050_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _12044_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _12037_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _12060_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _12056_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _12086_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _26860_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _26860_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _26860_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _26860_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _26860_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _26860_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _26860_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _26860_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _26887_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _26887_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _26887_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _26887_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _26887_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _26887_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _26887_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _26887_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _26897_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _26897_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _26897_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _26897_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _26897_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _26897_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _26897_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _26897_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _26867_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _26867_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _26868_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _26868_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _26868_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _26869_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _26869_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _26869_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _26870_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _26870_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _26871_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _26871_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _26871_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _26871_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _26872_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _26872_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _26873_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _26861_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _26861_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _26861_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _26862_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _26862_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _26862_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _26863_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _26863_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _26864_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _26864_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _26864_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _26864_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _26864_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _26864_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _26864_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _26864_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _26865_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _26866_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _26866_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _26912_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _26874_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _26874_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _26874_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _26874_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _26874_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _26874_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _26874_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _26874_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _26875_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _26875_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _26875_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _26875_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _26875_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _26875_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _26875_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _26875_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _26876_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _26876_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _26876_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _26876_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _26876_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _26876_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _26876_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _26876_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _26877_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _26877_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _26877_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _26877_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _26877_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _26877_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _26877_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _26877_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _26878_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _26878_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _26878_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _26878_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _26878_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _26878_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _26878_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _26878_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _26879_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _26879_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _26879_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _26879_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _26879_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _26879_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _26879_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _26879_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _26880_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _26880_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _26880_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _26880_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _26880_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _26880_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _26880_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _26880_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _26881_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _26881_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _26881_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _26881_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _26881_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _26881_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _26881_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _26881_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _26885_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _26885_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _26885_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _26885_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _26885_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _26882_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _26882_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _26882_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _26882_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _26882_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _26882_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _26882_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _26882_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _26882_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _26882_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _26882_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _26882_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _26882_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _26882_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _26882_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _26882_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _26883_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _26883_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _26883_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _26883_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _26883_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _26883_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _26883_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _26883_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _26883_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _26883_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _26883_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _26883_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _26883_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _26883_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _26883_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _26883_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _26903_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _26903_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _26903_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _26903_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _26903_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _26903_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _26903_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _26903_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _26903_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _26903_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _26903_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _26903_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _26903_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _26903_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _26903_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _26903_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _26903_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _26903_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _26903_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _26903_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _26903_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _26903_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _26903_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _26903_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _26903_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _26903_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _26903_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _26903_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _26903_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _26903_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _26903_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _26903_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _26884_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _26886_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _26886_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _26886_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _26886_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _26886_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _26886_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _26886_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _26886_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _26888_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _26889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _26890_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _26890_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _26890_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _26890_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _26890_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _26890_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _26890_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _26890_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _26890_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _26890_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _26890_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _26890_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _26890_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _26890_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _26890_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _26890_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _26891_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _26891_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _26891_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _26891_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _26891_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _26891_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _26891_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _26891_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _26891_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _26891_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _26891_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _26891_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _26891_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _26891_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _26891_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _26891_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _26892_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _26894_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _26893_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _26895_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _26895_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _26895_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _26895_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _26895_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _26895_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _26895_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _26895_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _26896_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _26896_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _26896_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _26898_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _26899_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _26899_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _26899_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _26899_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _26899_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _26899_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _26899_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _26899_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _26900_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _26901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _26902_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _26902_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _26902_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _26902_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _26904_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _26904_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _26904_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _26904_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _26904_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _26904_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _26904_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _26904_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _26904_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _26904_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _26904_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _26904_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _26904_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _26904_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _26904_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _26904_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _26904_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _26904_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _26904_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _26904_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _26904_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _26904_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _26904_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _26904_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _26904_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _26904_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _26904_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _26904_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _26904_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _26904_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _26904_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _26904_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _26905_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _26906_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _26907_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _26908_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _26908_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _26908_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _26908_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _26909_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _26910_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _26911_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _26911_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _26911_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _26911_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _26911_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _26911_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _26911_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _26911_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _26913_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _26913_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _26913_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _22681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _22683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _22682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _22703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _22701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _26992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _11711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _22673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _22880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _22863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _11715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _26978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _22705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _22740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _22727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _22726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _22959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _12237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _23125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _23119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _12234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _11791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _22759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _22758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _12226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _11793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _26942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _23210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _12232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _23297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _12228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _22993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _27008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _22675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _22677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _22676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _12241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _27009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _11867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _22656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _23507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _23513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _12224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _23566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _27301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _23406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _27302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _23388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _04653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _04647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _04638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _27156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _04733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _04716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _22694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _04697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _23723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _27138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _04779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _27139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _22697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _04818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _04847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _27140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _05321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _23410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _05465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _05456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _05451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _05503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _05498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _23650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _27199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _27200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _23685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _10452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _26771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _22715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _23162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _27201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _27196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _27197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _10416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _02571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _03365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _27198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _08203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _06170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _10399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _10737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _10390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _08205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _05707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _10406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _07531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _27195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _12185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _08175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _08442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _11698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _11783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _23426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _10377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _09523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _27193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _10342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _08208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _08909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _27194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _10355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _12101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _12292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _08210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _22714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _22723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _10336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _27192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _18519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _08749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _08765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _22704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _10310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _27191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _10770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _08179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _01784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _07708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _02210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _27189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _10280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _07185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _27190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _22925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _10297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _07402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _08181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _11617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _10015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _10138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _11458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _10291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _11456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _27188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _11615_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _11539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _27186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _09680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _27187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _11463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _09958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _11460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _09981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _09490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _11543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _09519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _11471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _27185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _11541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _09609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _09650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _10349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _10368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _09368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _10100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _10379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _09366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _27297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _10403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _09375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _10287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _10301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _27295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _09373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _27296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _10345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _09370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _11258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _11246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _27292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _27293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _27294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _11307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _11331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _11312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _27289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _11134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _09094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _27290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _27291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _11408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _11364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _11388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _11071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _08963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _11077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _27287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _08959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _09202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _11106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _27288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _27282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _27283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _08971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _27284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _08969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _27285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _09110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _27286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _09270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _10973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _27279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _08977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _27280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _08975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _27281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _09114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _09206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _10892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _10915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _08983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _10945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _08981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _10955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _09118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _10055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _11092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _12266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _11193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _11080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _12256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _12243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _12239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _10830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _09014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _10834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _10864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _09011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _27277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _09010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _10876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _11104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _11124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _09945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _11127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _11139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _09274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _26934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _26935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _09954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _26930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _09282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _11057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _09950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _26931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _26932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _26933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _09966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _26924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _26925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _09956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _26926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _26927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _26928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _26929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _26922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _09974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _10928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _10960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _09305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _10083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _26923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _09299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _09022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _07507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _07705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _05661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _05784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _07564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _05659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _07569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _07529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _08162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _08170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _07635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _08172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _26945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _07520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _08965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _06543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _06913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _07644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _06926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _07567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _07532_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _07712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _07625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _06562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _02062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _06664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _27161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _27162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _27163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _06368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _06342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _25152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _06784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _27159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _06915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _06891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _25147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _25673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _27160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _07278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _07253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _02013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _25575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _06986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _02033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _07092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _07089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _25747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _07359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _07338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _02008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _07435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _02003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _07191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _27158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _01104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _25458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _12284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _01833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _25457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _11117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _27157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _01837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _27154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _01750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _25758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _01806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _06103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _01789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _27155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _01344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _22698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _01761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _10856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _11267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _01780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _27153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _25492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _23328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _27152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _07658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _07633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _07611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _01991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _25578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _25771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _11834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _25589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _07729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _07719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _07777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _07797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _07781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _25288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _07523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _09038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _27150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _27151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _08103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _08092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _01976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _08429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _08118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _09191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _27149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _09952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _09387_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _25295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _08882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _08463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _08458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _10623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _25298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _10147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _27146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _27147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _01946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _27148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _09225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _27239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _08538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _27240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _08931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _11074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _26828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _26769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _07775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _25366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _10982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _10952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _01933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _27145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _25357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _10397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _01943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _11863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _27143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _11454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _27144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _11595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _11216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _11207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _11265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _27141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _11964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _12002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _12230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _27142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _01885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _11733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _11724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _27136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _12706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _12704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _01866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _12282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _01881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _27137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _01878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _23300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _27134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _27135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _25440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _12741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _09327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _01860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _25632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _27130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _05849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _03160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _27131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _23620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _27132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _27133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _03439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _06601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _27128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _06642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _03164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _07408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _00995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _27129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _03333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _03346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _27125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _12632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _27126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _04117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _27127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _07203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _03168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _03357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _03441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _22902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _24357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _27123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _23234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _27124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _10574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _27120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _03362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _07744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _22633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _27121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _22756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _27122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _06787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _22691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _07800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _08427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _26642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _26649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _26667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _27237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _27238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _27115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _27116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _27117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _22689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _22688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _27118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _22687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _27119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _02876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _22699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _03222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _22696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _02874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _22695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _03211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _22692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _07282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _27233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _09860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _07820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _11538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _04364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _22641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _23255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _07250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _07011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _07805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _22709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _27235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _22707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _22690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _27236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _03114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _08487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _03294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _03433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _22713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _02882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _22711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _03225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _00203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _03129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _09638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _03139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _10966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _03125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _27114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _03310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _22725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _27111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _27112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _27113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _22720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _03227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _03418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _11998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _01296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _01285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _27227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _01393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _27228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _27229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _08195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _23698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _27230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _23703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _00874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _01020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _00921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _27231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _27232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _10013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _27222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _09002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _09059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _08090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _08432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _08476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _05389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _05306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _27223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _27224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _05639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _10980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _03995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _03969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _03676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _05179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _25585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _12028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _11803_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _25487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _25478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _25535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _27082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _11738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _10920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _10895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _08094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _09919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _09906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _09900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _10360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _10938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _26914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _25617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _25614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _12024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _25658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _25648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _11754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _26915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _27203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _24502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _24499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _24496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _12072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _24395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _27204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _24387_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _25347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _11734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _24547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _24557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _24551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _12070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _24590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _12068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _25392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _25452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _25436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _12063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _24681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _27172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _24638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _12066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _24205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _11726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _23996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _24002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _23999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _12111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _24099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _24097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _24321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _24314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _12105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _24133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _24183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _27234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _12109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _24202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _24423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _24419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _24413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _24410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _11728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _11849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _24281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _12107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _23826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _23815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _23763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _23931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _23928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _27278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _12116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _11795_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _26664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _27108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _02906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _25180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _27109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _25177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _27110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _23176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _26731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _02972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _26726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _03270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _26720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _27107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _02923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _03391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _27106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _26834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _03108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _26805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _03287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _26764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _26748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _03046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _24330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _24580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _05568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _24583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _05573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _05842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _24603_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _24609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _05557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _27105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _05625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _05584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _05643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _24571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _24311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _24327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _27103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _05108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _27104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _03936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _05788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _05804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _05754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _05543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _04238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _05010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _05046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _05059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _27102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _05071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _04140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _05078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _04932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _27100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _04954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _27101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _03987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _04990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _03984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _04997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _27097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _27098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _04889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _04174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _04906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _04921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _04171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _04923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _04784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _04195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _04796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _04824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _27096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _04258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _04837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _04868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _04203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _04722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _04731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _04750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _04031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _04755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _04199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _27095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _04422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _04456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _04120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _04664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _04672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _04045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _04692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _04713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _04209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _04345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _04359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _04332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _04133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _04385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _04412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _04125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _04217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _04580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _04614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _04214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _04620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _27093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _27094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _04655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _04534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _04098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _04548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _27091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _04553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _04275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _27092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _04573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _05577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _04468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _04114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _04472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _04225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _04489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _04502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _27090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _25522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _05622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _25351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _25344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _25124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _25428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _25424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _25413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _24306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _25567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _05598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _25463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _25471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _25465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _05633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _25513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _24468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _05542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _24278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _24233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _24227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _24398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _24390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _24355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _05769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _25951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _25944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _25999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _24416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _24433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _05549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _24465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _25606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _25600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _27088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _25655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _25643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _25637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _27089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _25819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _25149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _25107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _05115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _03724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _25670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _27087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _25768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _25767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _01277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _01130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _05112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _01396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _01348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _03453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _11483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _11156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _05570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _27086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _01542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _01538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _05106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _03524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _03448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _05103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _05854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _05076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _09331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _09061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _27085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _05225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _04419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _04379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _05043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _10021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _05062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _10606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _27084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _05056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _06131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _05905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _11568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _11755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _05015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _10975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _27083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _10930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _05051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _11100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _22642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _22708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _22898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _05004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _03742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _11396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _11358_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _11280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _03605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _23207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _22998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _22719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _04988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _12674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _12615_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _12543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _25454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _25732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _04975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _27078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _01521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _04971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _03748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _27079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _03505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _27077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _02348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _02338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _04963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _04687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _04592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _03894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _09258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _27076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _03509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _07086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _05964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _04951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _08939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _07688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _09652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _09626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _09737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _09731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _04916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _09049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _09047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _04930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _03846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _27075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _09839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _09818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _10947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _10810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _10710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _03518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _27071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _27072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _04875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _11515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _11400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _11270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _27073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _27074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _04841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _27069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _22702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _04870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _02098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _04865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _03763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _27070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _09823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _03557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _03849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _02539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _04912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _03304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _04844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _05479_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _11659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _23189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _04798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _08215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _08951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _08947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _04827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _10206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _27068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _08826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _08828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _03574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _12509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _19972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _12613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _04803_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _08771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _22710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _22761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _08522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _08526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _03577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _09140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _27067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _09681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _07741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _00562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _23819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _04759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _03768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _08773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _08740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _27066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _03209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _26068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _05423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _04753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _22916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _04747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _26706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _04902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _03539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _07818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _06925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _07244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _27065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _09421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _24298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _27275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _10679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _27276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _09025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _10735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _10750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _10791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _09018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _10157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _09219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _10201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _10225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _10253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _09086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _10260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _09179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _10436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _27271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _09172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _10559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _27272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _10179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _27273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _27274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _09071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _09215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _10375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _10395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _09174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _10401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _10413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _09035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _10308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _09079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _10314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _27269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _10346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _09075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _27270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _09074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _11341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _27265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _27266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _27267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _11299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _22757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _27268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _10293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _27258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _27259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _27260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _27261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _27262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _11322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _27263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _27264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _27254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _03117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _12009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _11273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _07690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _27255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _27256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _27257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _27252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _11262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _16236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _22627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _16455_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _11244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _27253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _22660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _11356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _03855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _03788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _11394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _04742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _04519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _27251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _05258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _02903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _11353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _27247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _27248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _11418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _27249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _27250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _01716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _11189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _11183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _11136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _08190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _27246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _02437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _11404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _03083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _11255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _27243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _11132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _11368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _27244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _07746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _27245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _04080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _27241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _07752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _11489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _11473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _27242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _11591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _11534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _07750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _11102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _22724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _22693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _07771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _11721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _11718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _11696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _11853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _04610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _23554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _09433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _27205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _08496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _04849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _10227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _22679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _09156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _11548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _27182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _27183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _27184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _09277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _11545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _09338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _10196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _07300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _08188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _22716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _18188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _10165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _09887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _10163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _27179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _08852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _27180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _08908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _11478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _09009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _27181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _09081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _10646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _11694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _11526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _11425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _08115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _10182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _09184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _27202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _08572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _27177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _11487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _11621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _27178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _11485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _08777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _11562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _08202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _11924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _11911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _12273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _12294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _12277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _11230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _11153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _11569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _08365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _08416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _11493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _11622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _08466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _08544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _11491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _06542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _11613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _06585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _27175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _11532_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _11628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _08161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _27176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _07925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _11505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _11625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _07944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _08032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _11502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _08086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _08131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _27173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _07490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _11510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _27174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _07528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _07737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _11506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _07894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _11524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _06977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _11522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _07034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _11609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _07208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _11519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _27171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _06777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _04899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _04933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _04960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _23319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _27169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _27170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _11528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _22774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _22671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _00828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _04699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _27166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _27167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _04910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _27168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _27165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _12113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _04999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _04986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _22659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _05082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _05069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _05048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _27164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _05232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _05155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _05150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _05136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _05123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _05202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _05198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _27033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _21247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _21419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _21348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _27034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _22629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _22542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _12247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _05418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _05408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _23659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _05287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _05280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _05274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _27099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _05341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _27300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _10110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _10197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _10231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _09384_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _10240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _09379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _10258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _22640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _22637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _22658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _04530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _27041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _21820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _04550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _04542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _27042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _04562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _20570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _03664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _03871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _12920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _12950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _15784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _06171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _27020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _26054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _26057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _27021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _26059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _26066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _06100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _26981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _26982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _06660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _26983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _10194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _26984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _10304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _10289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _09382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _09309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _09296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _10104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _10036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _09991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _06864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _09101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _11164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _05546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _09837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _09359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _06705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _06611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _01901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _26980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _11161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _01372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _06709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _06528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _22835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _06714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _06711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _26962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _27298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _10454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _10511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _10569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _10625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _09357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _10172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _27299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _04409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _07854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _01524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _01495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _27225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _02826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _02446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _27226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _27219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _27220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _27221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _11203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _11200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _10897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _10784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _10799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _11236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _11228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _27217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _11497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _11468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _08107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _08435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _27218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _10813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _04851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _27214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _09923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _02714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _22685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _22684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _22670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _12477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _12288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _11882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _27215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _12586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _12545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _27216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _11222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _10838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _25628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _26780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _22639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _19920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _22636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _22638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _08110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _27209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _08439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _05185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _05689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _05300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _07535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _07290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _10755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _27213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _01820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _01566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _24697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _24449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _10832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _25792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _25972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _27210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _02362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _10797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _27211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _04640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _10780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _27212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _00764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _10748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _10650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _27206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _09668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _10706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _09753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _09733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _27207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _09254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _10731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _09612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _09600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _27208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _08995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _08943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _10745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _05902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _05673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _05587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _10652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _10604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _12268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _05386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _05370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _27080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _12258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _11091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _11051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _27081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _12264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _11792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _11681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _17981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _18303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _12252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _19421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _20043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _27058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _11787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _14938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _14601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _14450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _17417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _17267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _12254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _12344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _12223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _12805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _22661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _22669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _22662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _11707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _22632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _22631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _12245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _22635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _04802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _04719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _08089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _04710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _03792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _05383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _22787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _22678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _03880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _22722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _22643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _27063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _27064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _07342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _05815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _04689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _13798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _04670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _22628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _17600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _24247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _19941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _10888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _03613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _23504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _03703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _27060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _04446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _03701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _23248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _27061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _27062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _27050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _27051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _27052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _27053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _27054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _27055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _04651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _03802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _24200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _04330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _03883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _04400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _23586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _27059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _23477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _23517_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _04352_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _24091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _27056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _04382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _23891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _03713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _27057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _24106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _03542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _27046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _27047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _27048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _27049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _04645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _02060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _01953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _04361_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _04416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _04626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _27045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _05825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _03638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _02867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _02582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _04583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _08380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _08049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _07629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _04617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _09056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _09393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _04597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _22700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _04503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _27038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _22672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _27039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _27040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _22674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _04512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _03656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _11987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _04577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _27043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _27044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _03809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _10628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _04587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _03341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _06116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _25580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _23037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _23136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _27031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _27032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _22818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _22936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _27035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _22718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _22717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _27036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _22754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _04492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _27037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _03282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _03289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _27027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _27028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _03291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _03326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _27029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _27030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _03231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _05915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _03233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _06123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _06289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _03244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _27026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _05907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _05968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _03175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _05956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _03177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _06134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _03194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _05949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _03199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _02893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _02908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _05995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _02911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _27024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _05987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _06257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _02996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _03052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _06151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _03069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _03123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _27025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _06254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _03144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _05974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _06163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _01694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _06016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _01696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _27023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _02844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _02880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _06009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _00090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _00200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _27018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _06273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _00206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _00269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _06051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _00275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _26050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _06112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _00617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _06023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _00626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _06168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _27022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _01690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _00279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _06184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _00296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _27019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _00299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _06180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _00309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _00385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _06205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _26081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _26087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _06085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _06276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _26093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _26132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _06077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _27015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _04025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _27016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _07425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _03751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _07416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _26071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _27017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _03436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _03608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _27013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _07055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _26025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _27014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _03398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _03371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _03710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _03683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _03680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _07053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _03775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _03765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _06332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _03463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _06446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _06470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _02068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _25569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _06141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _06178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _06160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _02085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _04193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _04212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _06338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _03878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _03865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _04007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _04003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _03980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _04270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _27012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _04371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _04355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _06360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _04049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _04111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _04090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _04662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _04649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _04635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _04777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _04765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _04739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _07018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _04482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _27010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _04450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _04566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _27011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _04539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _07022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _06546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _04246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _05094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _06370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _04815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _04808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _04884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _04904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _04893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _06364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _27007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _06999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _06549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _05040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _05021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _05002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _05092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _05124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _06994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _05421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _05406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _27004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _27005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _05220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _27006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _05312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _06391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _05991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _05971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _05589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _26998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _06041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _06031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _06974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _05476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _05473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _26999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _27000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _27001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _27002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _06631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _27003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _06264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _06969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _26997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _06395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _06109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _06098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _06972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _06176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _06403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _06401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _06386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _06492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _06473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _06398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _06633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _06271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _06938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _06571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _06556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _06565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _06560_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _06965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _06617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _06640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _07061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _26994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _26995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _06635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _06869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _06859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _06837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _06932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _06917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _06911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _06415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _06707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _06695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _26996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _06758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _06765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _07195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _26993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _07173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _07150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _06430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _07013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _06929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _07081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _06923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _07287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _07310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _07305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _26991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _07098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _07110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _07106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _07396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _07390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _07363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _26989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _26990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _07428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _06440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _07246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _07739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _07851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _07823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _06450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _07640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _07638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _07617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _06901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _07694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _26987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _07495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _07491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _07485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _26988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _07561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _07538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _06457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _06638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _08100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _06887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _08424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _08421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _06885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _07765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _26985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _09228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _09194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _06461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _08454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _08449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _08988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _26986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _06684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _25285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _06679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _11884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _12672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _06689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _26979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _06702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _06824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _26976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _10370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _06833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _10599_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _26977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _06468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _06645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _11195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _26972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _26973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _06591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _10701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _26974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _06831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _26975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _06782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _06595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _11723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _26969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _11855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _06793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _26970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _11499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _11645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _06802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _06648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _11286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _06812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _11414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _06484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _26971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _12617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _06512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _26967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _12260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _12280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _26968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _11962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _06790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _12681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _12679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _06770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _26966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _12711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _06516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _12569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _12565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _06721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _26963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _26964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _11335_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _06748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _12249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _06523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _01928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _06754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _05700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _06121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _06521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _26965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _11684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _11410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _06519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _11119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _26961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _11141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _07445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _11147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _07441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _11149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _11159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _07587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _11062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _26959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _11083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _07453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _11094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _26960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _11109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _26952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _07607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _10958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _07487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _10968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _07604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _26953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _26954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _07602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _07724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _26955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _07481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _26956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _07598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _26957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _26958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _10192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _26950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _26951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _10221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _07498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _10806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _07614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _10902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _09167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _07627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _09291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _10089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _26948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _07702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _26949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _10188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _05862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _05899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _06088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _26946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _06093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _07680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _26947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _09112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _26943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _11349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _26944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _06526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _06535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _07540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _06537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _07654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _11289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _24175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _11296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _22746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _26939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _26940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _11346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _26941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _11315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _11329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _11317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _22866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _11242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _22680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _07579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _26938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _09340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _10844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _09988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _26920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _10880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _09334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _26921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _10886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _10239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _22686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _03822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _06233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _08183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _08451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _09854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _09821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _11406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _11374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _11376_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _24383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _11252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _26936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _26937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _11319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _26917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _09347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _10775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _26918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _26919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _10826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _09343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _10114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _10108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _10660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _09354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _10677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _10007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _26916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _10742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _09350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _22712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _11797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _04499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _03400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _04033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _22721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _11175_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _27303_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _27304_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _27304_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _27304_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _27304_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _27305_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _27306_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _27307_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _27307_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _27307_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _27307_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _27307_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _27307_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _27307_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _27307_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _10657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _10641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _10471_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _10500_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _10550_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _10516_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _10431_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _10353_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _06742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _06745_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _06744_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _06752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _06762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _06760_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _06767_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _05678_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _10133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _10132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _10097_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _10085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _10074_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _09940_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _10169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _09964_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _09976_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _10125_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _10050_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _10005_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _10130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _10128_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _10048_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _10143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _11762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _22664_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _09728_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _09843_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _09791_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _09772_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _09750_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22663_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _11828_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _09190_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _11565_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _11704_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _09127_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _22666_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _11663_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _09413_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _22665_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _11656_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _08672_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _08926_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _11683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _11577_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _11677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _11637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _08258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _08240_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _08221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _11651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _07683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _07512_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _07661_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _07595_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _07548_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _22667_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _07995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _11710_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _06934_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _06909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _06893_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _06844_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _22668_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _07281_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _07234_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _11687_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _12192_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _12170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _12139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _06267_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _12529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _12395_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _12507_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _11111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _11583_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _11558_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _11482_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _11413_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _06280_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _11954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _11878_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _11086_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _10891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _10718_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _10855_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _10829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _10779_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _10757_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _06293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _10940_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _10236_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _10212_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _10186_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _10161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _06326_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _10540_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _10409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _11053_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _10364_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _10338_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10329_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _10317_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _10330_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _10341_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _10039_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _06939_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _07222_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _07218_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _07231_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _07226_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _07228_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _07241_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _07237_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _06960_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _22634_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _01412_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _04590_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _11690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _11512_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _04585_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _00832_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _05875_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _03997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _06794_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _04624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _00740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _09365_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _15153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _12540_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _18600_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _26774_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _02663_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _22657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _10382_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _05196_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _03628_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _02555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _04642_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _10788_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _11085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _10873_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _22630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _12736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _12731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _04657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _23032_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _26617_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _26690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _09769_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _23573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _04338_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _12720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _12717_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _04659_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _26382_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _08395_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _15132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _17294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _06866_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _22655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _22654_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _04546_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _22653_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _07802_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _03406_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _07838_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _07834_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _07832_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _07830_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _07828_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _11891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _07779_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _07773_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _07769_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _07767_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _03409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _10384_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _07716_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _22652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _22648_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _03444_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _07656_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _07651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _07646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _03477_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _07699_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _07697_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _22647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _07596_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _07593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _03486_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _07630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _07609_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _07622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _07620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _22645_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _22644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _07549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _07546_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _03500_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _07575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _07565_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _07573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _07571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01438_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _23001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _23013_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _23010_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _23007_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _22760_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _22873_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _22752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _22753_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _22755_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _22776_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22790_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01419_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _01386_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _25815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _25814_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _01455_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _25874_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _25872_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _22851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _01452_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _22779_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _22792_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _22911_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _01384_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _22650_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _22651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _22955_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _22649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _22988_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _22933_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _22965_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _01407_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _25786_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _25778_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _25781_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _01466_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _22831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _22856_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _22858_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _25800_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _22751_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _22750_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _22749_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _22748_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _22747_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _22745_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _22744_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _22743_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _22742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _22741_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _25796_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _22739_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _22738_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _22646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _22737_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _04622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _22736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _22735_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _01457_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _22734_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _22733_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _22732_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _22731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _22730_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _22729_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _22728_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _01382_);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
endmodule
